
module alu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n226, n227, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621;

  HS65_LH_AND2X4 U157 ( .A(A[23]), .B(n587), .Z(n284) );
  HS65_LH_IVX9 U158 ( .A(B[1]), .Z(n580) );
  HS65_LH_OR2X9 U159 ( .A(B[29]), .B(n599), .Z(n294) );
  HS65_LH_IVX9 U160 ( .A(B[2]), .Z(n581) );
  HS65_LH_IVX9 U161 ( .A(B[23]), .Z(n587) );
  HS65_LH_IVX9 U162 ( .A(B[3]), .Z(n582) );
  HS65_LH_IVX9 U163 ( .A(B[22]), .Z(n586) );
  HS65_LH_IVX9 U164 ( .A(B[30]), .Z(n592) );
  HS65_LH_IVX9 U165 ( .A(A[14]), .Z(n596) );
  HS65_LH_IVX9 U166 ( .A(n304), .Z(n609) );
  HS65_LH_IVX9 U167 ( .A(A[8]), .Z(n594) );
  HS65_LH_IVX9 U168 ( .A(A[5]), .Z(n593) );
  HS65_LH_IVX9 U169 ( .A(A[17]), .Z(n597) );
  HS65_LH_IVX9 U170 ( .A(A[29]), .Z(n599) );
  HS65_LH_IVX9 U171 ( .A(A[20]), .Z(n598) );
  HS65_LH_IVX9 U172 ( .A(A[11]), .Z(n595) );
  HS65_LH_OAI32X5 U173 ( .A(n273), .B(n274), .C(n275), .D(n276), .E(n273), .Z(
        n272) );
  HS65_LH_OA22X9 U174 ( .A(n226), .B(n227), .C(n227), .D(n283), .Z(n274) );
  HS65_LH_CBI4I1X5 U175 ( .A(n600), .B(n601), .C(n286), .D(n287), .Z(n273) );
  HS65_LH_AOI212X4 U176 ( .A(n277), .B(n278), .C(n278), .D(n605), .E(n279), 
        .Z(n275) );
  HS65_LH_OAI21X3 U177 ( .A(n270), .B(n271), .C(n272), .Z(GE_LT_GT_LE) );
  HS65_LH_AOI312X4 U178 ( .A(n294), .B(n603), .C(B[28]), .D(B[29]), .E(n599), 
        .F(n295), .Z(n286) );
  HS65_LH_OAI212X5 U179 ( .A(n299), .B(n300), .C(n301), .D(n299), .E(n302), 
        .Z(n270) );
  HS65_LH_OA12X9 U180 ( .A(n606), .B(B[16]), .C(n282), .Z(n302) );
  HS65_LH_CBI4I1X5 U181 ( .A(n307), .B(n308), .C(n309), .D(n310), .Z(n300) );
  HS65_LH_NOR3X4 U182 ( .A(n303), .B(n304), .C(n305), .Z(n301) );
  HS65_LH_CBI4I1X5 U183 ( .A(n319), .B(n320), .C(n321), .D(n322), .Z(n299) );
  HS65_LH_OAI212X5 U184 ( .A(n323), .B(n324), .C(n613), .D(n323), .E(n609), 
        .Z(n322) );
  HS65_LH_AOI312X4 U185 ( .A(n325), .B(n612), .C(B[12]), .D(B[13]), .E(n611), 
        .F(n607), .Z(n321) );
  HS65_LH_IVX9 U186 ( .A(n305), .Z(n613) );
  HS65_LH_OAI211X5 U187 ( .A(B[12]), .B(n612), .C(n325), .D(n610), .Z(n304) );
  HS65_LH_IVX9 U188 ( .A(n320), .Z(n610) );
  HS65_LH_AOI32X5 U189 ( .A(n282), .B(n606), .C(B[16]), .D(B[17]), .E(n597), 
        .Z(n277) );
  HS65_LH_AOI12X2 U190 ( .A(n590), .B(A[26]), .C(n293), .Z(n290) );
  HS65_LH_OAI21X3 U191 ( .A(B[14]), .B(n596), .C(n327), .Z(n320) );
  HS65_LH_OAI211X5 U192 ( .A(B[20]), .B(n598), .C(n285), .D(n283), .Z(n279) );
  HS65_LH_OAI21X3 U193 ( .A(B[10]), .B(n614), .C(n326), .Z(n305) );
  HS65_LH_OAI21X3 U194 ( .A(B[6]), .B(n618), .C(n318), .Z(n308) );
  HS65_LH_NOR2X6 U195 ( .A(n593), .B(B[5]), .Z(n315) );
  HS65_LH_NAND3AX6 U196 ( .A(n279), .B(n280), .C(n276), .Z(n271) );
  HS65_LH_OA112X9 U197 ( .A(B[28]), .B(n603), .C(n294), .D(n296), .Z(n291) );
  HS65_LH_OAI21X3 U198 ( .A(B[8]), .B(n594), .C(n306), .Z(n303) );
  HS65_LH_AO32X4 U199 ( .A(B[10]), .B(n614), .C(n326), .D(n595), .E(B[11]), 
        .Z(n323) );
  HS65_LH_OR2X9 U200 ( .A(B[13]), .B(n611), .Z(n325) );
  HS65_LH_IVX9 U201 ( .A(n295), .Z(n600) );
  HS65_LH_AND2X4 U202 ( .A(B[31]), .B(n602), .Z(n297) );
  HS65_LH_OR2X9 U203 ( .A(B[17]), .B(n597), .Z(n282) );
  HS65_LH_OR2X9 U204 ( .A(B[21]), .B(n604), .Z(n285) );
  HS65_LH_AO32X4 U205 ( .A(n285), .B(n598), .C(B[20]), .D(B[21]), .E(n604), 
        .Z(n226) );
  HS65_LH_OR2X9 U206 ( .A(B[11]), .B(n595), .Z(n326) );
  HS65_LH_IVX9 U207 ( .A(B[4]), .Z(n583) );
  HS65_LH_IVX9 U208 ( .A(n319), .Z(n607) );
  HS65_LH_IVX9 U209 ( .A(n307), .Z(n616) );
  HS65_LH_IVX9 U210 ( .A(B[27]), .Z(n591) );
  HS65_LH_IVX9 U211 ( .A(B[26]), .Z(n590) );
  HS65_LH_IVX9 U212 ( .A(B[24]), .Z(n588) );
  HS65_LH_IVX9 U213 ( .A(B[19]), .Z(n585) );
  HS65_LH_IVX9 U214 ( .A(B[18]), .Z(n584) );
  HS65_LH_IVX9 U215 ( .A(n280), .Z(n605) );
  HS65_LH_IVX9 U216 ( .A(n296), .Z(n601) );
  HS65_LH_OAI32X5 U217 ( .A(n592), .B(A[30]), .C(n297), .D(B[31]), .E(n602), 
        .Z(n295) );
  HS65_LH_OAI32X5 U218 ( .A(n586), .B(A[22]), .C(n284), .D(A[23]), .E(n587), 
        .Z(n227) );
  HS65_LH_AOI312X4 U219 ( .A(n619), .B(n620), .C(B[4]), .D(B[5]), .E(n593), 
        .F(n616), .Z(n309) );
  HS65_LH_IVX9 U220 ( .A(A[4]), .Z(n620) );
  HS65_LH_IVX9 U221 ( .A(n315), .Z(n619) );
  HS65_LH_OAI212X5 U222 ( .A(n288), .B(n289), .C(n290), .D(n288), .E(n291), 
        .Z(n287) );
  HS65_LH_OAI32X5 U223 ( .A(n588), .B(A[24]), .C(n292), .D(A[25]), .E(n589), 
        .Z(n289) );
  HS65_LH_OAI32X5 U224 ( .A(n590), .B(A[26]), .C(n293), .D(A[27]), .E(n591), 
        .Z(n288) );
  HS65_LH_IVX9 U225 ( .A(B[25]), .Z(n589) );
  HS65_LH_AOI32X5 U226 ( .A(B[14]), .B(n596), .C(n327), .D(n608), .E(B[15]), 
        .Z(n319) );
  HS65_LH_IVX9 U227 ( .A(A[15]), .Z(n608) );
  HS65_LH_AOI32X5 U228 ( .A(B[6]), .B(n618), .C(n318), .D(n617), .E(B[7]), .Z(
        n307) );
  HS65_LH_IVX9 U229 ( .A(A[7]), .Z(n617) );
  HS65_LH_AOI12X2 U230 ( .A(n584), .B(A[18]), .C(n281), .Z(n280) );
  HS65_LH_AOI22X6 U231 ( .A(B[1]), .B(n621), .C(n316), .D(B[0]), .Z(n313) );
  HS65_LH_IVX9 U232 ( .A(A[1]), .Z(n621) );
  HS65_LH_AOI12X2 U233 ( .A(A[1]), .B(n580), .C(A[0]), .Z(n316) );
  HS65_LH_AOI12X2 U234 ( .A(n586), .B(A[22]), .C(n284), .Z(n283) );
  HS65_LH_NOR2AX3 U235 ( .A(A[25]), .B(B[25]), .Z(n292) );
  HS65_LH_NAND3AX6 U236 ( .A(n308), .B(n311), .C(n312), .Z(n310) );
  HS65_LH_CBI4I1X5 U237 ( .A(A[2]), .B(n581), .C(n317), .D(n314), .Z(n311) );
  HS65_LH_AOI212X4 U238 ( .A(n313), .B(n314), .C(A[4]), .D(n583), .E(n315), 
        .Z(n312) );
  HS65_LH_OA32X4 U239 ( .A(n581), .B(A[2]), .C(n317), .D(A[3]), .E(n582), .Z(
        n314) );
  HS65_LH_AOI12X2 U240 ( .A(n592), .B(A[30]), .C(n297), .Z(n296) );
  HS65_LH_OA32X4 U241 ( .A(n584), .B(A[18]), .C(n281), .D(A[19]), .E(n585), 
        .Z(n278) );
  HS65_LH_NAND2AX7 U242 ( .A(B[15]), .B(A[15]), .Z(n327) );
  HS65_LH_NAND2AX7 U243 ( .A(B[7]), .B(A[7]), .Z(n318) );
  HS65_LH_NAND2AX7 U244 ( .A(B[9]), .B(A[9]), .Z(n306) );
  HS65_LH_AND2X4 U245 ( .A(A[27]), .B(n591), .Z(n293) );
  HS65_LH_AO32X4 U246 ( .A(B[8]), .B(n594), .C(n306), .D(n615), .E(B[9]), .Z(
        n324) );
  HS65_LH_IVX9 U247 ( .A(A[9]), .Z(n615) );
  HS65_LH_AND3X9 U248 ( .A(n290), .B(n291), .C(n298), .Z(n276) );
  HS65_LH_AOI12X2 U249 ( .A(A[24]), .B(n588), .C(n292), .Z(n298) );
  HS65_LH_AND2X4 U250 ( .A(A[3]), .B(n582), .Z(n317) );
  HS65_LH_AND2X4 U251 ( .A(A[19]), .B(n585), .Z(n281) );
  HS65_LH_IVX9 U252 ( .A(A[12]), .Z(n612) );
  HS65_LH_IVX9 U253 ( .A(A[6]), .Z(n618) );
  HS65_LH_IVX9 U254 ( .A(A[13]), .Z(n611) );
  HS65_LH_IVX9 U255 ( .A(A[16]), .Z(n606) );
  HS65_LH_IVX9 U256 ( .A(A[31]), .Z(n602) );
  HS65_LH_IVX9 U257 ( .A(A[10]), .Z(n614) );
  HS65_LH_IVX9 U258 ( .A(A[28]), .Z(n603) );
  HS65_LH_IVX9 U259 ( .A(A[21]), .Z(n604) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253;
  wire   [32:0] carry;

  HS65_LH_FA1X4 U2_30 ( .A0(A[30]), .B0(n252), .CI(carry[30]), .CO(carry[31]), 
        .S0(DIFF[30]) );
  HS65_LH_FA1X4 U2_28 ( .A0(A[28]), .B0(n250), .CI(carry[28]), .CO(carry[29]), 
        .S0(DIFF[28]) );
  HS65_LH_FA1X4 U2_27 ( .A0(A[27]), .B0(n249), .CI(carry[27]), .CO(carry[28]), 
        .S0(DIFF[27]) );
  HS65_LH_FA1X4 U2_22 ( .A0(A[22]), .B0(n244), .CI(carry[22]), .CO(carry[23]), 
        .S0(DIFF[22]) );
  HS65_LH_FA1X4 U2_19 ( .A0(A[19]), .B0(n241), .CI(carry[19]), .CO(carry[20]), 
        .S0(DIFF[19]) );
  HS65_LH_FA1X4 U2_18 ( .A0(A[18]), .B0(n240), .CI(carry[18]), .CO(carry[19]), 
        .S0(DIFF[18]) );
  HS65_LH_FA1X4 U2_16 ( .A0(A[16]), .B0(n238), .CI(carry[16]), .CO(carry[17]), 
        .S0(DIFF[16]) );
  HS65_LH_FA1X4 U2_15 ( .A0(A[15]), .B0(n237), .CI(carry[15]), .CO(carry[16]), 
        .S0(DIFF[15]) );
  HS65_LH_FA1X4 U2_13 ( .A0(A[13]), .B0(n235), .CI(carry[13]), .CO(carry[14]), 
        .S0(DIFF[13]) );
  HS65_LH_FA1X4 U2_12 ( .A0(A[12]), .B0(n234), .CI(carry[12]), .CO(carry[13]), 
        .S0(DIFF[12]) );
  HS65_LH_FA1X4 U2_10 ( .A0(A[10]), .B0(n232), .CI(carry[10]), .CO(carry[11]), 
        .S0(DIFF[10]) );
  HS65_LH_FA1X4 U2_9 ( .A0(A[9]), .B0(n231), .CI(carry[9]), .CO(carry[10]), 
        .S0(DIFF[9]) );
  HS65_LH_FA1X4 U2_7 ( .A0(A[7]), .B0(n229), .CI(carry[7]), .CO(carry[8]), 
        .S0(DIFF[7]) );
  HS65_LH_FA1X4 U2_6 ( .A0(A[6]), .B0(n228), .CI(carry[6]), .CO(carry[7]), 
        .S0(DIFF[6]) );
  HS65_LH_FA1X4 U2_4 ( .A0(A[4]), .B0(n226), .CI(carry[4]), .CO(carry[5]), 
        .S0(DIFF[4]) );
  HS65_LH_FA1X4 U2_3 ( .A0(A[3]), .B0(n225), .CI(carry[3]), .CO(carry[4]), 
        .S0(DIFF[3]) );
  HS65_LH_FA1X4 U2_25 ( .A0(A[25]), .B0(n247), .CI(carry[25]), .CO(carry[26]), 
        .S0(DIFF[25]) );
  HS65_LH_FA1X4 U2_21 ( .A0(A[21]), .B0(n243), .CI(carry[21]), .CO(carry[22]), 
        .S0(DIFF[21]) );
  HS65_LH_FA1X4 U2_1 ( .A0(A[1]), .B0(n223), .CI(carry[1]), .CO(carry[2]), 
        .S0(DIFF[1]) );
  HS65_LH_FA1X4 U2_24 ( .A0(A[24]), .B0(n246), .CI(carry[24]), .CO(carry[25]), 
        .S0(DIFF[24]) );
  HS65_LH_FA1X4 U2_2 ( .A0(A[2]), .B0(n224), .CI(carry[2]), .CO(carry[3]), 
        .S0(DIFF[2]) );
  HS65_LH_FA1X4 U2_23 ( .A0(A[23]), .B0(n245), .CI(carry[23]), .CO(carry[24]), 
        .S0(DIFF[23]) );
  HS65_LH_FA1X4 U2_26 ( .A0(A[26]), .B0(n248), .CI(carry[26]), .CO(carry[27]), 
        .S0(DIFF[26]) );
  HS65_LH_FA1X4 U2_20 ( .A0(A[20]), .B0(n242), .CI(carry[20]), .CO(carry[21]), 
        .S0(DIFF[20]) );
  HS65_LH_FA1X4 U2_29 ( .A0(A[29]), .B0(n251), .CI(carry[29]), .CO(carry[30]), 
        .S0(DIFF[29]) );
  HS65_LH_FA1X4 U2_17 ( .A0(A[17]), .B0(n239), .CI(carry[17]), .CO(carry[18]), 
        .S0(DIFF[17]) );
  HS65_LH_FA1X4 U2_11 ( .A0(A[11]), .B0(n233), .CI(carry[11]), .CO(carry[12]), 
        .S0(DIFF[11]) );
  HS65_LH_FA1X4 U2_5 ( .A0(A[5]), .B0(n227), .CI(carry[5]), .CO(carry[6]), 
        .S0(DIFF[5]) );
  HS65_LH_FA1X4 U2_14 ( .A0(A[14]), .B0(n236), .CI(carry[14]), .CO(carry[15]), 
        .S0(DIFF[14]) );
  HS65_LH_FA1X4 U2_8 ( .A0(A[8]), .B0(n230), .CI(carry[8]), .CO(carry[9]), 
        .S0(DIFF[8]) );
  HS65_LH_IVX9 U1 ( .A(B[8]), .Z(n230) );
  HS65_LH_IVX9 U2 ( .A(B[14]), .Z(n236) );
  HS65_LH_IVX9 U3 ( .A(B[5]), .Z(n227) );
  HS65_LH_IVX9 U4 ( .A(B[11]), .Z(n233) );
  HS65_LH_IVX9 U5 ( .A(B[17]), .Z(n239) );
  HS65_LH_IVX9 U6 ( .A(B[29]), .Z(n251) );
  HS65_LH_IVX9 U7 ( .A(B[20]), .Z(n242) );
  HS65_LH_IVX9 U8 ( .A(B[26]), .Z(n248) );
  HS65_LH_IVX9 U9 ( .A(B[23]), .Z(n245) );
  HS65_LH_IVX9 U10 ( .A(B[2]), .Z(n224) );
  HS65_LHS_XNOR3X2 U11 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Z(DIFF[31]) );
  HS65_LHS_XOR2X6 U12 ( .A(A[0]), .B(B[0]), .Z(DIFF[0]) );
  HS65_LH_IVX9 U13 ( .A(B[24]), .Z(n246) );
  HS65_LH_IVX9 U14 ( .A(B[1]), .Z(n223) );
  HS65_LH_NAND2X7 U15 ( .A(n253), .B(B[0]), .Z(carry[1]) );
  HS65_LH_IVX9 U16 ( .A(A[0]), .Z(n253) );
  HS65_LH_IVX9 U17 ( .A(B[21]), .Z(n243) );
  HS65_LH_IVX9 U18 ( .A(B[25]), .Z(n247) );
  HS65_LH_IVX9 U19 ( .A(B[3]), .Z(n225) );
  HS65_LH_IVX9 U20 ( .A(B[4]), .Z(n226) );
  HS65_LH_IVX9 U21 ( .A(B[6]), .Z(n228) );
  HS65_LH_IVX9 U22 ( .A(B[7]), .Z(n229) );
  HS65_LH_IVX9 U23 ( .A(B[9]), .Z(n231) );
  HS65_LH_IVX9 U24 ( .A(B[10]), .Z(n232) );
  HS65_LH_IVX9 U25 ( .A(B[12]), .Z(n234) );
  HS65_LH_IVX9 U26 ( .A(B[13]), .Z(n235) );
  HS65_LH_IVX9 U27 ( .A(B[15]), .Z(n237) );
  HS65_LH_IVX9 U28 ( .A(B[16]), .Z(n238) );
  HS65_LH_IVX9 U29 ( .A(B[18]), .Z(n240) );
  HS65_LH_IVX9 U30 ( .A(B[19]), .Z(n241) );
  HS65_LH_IVX9 U31 ( .A(B[22]), .Z(n244) );
  HS65_LH_IVX9 U32 ( .A(B[27]), .Z(n249) );
  HS65_LH_IVX9 U33 ( .A(B[28]), .Z(n250) );
  HS65_LH_IVX9 U34 ( .A(B[30]), .Z(n252) );
endmodule


module alu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405;

  HS65_LH_NAND2X7 U1 ( .A(A[5]), .B(n366), .Z(n106) );
  HS65_LH_NAND2X7 U2 ( .A(A[29]), .B(n381), .Z(n62) );
  HS65_LH_NAND2X7 U3 ( .A(A[11]), .B(n369), .Z(n54) );
  HS65_LH_NAND2X7 U4 ( .A(A[20]), .B(n375), .Z(n74) );
  HS65_LH_NAND2X7 U5 ( .A(A[23]), .B(n377), .Z(n72) );
  HS65_LH_NAND2X7 U6 ( .A(A[17]), .B(n373), .Z(n69) );
  HS65_LH_IVX9 U7 ( .A(B[3]), .Z(n365) );
  HS65_LH_IVX9 U8 ( .A(B[2]), .Z(n364) );
  HS65_LH_IVX9 U9 ( .A(B[23]), .Z(n377) );
  HS65_LH_IVX9 U10 ( .A(B[29]), .Z(n381) );
  HS65_LH_IVX9 U11 ( .A(A[8]), .Z(n383) );
  HS65_LH_IVX9 U12 ( .A(B[31]), .Z(n382) );
  HS65_LH_IVX9 U13 ( .A(A[14]), .Z(n384) );
  HS65_LH_IVX9 U14 ( .A(A[26]), .Z(n385) );
  HS65_LH_IVX9 U15 ( .A(n115), .Z(n403) );
  HS65_LH_NOR4ABX2 U16 ( .A(n76), .B(n77), .C(n78), .D(LT), .Z(n43) );
  HS65_LH_AND2X4 U17 ( .A(n114), .B(n109), .Z(n77) );
  HS65_LH_NAND4ABX3 U18 ( .A(n115), .B(n401), .C(n106), .D(n105), .Z(n78) );
  HS65_LH_IVX9 U19 ( .A(n102), .Z(n401) );
  HS65_LH_NOR4ABX2 U20 ( .A(n55), .B(n56), .C(n57), .D(n58), .Z(n44) );
  HS65_LH_AND4X6 U21 ( .A(n72), .B(n73), .C(n74), .D(n75), .Z(n55) );
  HS65_LH_NAND4ABX3 U22 ( .A(n59), .B(n60), .C(n61), .D(n62), .Z(n58) );
  HS65_LH_NAND4ABX3 U23 ( .A(n64), .B(n390), .C(n65), .D(n66), .Z(n57) );
  HS65_LH_NOR4ABX2 U24 ( .A(n68), .B(n69), .C(n70), .D(n71), .Z(n56) );
  HS65_LH_NOR2X6 U25 ( .A(B[18]), .B(n395), .Z(n70) );
  HS65_LH_NAND4ABX3 U26 ( .A(n51), .B(n398), .C(n52), .D(n53), .Z(n45) );
  HS65_LH_IVX9 U27 ( .A(n54), .Z(n398) );
  HS65_LH_NOR2X6 U28 ( .A(n397), .B(B[16]), .Z(n71) );
  HS65_LH_NOR2X6 U29 ( .A(n389), .B(B[30]), .Z(n60) );
  HS65_LH_NOR2X6 U30 ( .A(n404), .B(B[4]), .Z(n115) );
  HS65_LH_NOR2X6 U31 ( .A(n392), .B(B[24]), .Z(n64) );
  HS65_LH_NOR2X6 U32 ( .A(n383), .B(B[8]), .Z(n51) );
  HS65_LH_IVX9 U33 ( .A(EQ), .Z(NE) );
  HS65_LH_NOR4ABX2 U34 ( .A(n43), .B(n44), .C(n45), .D(n46), .Z(EQ) );
  HS65_LH_OR2X9 U35 ( .A(B[26]), .B(n385), .Z(n66) );
  HS65_LH_NAND2X7 U36 ( .A(A[2]), .B(n364), .Z(n114) );
  HS65_LH_OR2X9 U37 ( .A(B[14]), .B(n384), .Z(n50) );
  HS65_LH_IVX9 U38 ( .A(B[19]), .Z(n374) );
  HS65_LH_IVX9 U39 ( .A(B[27]), .Z(n379) );
  HS65_LH_IVX9 U40 ( .A(B[25]), .Z(n378) );
  HS65_LH_IVX9 U41 ( .A(B[12]), .Z(n370) );
  HS65_LH_IVX9 U42 ( .A(B[15]), .Z(n372) );
  HS65_LH_IVX9 U43 ( .A(B[20]), .Z(n375) );
  HS65_LH_IVX9 U44 ( .A(B[13]), .Z(n371) );
  HS65_LH_IVX9 U45 ( .A(B[5]), .Z(n366) );
  HS65_LH_IVX9 U46 ( .A(B[17]), .Z(n373) );
  HS65_LH_IVX9 U47 ( .A(B[7]), .Z(n367) );
  HS65_LH_IVX9 U48 ( .A(B[11]), .Z(n369) );
  HS65_LH_IVX9 U49 ( .A(B[28]), .Z(n380) );
  HS65_LH_IVX9 U50 ( .A(B[21]), .Z(n376) );
  HS65_LH_IVX9 U51 ( .A(B[9]), .Z(n368) );
  HS65_LH_NAND4X9 U52 ( .A(n47), .B(n48), .C(n49), .D(n50), .Z(n46) );
  HS65_LH_IVX9 U53 ( .A(n67), .Z(n390) );
  HS65_LH_OAI22X6 U54 ( .A(A[31]), .B(n382), .C(n387), .D(n79), .Z(LT) );
  HS65_LH_IVX9 U55 ( .A(n76), .Z(n387) );
  HS65_LH_AOI32X5 U56 ( .A(n62), .B(n388), .C(n80), .D(B[30]), .E(n389), .Z(
        n79) );
  HS65_LH_IVX9 U57 ( .A(n60), .Z(n388) );
  HS65_LH_OAI212X5 U58 ( .A(A[2]), .B(n364), .C(A[3]), .D(n365), .E(n111), .Z(
        n110) );
  HS65_LH_OAI212X5 U59 ( .A(B[1]), .B(n112), .C(n113), .D(n405), .E(n114), .Z(
        n111) );
  HS65_LH_AND2X4 U60 ( .A(n113), .B(n405), .Z(n112) );
  HS65_LH_NOR2AX3 U61 ( .A(B[0]), .B(A[0]), .Z(n113) );
  HS65_LH_OAI212X5 U62 ( .A(A[12]), .B(n370), .C(A[13]), .D(n371), .E(n97), 
        .Z(n96) );
  HS65_LH_NAND3X5 U63 ( .A(n47), .B(n54), .C(n98), .Z(n97) );
  HS65_LH_OAI21X3 U64 ( .A(A[11]), .B(n369), .C(n99), .Z(n98) );
  HS65_LH_AOI32X5 U65 ( .A(n53), .B(n52), .C(n100), .D(B[10]), .E(n399), .Z(
        n99) );
  HS65_LH_OAI212X5 U66 ( .A(A[28]), .B(n380), .C(A[29]), .D(n381), .E(n81), 
        .Z(n80) );
  HS65_LH_NAND3X5 U67 ( .A(n61), .B(n67), .C(n82), .Z(n81) );
  HS65_LH_OAI21X3 U68 ( .A(A[27]), .B(n379), .C(n83), .Z(n82) );
  HS65_LH_AOI32X5 U69 ( .A(n66), .B(n65), .C(n84), .D(B[26]), .E(n385), .Z(n83) );
  HS65_LH_AOI32X5 U70 ( .A(n73), .B(n75), .C(n88), .D(B[22]), .E(n393), .Z(n87) );
  HS65_LH_IVX9 U71 ( .A(A[22]), .Z(n393) );
  HS65_LH_OAI212X5 U72 ( .A(A[20]), .B(n375), .C(A[21]), .D(n376), .E(n89), 
        .Z(n88) );
  HS65_LH_NAND3X5 U73 ( .A(n74), .B(n68), .C(n90), .Z(n89) );
  HS65_LH_AOI32X5 U74 ( .A(n396), .B(n49), .C(n94), .D(B[16]), .E(n397), .Z(
        n93) );
  HS65_LH_IVX9 U75 ( .A(n71), .Z(n396) );
  HS65_LH_OAI21X3 U76 ( .A(A[15]), .B(n372), .C(n95), .Z(n94) );
  HS65_LH_AOI32X5 U77 ( .A(n50), .B(n48), .C(n96), .D(B[14]), .E(n384), .Z(n95) );
  HS65_LH_AOI32X5 U78 ( .A(n105), .B(n106), .C(n107), .D(B[6]), .E(n402), .Z(
        n104) );
  HS65_LH_IVX9 U79 ( .A(A[6]), .Z(n402) );
  HS65_LH_OAI21X3 U80 ( .A(A[5]), .B(n366), .C(n108), .Z(n107) );
  HS65_LH_AOI32X5 U81 ( .A(n403), .B(n109), .C(n110), .D(B[4]), .E(n404), .Z(
        n108) );
  HS65_LH_AOI22X6 U82 ( .A(n405), .B(n63), .C(n63), .D(B[1]), .Z(n59) );
  HS65_LH_NAND2AX7 U83 ( .A(B[0]), .B(A[0]), .Z(n63) );
  HS65_LH_OAI21X3 U84 ( .A(A[25]), .B(n378), .C(n85), .Z(n84) );
  HS65_LH_AOI32X5 U85 ( .A(n391), .B(n72), .C(n86), .D(B[24]), .E(n392), .Z(
        n85) );
  HS65_LH_IVX9 U86 ( .A(n64), .Z(n391) );
  HS65_LH_OAI21X3 U87 ( .A(A[23]), .B(n377), .C(n87), .Z(n86) );
  HS65_LH_OAI21X3 U88 ( .A(A[9]), .B(n368), .C(n101), .Z(n100) );
  HS65_LH_AOI32X5 U89 ( .A(n400), .B(n102), .C(n103), .D(B[8]), .E(n383), .Z(
        n101) );
  HS65_LH_IVX9 U90 ( .A(n51), .Z(n400) );
  HS65_LH_OAI21X3 U91 ( .A(A[7]), .B(n367), .C(n104), .Z(n103) );
  HS65_LH_OAI21X3 U92 ( .A(A[19]), .B(n374), .C(n91), .Z(n90) );
  HS65_LH_AOI32X5 U93 ( .A(n394), .B(n69), .C(n92), .D(B[18]), .E(n395), .Z(
        n91) );
  HS65_LH_IVX9 U94 ( .A(n70), .Z(n394) );
  HS65_LH_OAI21X3 U95 ( .A(A[17]), .B(n373), .C(n93), .Z(n92) );
  HS65_LH_NAND2AX7 U96 ( .A(B[6]), .B(A[6]), .Z(n105) );
  HS65_LH_NAND2AX7 U97 ( .A(B[10]), .B(A[10]), .Z(n53) );
  HS65_LH_NAND2AX7 U98 ( .A(B[22]), .B(A[22]), .Z(n73) );
  HS65_LH_NAND2X7 U99 ( .A(A[28]), .B(n380), .Z(n61) );
  HS65_LH_NAND2X7 U100 ( .A(A[25]), .B(n378), .Z(n65) );
  HS65_LH_NAND2X7 U101 ( .A(A[9]), .B(n368), .Z(n52) );
  HS65_LH_NAND2X7 U102 ( .A(A[27]), .B(n379), .Z(n67) );
  HS65_LH_NAND2X7 U103 ( .A(A[7]), .B(n367), .Z(n102) );
  HS65_LH_NAND2X7 U104 ( .A(A[19]), .B(n374), .Z(n68) );
  HS65_LH_NAND2X7 U105 ( .A(A[3]), .B(n365), .Z(n109) );
  HS65_LH_NAND2X7 U106 ( .A(A[21]), .B(n376), .Z(n75) );
  HS65_LH_NAND2X7 U107 ( .A(A[31]), .B(n382), .Z(n76) );
  HS65_LH_NAND2X7 U108 ( .A(A[12]), .B(n370), .Z(n47) );
  HS65_LH_NAND2X7 U109 ( .A(A[13]), .B(n371), .Z(n48) );
  HS65_LH_NAND2X7 U110 ( .A(A[15]), .B(n372), .Z(n49) );
  HS65_LH_IVX9 U111 ( .A(A[1]), .Z(n405) );
  HS65_LH_IVX9 U112 ( .A(A[4]), .Z(n404) );
  HS65_LH_IVX9 U113 ( .A(A[16]), .Z(n397) );
  HS65_LH_IVX9 U114 ( .A(A[24]), .Z(n392) );
  HS65_LH_IVX9 U115 ( .A(A[30]), .Z(n389) );
  HS65_LH_IVX9 U116 ( .A(A[18]), .Z(n395) );
  HS65_LH_IVX9 U117 ( .A(A[10]), .Z(n399) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  HS65_LH_FA1X4 U1_30 ( .A0(A[30]), .B0(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S0(SUM[30]) );
  HS65_LH_FA1X4 U1_28 ( .A0(A[28]), .B0(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S0(SUM[28]) );
  HS65_LH_FA1X4 U1_27 ( .A0(A[27]), .B0(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S0(SUM[27]) );
  HS65_LH_FA1X4 U1_25 ( .A0(A[25]), .B0(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S0(SUM[25]) );
  HS65_LH_FA1X4 U1_24 ( .A0(A[24]), .B0(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S0(SUM[24]) );
  HS65_LH_FA1X4 U1_22 ( .A0(A[22]), .B0(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S0(SUM[22]) );
  HS65_LH_FA1X4 U1_21 ( .A0(A[21]), .B0(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S0(SUM[21]) );
  HS65_LH_FA1X4 U1_19 ( .A0(A[19]), .B0(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S0(SUM[19]) );
  HS65_LH_FA1X4 U1_18 ( .A0(A[18]), .B0(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S0(SUM[18]) );
  HS65_LH_FA1X4 U1_12 ( .A0(A[12]), .B0(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S0(SUM[12]) );
  HS65_LH_FA1X4 U1_10 ( .A0(A[10]), .B0(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S0(SUM[10]) );
  HS65_LH_FA1X4 U1_9 ( .A0(A[9]), .B0(B[9]), .CI(carry[9]), .CO(carry[10]), 
        .S0(SUM[9]) );
  HS65_LH_FA1X4 U1_7 ( .A0(A[7]), .B0(B[7]), .CI(carry[7]), .CO(carry[8]), 
        .S0(SUM[7]) );
  HS65_LH_FA1X4 U1_6 ( .A0(A[6]), .B0(B[6]), .CI(carry[6]), .CO(carry[7]), 
        .S0(SUM[6]) );
  HS65_LH_FA1X4 U1_4 ( .A0(A[4]), .B0(B[4]), .CI(carry[4]), .CO(carry[5]), 
        .S0(SUM[4]) );
  HS65_LH_FA1X4 U1_3 ( .A0(A[3]), .B0(B[3]), .CI(carry[3]), .CO(carry[4]), 
        .S0(SUM[3]) );
  HS65_LH_FA1X4 U1_16 ( .A0(A[16]), .B0(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S0(SUM[16]) );
  HS65_LH_FA1X4 U1_1 ( .A0(A[1]), .B0(B[1]), .CI(n1), .CO(carry[2]), .S0(
        SUM[1]) );
  HS65_LH_FA1X4 U1_15 ( .A0(A[15]), .B0(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S0(SUM[15]) );
  HS65_LH_FA1X4 U1_13 ( .A0(A[13]), .B0(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S0(SUM[13]) );
  HS65_LHS_XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Z(SUM[31]) );
  HS65_LH_FA1X4 U1_2 ( .A0(A[2]), .B0(B[2]), .CI(carry[2]), .CO(carry[3]), 
        .S0(SUM[2]) );
  HS65_LH_FA1X4 U1_23 ( .A0(A[23]), .B0(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S0(SUM[23]) );
  HS65_LH_FA1X4 U1_29 ( .A0(A[29]), .B0(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S0(SUM[29]) );
  HS65_LH_FA1X4 U1_26 ( .A0(A[26]), .B0(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S0(SUM[26]) );
  HS65_LH_FA1X4 U1_20 ( .A0(A[20]), .B0(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S0(SUM[20]) );
  HS65_LH_FA1X4 U1_17 ( .A0(A[17]), .B0(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S0(SUM[17]) );
  HS65_LH_FA1X4 U1_11 ( .A0(A[11]), .B0(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S0(SUM[11]) );
  HS65_LH_FA1X4 U1_5 ( .A0(A[5]), .B0(B[5]), .CI(carry[5]), .CO(carry[6]), 
        .S0(SUM[5]) );
  HS65_LH_FA1X4 U1_8 ( .A0(A[8]), .B0(B[8]), .CI(carry[8]), .CO(carry[9]), 
        .S0(SUM[8]) );
  HS65_LH_FA1X4 U1_14 ( .A0(A[14]), .B0(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S0(SUM[14]) );
  HS65_LHS_XOR2X6 U1 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  HS65_LH_AND2X4 U2 ( .A(A[0]), .B(B[0]), .Z(n1) );
endmodule


module alu_DW_mult_uns_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n7, n19, n31, n43, n55, n67, n79, n91, n103, n115, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n292, n293, n294, n295, n296, n297,
         n299, n300, n302, n303, n304, n305, n306, n307, n308, n309, n311,
         n312, n313, n314, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
         n360, n361, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n2417, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719;
  assign n7 = a[2];
  assign n19 = a[5];
  assign n31 = a[8];
  assign n43 = a[11];
  assign n55 = a[14];
  assign n67 = a[17];
  assign n79 = a[20];
  assign n91 = a[23];
  assign n103 = a[26];
  assign n115 = a[29];

  HS65_LH_NOR3AX2 U1941 ( .A(n2758), .B(n2754), .C(n2753), .Z(n2723) );
  HS65_LH_NOR3AX2 U1942 ( .A(n3058), .B(n3054), .C(n3053), .Z(n3023) );
  HS65_LH_NOR3AX2 U1943 ( .A(n3101), .B(n3097), .C(n3096), .Z(n3066) );
  HS65_LH_NOR3AX2 U1944 ( .A(n2929), .B(n2925), .C(n2924), .Z(n2894) );
  HS65_LH_NOR3AX2 U1945 ( .A(n2801), .B(n2797), .C(n2796), .Z(n2766) );
  HS65_LH_NOR3AX2 U1946 ( .A(n2843), .B(n2839), .C(n2838), .Z(n2808) );
  HS65_LH_NOR3AX2 U1947 ( .A(n2886), .B(n2882), .C(n2881), .Z(n2851) );
  HS65_LH_NOR3AX2 U1948 ( .A(n2972), .B(n2968), .C(n2967), .Z(n2937) );
  HS65_LH_NOR3AX2 U1949 ( .A(n3015), .B(n3011), .C(n3010), .Z(n2980) );
  HS65_LH_AND2X4 U1950 ( .A(n2753), .B(n2754), .Z(n2718) );
  HS65_LH_AND2X4 U1951 ( .A(n3010), .B(n3011), .Z(n2975) );
  HS65_LH_AND2X4 U1952 ( .A(n2796), .B(n2797), .Z(n2761) );
  HS65_LH_AND2X4 U1953 ( .A(n2838), .B(n2839), .Z(n2417) );
  HS65_LH_AND2X4 U1954 ( .A(n2881), .B(n2882), .Z(n2846) );
  HS65_LH_AND2X4 U1955 ( .A(n2924), .B(n2925), .Z(n2889) );
  HS65_LH_AND2X4 U1956 ( .A(n2967), .B(n2968), .Z(n2932) );
  HS65_LH_AND2X4 U1957 ( .A(n3053), .B(n3054), .Z(n3018) );
  HS65_LH_AND2X4 U1958 ( .A(n3096), .B(n3097), .Z(n3061) );
  HS65_LH_NOR3AX2 U1959 ( .A(a[31]), .B(n3104), .C(n3103), .Z(n2670) );
  HS65_LH_NOR3AX2 U1960 ( .A(n2711), .B(a[0]), .C(a[1]), .Z(n2681) );
  HS65_LH_IVX9 U1961 ( .A(n1007), .Z(n4719) );
  HS65_LH_FA1X4 U1962 ( .A0(n530), .B0(n546), .CI(n253), .CO(n252), .S0(
        product[37]) );
  HS65_LH_FA1X4 U1963 ( .A0(n480), .B0(n494), .CI(n250), .CO(n249), .S0(
        product[40]) );
  HS65_LH_FA1X4 U1964 ( .A0(n435), .B0(n448), .CI(n247), .CO(n246), .S0(
        product[43]) );
  HS65_LH_FA1X4 U1965 ( .A0(n397), .B0(n407), .CI(n244), .CO(n243), .S0(
        product[46]) );
  HS65_LH_FA1X4 U1966 ( .A0(n364), .B0(n373), .CI(n241), .CO(n240), .S0(
        product[49]) );
  HS65_LH_FA1X4 U1967 ( .A0(n338), .B0(n344), .CI(n238), .CO(n237), .S0(
        product[52]) );
  HS65_LH_FA1X4 U1968 ( .A0(n317), .B0(n322), .CI(n235), .CO(n234), .S0(
        product[55]) );
  HS65_LH_FA1X4 U1969 ( .A0(n303), .B0(n305), .CI(n232), .CO(n231), .S0(
        product[58]) );
  HS65_LH_HA1X4 U1970 ( .A0(n4678), .B0(n975), .CO(n1006), .S0(n1007) );
  HS65_LH_OAI22X6 U1971 ( .A(n4676), .B(n2757), .C(n4580), .D(n2757), .Z(n2756) );
  HS65_LH_AND2X4 U1972 ( .A(n4585), .B(n4679), .Z(n2757) );
  HS65_LH_OAI22X6 U1973 ( .A(n4676), .B(n3100), .C(n4495), .D(n3100), .Z(n3099) );
  HS65_LH_AND2X4 U1974 ( .A(n4500), .B(n4679), .Z(n3100) );
  HS65_LH_FA1X4 U1975 ( .A0(n1351), .B0(n1319), .CI(n549), .CO(n546), .S0(n547) );
  HS65_LHS_XOR2X6 U1976 ( .A(n4684), .B(n2759), .Z(n1351) );
  HS65_LHS_XOR2X6 U1977 ( .A(n31), .B(n2794), .Z(n1319) );
  HS65_LH_AOI22X6 U1978 ( .A(n4586), .B(n1006), .C(n4580), .D(n4678), .Z(n2759) );
  HS65_LH_FA1X4 U1979 ( .A0(n1281), .B0(n1249), .CI(n451), .CO(n448), .S0(n449) );
  HS65_LHS_XOR2X6 U1980 ( .A(n4690), .B(n2844), .Z(n1281) );
  HS65_LHS_XOR2X6 U1981 ( .A(n55), .B(n2879), .Z(n1249) );
  HS65_LH_AOI22X6 U1982 ( .A(n4567), .B(n1006), .C(n4561), .D(n4678), .Z(n2844) );
  HS65_LH_FA1X4 U1983 ( .A0(n1141), .B0(n1109), .CI(n325), .CO(n322), .S0(n323) );
  HS65_LHS_XOR2X6 U1984 ( .A(n4702), .B(n3016), .Z(n1141) );
  HS65_LHS_XOR2X6 U1985 ( .A(n4703), .B(n3051), .Z(n1109) );
  HS65_LH_AOI22X6 U1986 ( .A(n4523), .B(n1006), .C(n4517), .D(n4678), .Z(n3016) );
  HS65_LH_FA1X4 U1987 ( .A0(n1106), .B0(n1074), .CI(n308), .CO(n305), .S0(n306) );
  HS65_LHS_XOR2X6 U1988 ( .A(n4705), .B(n3059), .Z(n1106) );
  HS65_LHS_XOR2X6 U1989 ( .A(n4707), .B(n3094), .Z(n1074) );
  HS65_LH_AOI22X6 U1990 ( .A(n4512), .B(n1006), .C(n4506), .D(n4678), .Z(n3059) );
  HS65_LH_FA1X4 U1991 ( .A0(n1318), .B0(n532), .CI(n548), .CO(n529), .S0(n530)
         );
  HS65_LHS_XOR2X6 U1992 ( .A(n31), .B(n2795), .Z(n1318) );
  HS65_LH_MX41X7 U1993 ( .D0(n2762), .S0(n1008), .D1(n4570), .S1(n4675), .D2(
        n4574), .S2(n4677), .D3(n4579), .S3(n4678), .Z(n2795) );
  HS65_LH_FA1X4 U1994 ( .A0(n1316), .B0(n1284), .CI(n497), .CO(n494), .S0(n495) );
  HS65_LHS_XOR2X6 U1995 ( .A(n4687), .B(n2802), .Z(n1316) );
  HS65_LHS_XOR2X6 U1996 ( .A(n4689), .B(n2836), .Z(n1284) );
  HS65_LH_AOI22X6 U1997 ( .A(n4575), .B(n1006), .C(n4569), .D(n4678), .Z(n2802) );
  HS65_LH_FA1X4 U1998 ( .A0(n1283), .B0(n482), .CI(n496), .CO(n479), .S0(n480)
         );
  HS65_LHS_XOR2X6 U1999 ( .A(n43), .B(n2837), .Z(n1283) );
  HS65_LH_MX41X7 U2000 ( .D0(n2804), .S0(n1008), .D1(n4566), .S1(n4677), .D2(
        n4611), .S2(n4679), .D3(n4562), .S3(n4674), .Z(n2837) );
  HS65_LH_FA1X4 U2001 ( .A0(n1248), .B0(n437), .CI(n450), .CO(n434), .S0(n435)
         );
  HS65_LHS_XOR2X6 U2002 ( .A(n55), .B(n2880), .Z(n1248) );
  HS65_LH_MX41X7 U2003 ( .D0(n2847), .S0(n1008), .D1(n4551), .S1(n4675), .D2(
        n4555), .S2(n4677), .D3(n4560), .S3(n4678), .Z(n2880) );
  HS65_LH_FA1X4 U2004 ( .A0(n1246), .B0(n1214), .CI(n410), .CO(n407), .S0(n408) );
  HS65_LHS_XOR2X6 U2005 ( .A(n4693), .B(n2887), .Z(n1246) );
  HS65_LHS_XOR2X6 U2006 ( .A(n4694), .B(n2922), .Z(n1214) );
  HS65_LH_AOI22X6 U2007 ( .A(n4556), .B(n1006), .C(n4550), .D(n4678), .Z(n2887) );
  HS65_LH_FA1X4 U2008 ( .A0(n1213), .B0(n399), .CI(n409), .CO(n396), .S0(n397)
         );
  HS65_LHS_XOR2X6 U2009 ( .A(n67), .B(n2923), .Z(n1213) );
  HS65_LH_MX41X7 U2010 ( .D0(n2890), .S0(n1008), .D1(n4540), .S1(n4675), .D2(
        n4544), .S2(n4677), .D3(n4549), .S3(n4678), .Z(n2923) );
  HS65_LH_FA1X4 U2011 ( .A0(n1211), .B0(n1179), .CI(n376), .CO(n373), .S0(n374) );
  HS65_LHS_XOR2X6 U2012 ( .A(n4696), .B(n2930), .Z(n1211) );
  HS65_LHS_XOR2X6 U2013 ( .A(n4698), .B(n2965), .Z(n1179) );
  HS65_LH_AOI22X6 U2014 ( .A(n4545), .B(n1006), .C(n4539), .D(n4678), .Z(n2930) );
  HS65_LH_FA1X4 U2015 ( .A0(n1178), .B0(n366), .CI(n375), .CO(n363), .S0(n364)
         );
  HS65_LHS_XOR2X6 U2016 ( .A(n79), .B(n2966), .Z(n1178) );
  HS65_LH_MX41X7 U2017 ( .D0(n2933), .S0(n1008), .D1(n4529), .S1(n4675), .D2(
        n4533), .S2(n4677), .D3(n4538), .S3(n4678), .Z(n2966) );
  HS65_LH_FA1X4 U2018 ( .A0(n1176), .B0(n1144), .CI(n347), .CO(n344), .S0(n345) );
  HS65_LHS_XOR2X6 U2019 ( .A(n4699), .B(n2973), .Z(n1176) );
  HS65_LHS_XOR2X6 U2020 ( .A(n4701), .B(n3008), .Z(n1144) );
  HS65_LH_AOI22X6 U2021 ( .A(n4534), .B(n1006), .C(n4528), .D(n4678), .Z(n2973) );
  HS65_LH_FA1X4 U2022 ( .A0(n1143), .B0(n340), .CI(n346), .CO(n337), .S0(n338)
         );
  HS65_LHS_XOR2X6 U2023 ( .A(n91), .B(n3009), .Z(n1143) );
  HS65_LH_MX41X7 U2024 ( .D0(n2976), .S0(n1008), .D1(n4527), .S1(n4679), .D2(
        n4518), .S2(n4675), .D3(n4522), .S3(n4677), .Z(n3009) );
  HS65_LH_FA1X4 U2025 ( .A0(n1108), .B0(n319), .CI(n324), .CO(n316), .S0(n317)
         );
  HS65_LHS_XOR2X6 U2026 ( .A(n103), .B(n3052), .Z(n1108) );
  HS65_LH_MX41X7 U2027 ( .D0(n3019), .S0(n1008), .D1(n4507), .S1(n4674), .D2(
        n4511), .S2(n4677), .D3(n4516), .S3(n4679), .Z(n3052) );
  HS65_LH_FA1X4 U2028 ( .A0(n1073), .B0(n304), .CI(n307), .CO(n302), .S0(n303)
         );
  HS65_LHS_XOR2X6 U2029 ( .A(n115), .B(n3095), .Z(n1073) );
  HS65_LH_MX41X7 U2030 ( .D0(n3062), .S0(n1008), .D1(n4495), .S1(n4674), .D2(
        n4500), .S2(n4677), .D3(n4505), .S3(n4679), .Z(n3095) );
  HS65_LH_FA1X4 U2031 ( .A0(n585), .B0(n602), .CI(n1353), .CO(n582), .S0(n583)
         );
  HS65_LHS_XOR2X6 U2032 ( .A(n19), .B(n2752), .Z(n1353) );
  HS65_LH_MX41X7 U2033 ( .D0(n2719), .S0(n1008), .D1(n4581), .S1(n4675), .D2(
        n4585), .S2(n4677), .D3(n4590), .S3(n4678), .Z(n2752) );
  HS65_LH_HA1X4 U2034 ( .A0(n31), .B0(n1349), .CO(n934), .S0(n935) );
  HS65_LHS_XOR2X6 U2035 ( .A(n31), .B(n2760), .Z(n1349) );
  HS65_LH_AO22X9 U2036 ( .A(n4616), .B(n4579), .C(n4615), .D(n2762), .Z(n2760)
         );
  HS65_LH_HA1X4 U2037 ( .A0(n19), .B0(n1384), .CO(n940), .S0(n941) );
  HS65_LHS_XOR2X6 U2038 ( .A(n19), .B(n2717), .Z(n1384) );
  HS65_LH_AO22X9 U2039 ( .A(n4616), .B(n4590), .C(n4615), .D(n2719), .Z(n2717)
         );
  HS65_LH_HA1X4 U2040 ( .A0(n43), .B0(n1314), .CO(n922), .S0(n923) );
  HS65_LHS_XOR2X6 U2041 ( .A(n43), .B(n2803), .Z(n1314) );
  HS65_LH_AO22X9 U2042 ( .A(n4616), .B(n4613), .C(n4615), .D(n2804), .Z(n2803)
         );
  HS65_LH_HA1X4 U2043 ( .A0(n55), .B0(n1279), .CO(n904), .S0(n905) );
  HS65_LHS_XOR2X6 U2044 ( .A(n55), .B(n2845), .Z(n1279) );
  HS65_LH_AO22X9 U2045 ( .A(n4615), .B(n4560), .C(n4615), .D(n2847), .Z(n2845)
         );
  HS65_LH_HA1X4 U2046 ( .A0(n67), .B0(n1244), .CO(n880), .S0(n881) );
  HS65_LHS_XOR2X6 U2047 ( .A(n67), .B(n2888), .Z(n1244) );
  HS65_LH_AO22X9 U2048 ( .A(n4616), .B(n4549), .C(n4615), .D(n2890), .Z(n2888)
         );
  HS65_LH_HA1X4 U2049 ( .A0(n79), .B0(n1209), .CO(n850), .S0(n851) );
  HS65_LHS_XOR2X6 U2050 ( .A(n79), .B(n2931), .Z(n1209) );
  HS65_LH_AO22X9 U2051 ( .A(n4616), .B(n4538), .C(n4615), .D(n2933), .Z(n2931)
         );
  HS65_LH_HA1X4 U2052 ( .A0(n4700), .B0(n1174), .CO(n814), .S0(n815) );
  HS65_LHS_XOR2X6 U2053 ( .A(n91), .B(n2974), .Z(n1174) );
  HS65_LH_AO22X9 U2054 ( .A(n4616), .B(n4527), .C(n4615), .D(n2976), .Z(n2974)
         );
  HS65_LH_HA1X4 U2055 ( .A0(n4703), .B0(n1139), .CO(n772), .S0(n773) );
  HS65_LHS_XOR2X6 U2056 ( .A(n103), .B(n3017), .Z(n1139) );
  HS65_LH_AO22X9 U2057 ( .A(n4616), .B(n4516), .C(n4615), .D(n3019), .Z(n3017)
         );
  HS65_LH_HA1X4 U2058 ( .A0(n115), .B0(n1104), .CO(n724), .S0(n725) );
  HS65_LHS_XOR2X6 U2059 ( .A(n115), .B(n3060), .Z(n1104) );
  HS65_LH_AO22X9 U2060 ( .A(n4616), .B(n4505), .C(n4615), .D(n3062), .Z(n3060)
         );
  HS65_LH_HA1X4 U2061 ( .A0(n1383), .B0(n940), .CO(n938), .S0(n939) );
  HS65_LHS_XOR2X6 U2062 ( .A(n19), .B(n2720), .Z(n1383) );
  HS65_LH_AO222X4 U2063 ( .A(n4619), .B(n4590), .C(n4615), .D(n4585), .E(n1038), .F(n2719), .Z(n2720) );
  HS65_LH_HA1X4 U2064 ( .A0(n1348), .B0(n934), .CO(n930), .S0(n931) );
  HS65_LHS_XOR2X6 U2065 ( .A(n4685), .B(n2763), .Z(n1348) );
  HS65_LH_AO222X4 U2066 ( .A(n4619), .B(n4579), .C(n4615), .D(n4574), .E(n1038), .F(n2762), .Z(n2763) );
  HS65_LH_HA1X4 U2067 ( .A0(n1313), .B0(n922), .CO(n916), .S0(n917) );
  HS65_LHS_XOR2X6 U2068 ( .A(n4688), .B(n2805), .Z(n1313) );
  HS65_LH_AO222X4 U2069 ( .A(n4619), .B(n4613), .C(n4615), .D(n4566), .E(n1038), .F(n2804), .Z(n2805) );
  HS65_LH_HA1X4 U2070 ( .A0(n1278), .B0(n904), .CO(n896), .S0(n897) );
  HS65_LHS_XOR2X6 U2071 ( .A(n4691), .B(n2848), .Z(n1278) );
  HS65_LH_AO222X4 U2072 ( .A(n4619), .B(n4560), .C(n4615), .D(n4555), .E(n1038), .F(n2847), .Z(n2848) );
  HS65_LH_HA1X4 U2073 ( .A0(n1243), .B0(n880), .CO(n870), .S0(n871) );
  HS65_LHS_XOR2X6 U2074 ( .A(n4694), .B(n2891), .Z(n1243) );
  HS65_LH_AO222X4 U2075 ( .A(n4619), .B(n4549), .C(n4615), .D(n4544), .E(n1038), .F(n2890), .Z(n2891) );
  HS65_LH_HA1X4 U2076 ( .A0(n1208), .B0(n850), .CO(n838), .S0(n839) );
  HS65_LHS_XOR2X6 U2077 ( .A(n4697), .B(n2934), .Z(n1208) );
  HS65_LH_AO222X4 U2078 ( .A(n4619), .B(n4538), .C(n4615), .D(n4533), .E(n1038), .F(n2933), .Z(n2934) );
  HS65_LH_HA1X4 U2079 ( .A0(n1173), .B0(n814), .CO(n800), .S0(n801) );
  HS65_LHS_XOR2X6 U2080 ( .A(n4700), .B(n2977), .Z(n1173) );
  HS65_LH_AO222X4 U2081 ( .A(n4619), .B(n4527), .C(n4615), .D(n4522), .E(n1038), .F(n2976), .Z(n2977) );
  HS65_LH_HA1X4 U2082 ( .A0(n1138), .B0(n772), .CO(n756), .S0(n757) );
  HS65_LHS_XOR2X6 U2083 ( .A(n4703), .B(n3020), .Z(n1138) );
  HS65_LH_AO222X4 U2084 ( .A(n4619), .B(n4516), .C(n4615), .D(n4511), .E(n1038), .F(n3019), .Z(n3020) );
  HS65_LH_HA1X4 U2085 ( .A0(n1103), .B0(n724), .CO(n706), .S0(n707) );
  HS65_LHS_XOR2X6 U2086 ( .A(n4706), .B(n3063), .Z(n1103) );
  HS65_LH_AO222X4 U2087 ( .A(n4619), .B(n4505), .C(n4615), .D(n4500), .E(n1038), .F(n3062), .Z(n3063) );
  HS65_LH_HA1X4 U2088 ( .A0(n1382), .B0(n938), .CO(n936), .S0(n937) );
  HS65_LHS_XOR2X6 U2089 ( .A(n19), .B(n2722), .Z(n1382) );
  HS65_LH_MX41X7 U2090 ( .D0(n2719), .S0(n1037), .D1(n4581), .S1(n4616), .D2(
        n4585), .S2(n4618), .D3(n4590), .S3(n4620), .Z(n2722) );
  HS65_LH_HA1X4 U2091 ( .A0(n1347), .B0(n930), .CO(n926), .S0(n927) );
  HS65_LHS_XOR2X6 U2092 ( .A(n31), .B(n2765), .Z(n1347) );
  HS65_LH_MX41X7 U2093 ( .D0(n2762), .S0(n1037), .D1(n4570), .S1(n4616), .D2(
        n4574), .S2(n4618), .D3(n4579), .S3(n4620), .Z(n2765) );
  HS65_LH_HA1X4 U2094 ( .A0(n1312), .B0(n916), .CO(n910), .S0(n911) );
  HS65_LHS_XOR2X6 U2095 ( .A(n43), .B(n2807), .Z(n1312) );
  HS65_LH_MX41X7 U2096 ( .D0(n2804), .S0(n1037), .D1(n4613), .S1(n4620), .D2(
        n4565), .S2(n4618), .D3(n4562), .S3(n4616), .Z(n2807) );
  HS65_LH_HA1X4 U2097 ( .A0(n1277), .B0(n896), .CO(n888), .S0(n889) );
  HS65_LHS_XOR2X6 U2098 ( .A(n55), .B(n2850), .Z(n1277) );
  HS65_LH_MX41X7 U2099 ( .D0(n2847), .S0(n1037), .D1(n4551), .S1(n4616), .D2(
        n4555), .S2(n4618), .D3(n4560), .S3(n4620), .Z(n2850) );
  HS65_LH_HA1X4 U2100 ( .A0(n1242), .B0(n870), .CO(n860), .S0(n861) );
  HS65_LHS_XOR2X6 U2101 ( .A(n67), .B(n2893), .Z(n1242) );
  HS65_LH_MX41X7 U2102 ( .D0(n2890), .S0(n1037), .D1(n4540), .S1(n4616), .D2(
        n4544), .S2(n4618), .D3(n4549), .S3(n4620), .Z(n2893) );
  HS65_LH_HA1X4 U2103 ( .A0(n1207), .B0(n838), .CO(n826), .S0(n827) );
  HS65_LHS_XOR2X6 U2104 ( .A(n79), .B(n2936), .Z(n1207) );
  HS65_LH_MX41X7 U2105 ( .D0(n2933), .S0(n1037), .D1(n4529), .S1(n4616), .D2(
        n4533), .S2(n4619), .D3(n4538), .S3(n4620), .Z(n2936) );
  HS65_LH_HA1X4 U2106 ( .A0(n1172), .B0(n800), .CO(n786), .S0(n787) );
  HS65_LHS_XOR2X6 U2107 ( .A(n91), .B(n2979), .Z(n1172) );
  HS65_LH_MX41X7 U2108 ( .D0(n2976), .S0(n1037), .D1(n4527), .S1(n4620), .D2(
        n4518), .S2(n4617), .D3(n4522), .S3(n4618), .Z(n2979) );
  HS65_LH_HA1X4 U2109 ( .A0(n1137), .B0(n756), .CO(n740), .S0(n741) );
  HS65_LHS_XOR2X6 U2110 ( .A(n103), .B(n3022), .Z(n1137) );
  HS65_LH_MX41X7 U2111 ( .D0(n3019), .S0(n1037), .D1(n4507), .S1(n4616), .D2(
        n4511), .S2(n4619), .D3(n4516), .S3(n4620), .Z(n3022) );
  HS65_LH_HA1X4 U2112 ( .A0(n1102), .B0(n706), .CO(n688), .S0(n689) );
  HS65_LHS_XOR2X6 U2113 ( .A(n115), .B(n3065), .Z(n1102) );
  HS65_LH_MX41X7 U2114 ( .D0(n3062), .S0(n1037), .D1(n4496), .S1(n4616), .D2(
        n4500), .S2(n4618), .D3(n4505), .S3(n4620), .Z(n3065) );
  HS65_LH_FA1X4 U2115 ( .A0(n1381), .B0(n935), .CI(n936), .CO(n932), .S0(n933)
         );
  HS65_LHS_XOR2X6 U2116 ( .A(n19), .B(n2724), .Z(n1381) );
  HS65_LH_MX41X7 U2117 ( .D0(n2719), .S0(n1036), .D1(n4581), .S1(n4618), .D2(
        n4585), .S2(n4621), .D3(n4590), .S3(n4622), .Z(n2724) );
  HS65_LH_FA1X4 U2118 ( .A0(n1346), .B0(n923), .CI(n926), .CO(n920), .S0(n921)
         );
  HS65_LHS_XOR2X6 U2119 ( .A(n31), .B(n2767), .Z(n1346) );
  HS65_LH_MX41X7 U2120 ( .D0(n2762), .S0(n1036), .D1(n4570), .S1(n4618), .D2(
        n4574), .S2(n4621), .D3(n4579), .S3(n4622), .Z(n2767) );
  HS65_LH_FA1X4 U2121 ( .A0(n1276), .B0(n881), .CI(n888), .CO(n878), .S0(n879)
         );
  HS65_LHS_XOR2X6 U2122 ( .A(n55), .B(n2852), .Z(n1276) );
  HS65_LH_MX41X7 U2123 ( .D0(n2847), .S0(n1036), .D1(n4551), .S1(n4618), .D2(
        n4555), .S2(n4621), .D3(n4560), .S3(n4622), .Z(n2852) );
  HS65_LH_FA1X4 U2124 ( .A0(n1241), .B0(n851), .CI(n860), .CO(n848), .S0(n849)
         );
  HS65_LHS_XOR2X6 U2125 ( .A(n67), .B(n2895), .Z(n1241) );
  HS65_LH_MX41X7 U2126 ( .D0(n2890), .S0(n1036), .D1(n4540), .S1(n4618), .D2(
        n4544), .S2(n4621), .D3(n4549), .S3(n4622), .Z(n2895) );
  HS65_LH_FA1X4 U2127 ( .A0(n1206), .B0(n815), .CI(n826), .CO(n812), .S0(n813)
         );
  HS65_LHS_XOR2X6 U2128 ( .A(n79), .B(n2938), .Z(n1206) );
  HS65_LH_MX41X7 U2129 ( .D0(n2933), .S0(n1036), .D1(n4529), .S1(n4618), .D2(
        n4532), .S2(n4621), .D3(n4538), .S3(n4622), .Z(n2938) );
  HS65_LH_FA1X4 U2130 ( .A0(n1171), .B0(n773), .CI(n786), .CO(n770), .S0(n771)
         );
  HS65_LHS_XOR2X6 U2131 ( .A(n91), .B(n2981), .Z(n1171) );
  HS65_LH_MX41X7 U2132 ( .D0(n2976), .S0(n1036), .D1(n4527), .S1(n4622), .D2(
        n4518), .S2(n4619), .D3(n4522), .S3(n4620), .Z(n2981) );
  HS65_LH_FA1X4 U2133 ( .A0(n1136), .B0(n725), .CI(n740), .CO(n722), .S0(n723)
         );
  HS65_LHS_XOR2X6 U2134 ( .A(n103), .B(n3024), .Z(n1136) );
  HS65_LH_MX41X7 U2135 ( .D0(n3019), .S0(n1036), .D1(n4507), .S1(n4618), .D2(
        n4510), .S2(n4621), .D3(n4516), .S3(n4622), .Z(n3024) );
  HS65_LH_FA1X4 U2136 ( .A0(n1311), .B0(n905), .CI(n910), .CO(n902), .S0(n903)
         );
  HS65_LHS_XOR2X6 U2137 ( .A(n43), .B(n2809), .Z(n1311) );
  HS65_LH_MX41X7 U2138 ( .D0(n2804), .S0(n1036), .D1(n4613), .S1(n4623), .D2(
        n4565), .S2(n4621), .D3(n4562), .S3(n4618), .Z(n2809) );
  HS65_LH_FA1X4 U2139 ( .A0(n507), .B0(n524), .CI(n522), .CO(n504), .S0(n505)
         );
  HS65_LH_FA1X4 U2140 ( .A0(n583), .B0(n600), .CI(n256), .CO(n255), .S0(
        product[34]) );
  HS65_LH_FA1X4 U2141 ( .A0(n565), .B0(n582), .CI(n255), .CO(n254), .S0(
        product[35]) );
  HS65_LH_FA1X4 U2142 ( .A0(n503), .B0(n520), .CI(n518), .CO(n500), .S0(n501)
         );
  HS65_LH_FA1X4 U2143 ( .A0(n513), .B0(n529), .CI(n252), .CO(n251), .S0(
        product[38]) );
  HS65_LH_FA1X4 U2144 ( .A0(n457), .B0(n472), .CI(n470), .CO(n454), .S0(n455)
         );
  HS65_LH_FA1X4 U2145 ( .A0(n465), .B0(n479), .CI(n249), .CO(n248), .S0(
        product[41]) );
  HS65_LH_FA1X4 U2146 ( .A0(n416), .B0(n429), .CI(n427), .CO(n413), .S0(n414)
         );
  HS65_LH_FA1X4 U2147 ( .A0(n577), .B0(n594), .CI(n592), .CO(n574), .S0(n575)
         );
  HS65_LH_FA1X4 U2148 ( .A0(n559), .B0(n576), .CI(n574), .CO(n556), .S0(n557)
         );
  HS65_LH_FA1X4 U2149 ( .A0(n573), .B0(n590), .CI(n588), .CO(n570), .S0(n571)
         );
  HS65_LH_FA1X4 U2150 ( .A0(n547), .B0(n564), .CI(n254), .CO(n253), .S0(
        product[36]) );
  HS65_LH_FA1X4 U2151 ( .A0(n461), .B0(n476), .CI(n474), .CO(n458), .S0(n459)
         );
  HS65_LH_FA1X4 U2152 ( .A0(n499), .B0(n516), .CI(n514), .CO(n496), .S0(n497)
         );
  HS65_LH_FA1X4 U2153 ( .A0(n495), .B0(n512), .CI(n251), .CO(n250), .S0(
        product[39]) );
  HS65_LH_FA1X4 U2154 ( .A0(n453), .B0(n468), .CI(n466), .CO(n450), .S0(n451)
         );
  HS65_LH_FA1X4 U2155 ( .A0(n449), .B0(n464), .CI(n248), .CO(n247), .S0(
        product[42]) );
  HS65_LH_FA1X4 U2156 ( .A0(n412), .B0(n425), .CI(n423), .CO(n409), .S0(n410)
         );
  HS65_LH_FA1X4 U2157 ( .A0(n422), .B0(n434), .CI(n246), .CO(n245), .S0(
        product[44]) );
  HS65_LH_FA1X4 U2158 ( .A0(n382), .B0(n393), .CI(n391), .CO(n379), .S0(n380)
         );
  HS65_LH_FA1X4 U2159 ( .A0(n408), .B0(n421), .CI(n245), .CO(n244), .S0(
        product[45]) );
  HS65_LH_FA1X4 U2160 ( .A0(n378), .B0(n389), .CI(n387), .CO(n375), .S0(n376)
         );
  HS65_LH_FA1X4 U2161 ( .A0(n386), .B0(n396), .CI(n243), .CO(n242), .S0(
        product[47]) );
  HS65_LH_FA1X4 U2162 ( .A0(n374), .B0(n385), .CI(n242), .CO(n241), .S0(
        product[48]) );
  HS65_LH_FA1X4 U2163 ( .A0(n349), .B0(n358), .CI(n356), .CO(n346), .S0(n347)
         );
  HS65_LH_FA1X4 U2164 ( .A0(n355), .B0(n363), .CI(n240), .CO(n239), .S0(
        product[50]) );
  HS65_LH_FA1X4 U2165 ( .A0(n345), .B0(n354), .CI(n239), .CO(n238), .S0(
        product[51]) );
  HS65_LH_FA1X4 U2166 ( .A0(n327), .B0(n334), .CI(n332), .CO(n324), .S0(n325)
         );
  HS65_LH_FA1X4 U2167 ( .A0(n331), .B0(n337), .CI(n237), .CO(n236), .S0(
        product[53]) );
  HS65_LH_FA1X4 U2168 ( .A0(n312), .B0(n316), .CI(n234), .CO(n233), .S0(
        product[56]) );
  HS65_LH_FA1X4 U2169 ( .A0(n296), .B0(n299), .CI(n230), .CO(n229), .S0(
        product[60]) );
  HS65_LH_FA1X4 U2170 ( .A0(n555), .B0(n572), .CI(n570), .CO(n552), .S0(n553)
         );
  HS65_LH_FA1X4 U2171 ( .A0(n323), .B0(n330), .CI(n236), .CO(n235), .S0(
        product[54]) );
  HS65_LH_FA1X4 U2172 ( .A0(n306), .B0(n311), .CI(n233), .CO(n232), .S0(
        product[57]) );
  HS65_LH_FA1X4 U2173 ( .A0(n300), .B0(n302), .CI(n231), .CO(n230), .S0(
        product[59]) );
  HS65_LH_FA1X4 U2174 ( .A0(n295), .B0(n294), .CI(n229), .CO(n228), .S0(
        product[61]) );
  HS65_LH_FA1X4 U2175 ( .A0(n4618), .B0(n4620), .CI(n1005), .CO(n1004), .S0(
        n1037) );
  HS65_LH_FA1X4 U2176 ( .A0(n4620), .B0(n4622), .CI(n1004), .CO(n1003), .S0(
        n1036) );
  HS65_LH_FA1X4 U2177 ( .A0(n4660), .B0(n4662), .CI(n984), .CO(n983), .S0(
        n1016) );
  HS65_LH_FA1X4 U2178 ( .A0(n4674), .B0(n4676), .CI(n977), .CO(n976), .S0(
        n1009) );
  HS65_LH_IVX9 U2179 ( .A(n462), .Z(n4710) );
  HS65_LH_IVX9 U2180 ( .A(n383), .Z(n4711) );
  HS65_LH_IVX9 U2181 ( .A(n328), .Z(n4712) );
  HS65_LH_IVX9 U2182 ( .A(n297), .Z(n4716) );
  HS65_LH_IVX9 U2183 ( .A(n510), .Z(n4709) );
  HS65_LH_IVX9 U2184 ( .A(n419), .Z(n4713) );
  HS65_LH_IVX9 U2185 ( .A(n352), .Z(n4714) );
  HS65_LH_IVX9 U2186 ( .A(n309), .Z(n4715) );
  HS65_LH_FA1X4 U2187 ( .A0(n4676), .B0(n4678), .CI(n976), .CO(n975), .S0(
        n1008) );
  HS65_LH_AND2X4 U2188 ( .A(n4574), .B(n4679), .Z(n2800) );
  HS65_LH_AND2X4 U2189 ( .A(n4566), .B(n4679), .Z(n2842) );
  HS65_LH_AND2X4 U2190 ( .A(n4555), .B(n4679), .Z(n2885) );
  HS65_LH_AND2X4 U2191 ( .A(n4544), .B(n4679), .Z(n2928) );
  HS65_LH_AND2X4 U2192 ( .A(n4533), .B(n4679), .Z(n2971) );
  HS65_LH_AND2X4 U2193 ( .A(n4520), .B(n4679), .Z(n3014) );
  HS65_LH_AND2X4 U2194 ( .A(n4511), .B(n4679), .Z(n3057) );
  HS65_LH_BFX9 U2195 ( .A(n4614), .Z(n4615) );
  HS65_LH_BFX9 U2196 ( .A(n4614), .Z(n4616) );
  HS65_LH_HA1X4 U2197 ( .A0(n4618), .B0(n4615), .CO(n1005), .S0(n1038) );
  HS65_LH_BFX9 U2198 ( .A(n4614), .Z(n4617) );
  HS65_LH_FA1X4 U2199 ( .A0(n510), .B0(n4687), .CI(n1059), .CO(n462), .S0(n493) );
  HS65_LH_MX41X7 U2200 ( .D0(n1029), .S0(n4491), .D1(n4636), .S1(n4607), .D2(
        n4634), .S2(n4603), .D3(n4632), .S3(n4609), .Z(n1059) );
  HS65_LH_FA1X4 U2201 ( .A0(n4684), .B0(n4682), .CI(n1062), .CO(n510), .S0(
        n545) );
  HS65_LH_MX41X7 U2202 ( .D0(n1032), .S0(n4492), .D1(n4630), .S1(n4607), .D2(
        n4628), .S2(n4603), .D3(n4626), .S3(n4609), .Z(n1062) );
  HS65_LH_FA1X4 U2203 ( .A0(n419), .B0(n4693), .CI(n1054), .CO(n383), .S0(n406) );
  HS65_LH_MX41X7 U2204 ( .D0(n1023), .S0(n4491), .D1(n4644), .S1(n4610), .D2(
        n4646), .S2(n4603), .D3(n4648), .S3(n4607), .Z(n1054) );
  HS65_LH_FA1X4 U2205 ( .A0(n352), .B0(n4699), .CI(n1049), .CO(n328), .S0(n343) );
  HS65_LH_MX41X7 U2206 ( .D0(n1017), .S0(n4491), .D1(n4656), .S1(n4610), .D2(
        n4658), .S2(n4603), .D3(n4660), .S3(n4607), .Z(n1049) );
  HS65_LH_FA1X4 U2207 ( .A0(n309), .B0(n4705), .CI(n1044), .CO(n297), .S0(n304) );
  HS65_LH_MX41X7 U2208 ( .D0(n1011), .S0(n4490), .D1(n4668), .S1(n4609), .D2(
        n4670), .S2(n4603), .D3(n4672), .S3(n4607), .Z(n1044) );
  HS65_LH_FA1X4 U2209 ( .A0(n462), .B0(n4690), .CI(n1056), .CO(n446), .S0(n447) );
  HS65_LH_MX41X7 U2210 ( .D0(n1026), .S0(n4490), .D1(n4606), .S1(n4642), .D2(
        n4640), .S2(n4602), .D3(n4638), .S3(n4609), .Z(n1056) );
  HS65_LH_FA1X4 U2211 ( .A0(n383), .B0(n4696), .CI(n1051), .CO(n371), .S0(n372) );
  HS65_LH_MX41X7 U2212 ( .D0(n1020), .S0(n4491), .D1(n4650), .S1(n4610), .D2(
        n4652), .S2(n4603), .D3(n4654), .S3(n4607), .Z(n1051) );
  HS65_LH_FA1X4 U2213 ( .A0(n328), .B0(n4702), .CI(n1046), .CO(n320), .S0(n321) );
  HS65_LH_MX41X7 U2214 ( .D0(n1014), .S0(n4490), .D1(n4662), .S1(n4609), .D2(
        n4664), .S2(n4602), .D3(n4666), .S3(n4606), .Z(n1046) );
  HS65_LH_FA1X4 U2215 ( .A0(n1194), .B0(n613), .CI(n628), .CO(n610), .S0(n611)
         );
  HS65_LHS_XOR2X6 U2216 ( .A(n4697), .B(n2950), .Z(n1194) );
  HS65_LH_MX41X7 U2217 ( .D0(n4534), .S0(n1024), .D1(n4528), .S1(n4642), .D2(
        n4531), .S2(n4645), .D3(n4536), .S3(n4646), .Z(n2950) );
  HS65_LH_FA1X4 U2218 ( .A0(n1226), .B0(n611), .CI(n626), .CO(n608), .S0(n609)
         );
  HS65_LHS_XOR2X6 U2219 ( .A(n4695), .B(n2910), .Z(n1226) );
  HS65_LH_MX41X7 U2220 ( .D0(n2890), .S0(n1021), .D1(n4540), .S1(n4649), .D2(
        n4543), .S2(n4651), .D3(n4548), .S3(n4652), .Z(n2910) );
  HS65_LH_FA1X4 U2221 ( .A0(n1258), .B0(n609), .CI(n624), .CO(n606), .S0(n607)
         );
  HS65_LHS_XOR2X6 U2222 ( .A(n4691), .B(n2870), .Z(n1258) );
  HS65_LH_MX41X7 U2223 ( .D0(n4556), .S0(n1018), .D1(n4550), .S1(n4654), .D2(
        n4553), .S2(n4657), .D3(n4558), .S3(n4658), .Z(n2870) );
  HS65_LH_FA1X4 U2224 ( .A0(n1290), .B0(n607), .CI(n622), .CO(n604), .S0(n605)
         );
  HS65_LHS_XOR2X6 U2225 ( .A(n4689), .B(n2830), .Z(n1290) );
  HS65_LH_MX41X7 U2226 ( .D0(n4567), .S0(n1015), .D1(n4612), .S1(n4665), .D2(
        n4564), .S2(n4663), .D3(n4561), .S3(n4660), .Z(n2830) );
  HS65_LH_FA1X4 U2227 ( .A0(n1126), .B0(n544), .CI(n560), .CO(n541), .S0(n542)
         );
  HS65_LHS_XOR2X6 U2228 ( .A(n4704), .B(n3034), .Z(n1126) );
  HS65_LH_MX41X7 U2229 ( .D0(n3019), .S0(n1026), .D1(n4507), .S1(n4639), .D2(
        n4510), .S2(n4641), .D3(n4515), .S3(n4642), .Z(n3034) );
  HS65_LH_FA1X4 U2230 ( .A0(n1322), .B0(n605), .CI(n620), .CO(n602), .S0(n603)
         );
  HS65_LHS_XOR2X6 U2231 ( .A(n4686), .B(n2791), .Z(n1322) );
  HS65_LH_MX41X7 U2232 ( .D0(n4575), .S0(n1012), .D1(n4569), .S1(n4667), .D2(
        n4572), .S2(n4669), .D3(n4577), .S3(n4670), .Z(n2791) );
  HS65_LH_FA1X4 U2233 ( .A0(n1158), .B0(n542), .CI(n558), .CO(n539), .S0(n540)
         );
  HS65_LHS_XOR2X6 U2234 ( .A(n4701), .B(n2994), .Z(n1158) );
  HS65_LH_MX41X7 U2235 ( .D0(n2976), .S0(n1023), .D1(n4526), .S1(n4648), .D2(
        n4518), .S2(n4645), .D3(n4521), .S3(n4646), .Z(n2994) );
  HS65_LH_FA1X4 U2236 ( .A0(n1091), .B0(n493), .CI(n508), .CO(n491), .S0(n492)
         );
  HS65_LHS_XOR2X6 U2237 ( .A(n4707), .B(n3077), .Z(n1091) );
  HS65_LH_MX41X7 U2238 ( .D0(n4501), .S0(n1026), .D1(n4495), .S1(n4639), .D2(
        n4498), .S2(n4641), .D3(n4504), .S3(n4642), .Z(n3077) );
  HS65_LH_FA1X4 U2239 ( .A0(n1254), .B0(n536), .CI(n552), .CO(n533), .S0(n534)
         );
  HS65_LHS_XOR2X6 U2240 ( .A(n4691), .B(n2874), .Z(n1254) );
  HS65_LH_MX41X7 U2241 ( .D0(n4556), .S0(n1014), .D1(n4550), .S1(n4662), .D2(
        n4553), .S2(n4665), .D3(n4558), .S3(n4666), .Z(n2874) );
  HS65_LH_FA1X4 U2242 ( .A0(n1155), .B0(n490), .CI(n504), .CO(n487), .S0(n488)
         );
  HS65_LHS_XOR2X6 U2243 ( .A(n4701), .B(n2997), .Z(n1155) );
  HS65_LH_MX41X7 U2244 ( .D0(n4523), .S0(n1020), .D1(n4526), .S1(n4655), .D2(
        n4518), .S2(n4651), .D3(n4521), .S3(n4652), .Z(n2997) );
  HS65_LH_FA1X4 U2245 ( .A0(n1098), .B0(n1066), .CI(n634), .CO(n616), .S0(n617) );
  HS65_LH_MX41X7 U2246 ( .D0(n1036), .S0(n4492), .D1(n4622), .S1(n4608), .D2(
        n4620), .S2(n4604), .D3(n4618), .S3(n4609), .Z(n1066) );
  HS65_LHS_XOR2X6 U2247 ( .A(n115), .B(n3070), .Z(n1098) );
  HS65_LH_MX41X7 U2248 ( .D0(n3062), .S0(n1033), .D1(n4496), .S1(n4625), .D2(
        n4499), .S2(n4627), .D3(n4504), .S3(n4628), .Z(n3070) );
  HS65_LH_FA1X4 U2249 ( .A0(n1130), .B0(n617), .CI(n632), .CO(n614), .S0(n615)
         );
  HS65_LHS_XOR2X6 U2250 ( .A(n4704), .B(n3030), .Z(n1130) );
  HS65_LH_MX41X7 U2251 ( .D0(n3019), .S0(n1030), .D1(n4507), .S1(n4630), .D2(
        n4510), .S2(n4633), .D3(n4515), .S3(n4634), .Z(n3030) );
  HS65_LH_FA1X4 U2252 ( .A0(n1162), .B0(n615), .CI(n630), .CO(n612), .S0(n613)
         );
  HS65_LHS_XOR2X6 U2253 ( .A(n4701), .B(n2990), .Z(n1162) );
  HS65_LH_MX41X7 U2254 ( .D0(n2976), .S0(n1027), .D1(n4526), .S1(n4640), .D2(
        n4518), .S2(n4637), .D3(n4521), .S3(n4638), .Z(n2990) );
  HS65_LH_FA1X4 U2255 ( .A0(n1354), .B0(n603), .CI(n618), .CO(n600), .S0(n601)
         );
  HS65_LHS_XOR2X6 U2256 ( .A(n19), .B(n2751), .Z(n1354) );
  HS65_LH_MX41X7 U2257 ( .D0(n4586), .S0(n1009), .D1(n4580), .S1(n4672), .D2(
        n4583), .S2(n4675), .D3(n4588), .S3(n4677), .Z(n2751) );
  HS65_LH_FA1X4 U2258 ( .A0(n1190), .B0(n540), .CI(n556), .CO(n537), .S0(n538)
         );
  HS65_LHS_XOR2X6 U2259 ( .A(n4698), .B(n2954), .Z(n1190) );
  HS65_LH_MX41X7 U2260 ( .D0(n4534), .S0(n1020), .D1(n4529), .S1(n4651), .D2(
        n4532), .S2(n4653), .D3(n4537), .S3(n4654), .Z(n2954) );
  HS65_LH_FA1X4 U2261 ( .A0(n1219), .B0(n486), .CI(n500), .CO(n483), .S0(n484)
         );
  HS65_LHS_XOR2X6 U2262 ( .A(n4694), .B(n2917), .Z(n1219) );
  HS65_LH_MX41X7 U2263 ( .D0(n4545), .S0(n1014), .D1(n4539), .S1(n4663), .D2(
        n4542), .S2(n4665), .D3(n4547), .S3(n4666), .Z(n2917) );
  HS65_LH_FA1X4 U2264 ( .A0(n1120), .B0(n445), .CI(n458), .CO(n442), .S0(n443)
         );
  HS65_LHS_XOR2X6 U2265 ( .A(n4704), .B(n3040), .Z(n1120) );
  HS65_LH_MX41X7 U2266 ( .D0(n3019), .S0(n1020), .D1(n4507), .S1(n4650), .D2(
        n4510), .S2(n4653), .D3(n4515), .S3(n4654), .Z(n3040) );
  HS65_LH_FA1X4 U2267 ( .A0(n1184), .B0(n441), .CI(n454), .CO(n438), .S0(n439)
         );
  HS65_LHS_XOR2X6 U2268 ( .A(n4697), .B(n2960), .Z(n1184) );
  HS65_LH_MX41X7 U2269 ( .D0(n4534), .S0(n1014), .D1(n4528), .S1(n4663), .D2(
        n4531), .S2(n4665), .D3(n4536), .S3(n4666), .Z(n2960) );
  HS65_LH_FA1X4 U2270 ( .A0(n1085), .B0(n406), .CI(n417), .CO(n404), .S0(n405)
         );
  HS65_LHS_XOR2X6 U2271 ( .A(n4706), .B(n3083), .Z(n1085) );
  HS65_LH_MX41X7 U2272 ( .D0(n4501), .S0(n1020), .D1(n4495), .S1(n4651), .D2(
        n4498), .S2(n4653), .D3(n4503), .S3(n4654), .Z(n3083) );
  HS65_LH_FA1X4 U2273 ( .A0(n1149), .B0(n403), .CI(n413), .CO(n400), .S0(n401)
         );
  HS65_LHS_XOR2X6 U2274 ( .A(n4701), .B(n3003), .Z(n1149) );
  HS65_LH_MX41X7 U2275 ( .D0(n2976), .S0(n1014), .D1(n4526), .S1(n4667), .D2(
        n4518), .S2(n4663), .D3(n4521), .S3(n4664), .Z(n3003) );
  HS65_LH_FA1X4 U2276 ( .A0(n1114), .B0(n370), .CI(n379), .CO(n367), .S0(n368)
         );
  HS65_LHS_XOR2X6 U2277 ( .A(n4703), .B(n3046), .Z(n1114) );
  HS65_LH_MX41X7 U2278 ( .D0(n4512), .S0(n1014), .D1(n4506), .S1(n4663), .D2(
        n4509), .S2(n4665), .D3(n4514), .S3(n4666), .Z(n3046) );
  HS65_LH_FA1X4 U2279 ( .A0(n1079), .B0(n343), .CI(n350), .CO(n341), .S0(n342)
         );
  HS65_LHS_XOR2X6 U2280 ( .A(n4706), .B(n3089), .Z(n1079) );
  HS65_LH_MX41X7 U2281 ( .D0(n4501), .S0(n1014), .D1(n4495), .S1(n4663), .D2(
        n4499), .S2(n4665), .D3(n4503), .S3(n4666), .Z(n3089) );
  HS65_LH_FA1X4 U2282 ( .A0(n597), .B0(n614), .CI(n1161), .CO(n594), .S0(n595)
         );
  HS65_LHS_XOR2X6 U2283 ( .A(n4700), .B(n2991), .Z(n1161) );
  HS65_LH_MX41X7 U2284 ( .D0(n4523), .S0(n1026), .D1(n4525), .S1(n4642), .D2(
        n4517), .S2(n4639), .D3(n4520), .S3(n4640), .Z(n2991) );
  HS65_LH_FA1X4 U2285 ( .A0(n579), .B0(n1128), .CI(n1160), .CO(n576), .S0(n577) );
  HS65_LHS_XOR2X6 U2286 ( .A(n4700), .B(n2992), .Z(n1160) );
  HS65_LHS_XOR2X6 U2287 ( .A(n4704), .B(n3032), .Z(n1128) );
  HS65_LH_MX41X7 U2288 ( .D0(n4523), .S0(n1025), .D1(n4525), .S1(n4644), .D2(
        n4517), .S2(n4641), .D3(n4520), .S3(n4642), .Z(n2992) );
  HS65_LH_FA1X4 U2289 ( .A0(n593), .B0(n610), .CI(n1225), .CO(n590), .S0(n591)
         );
  HS65_LHS_XOR2X6 U2290 ( .A(n4694), .B(n2911), .Z(n1225) );
  HS65_LH_MX41X7 U2291 ( .D0(n4545), .S0(n1020), .D1(n4539), .S1(n4650), .D2(
        n4542), .S2(n4653), .D3(n4547), .S3(n4654), .Z(n2911) );
  HS65_LH_FA1X4 U2292 ( .A0(n562), .B0(n545), .CI(n1094), .CO(n543), .S0(n544)
         );
  HS65_LHS_XOR2X6 U2293 ( .A(n115), .B(n3074), .Z(n1094) );
  HS65_LH_MX41X7 U2294 ( .D0(n3062), .S0(n1029), .D1(n4496), .S1(n4632), .D2(
        n4500), .S2(n4635), .D3(n4505), .S3(n4636), .Z(n3074) );
  HS65_LH_FA1X4 U2295 ( .A0(n575), .B0(n1192), .CI(n1224), .CO(n572), .S0(n573) );
  HS65_LHS_XOR2X6 U2296 ( .A(n4694), .B(n2912), .Z(n1224) );
  HS65_LHS_XOR2X6 U2297 ( .A(n4697), .B(n2952), .Z(n1192) );
  HS65_LH_MX41X7 U2298 ( .D0(n4545), .S0(n1019), .D1(n4539), .S1(n4653), .D2(
        n4542), .S2(n4655), .D3(n4547), .S3(n4656), .Z(n2912) );
  HS65_LH_FA1X4 U2299 ( .A0(n527), .B0(n543), .CI(n1125), .CO(n524), .S0(n525)
         );
  HS65_LHS_XOR2X6 U2300 ( .A(n4704), .B(n3035), .Z(n1125) );
  HS65_LH_MX41X7 U2301 ( .D0(n4512), .S0(n1025), .D1(n4507), .S1(n4640), .D2(
        n4510), .S2(n4643), .D3(n4515), .S3(n4644), .Z(n3035) );
  HS65_LH_FA1X4 U2302 ( .A0(n554), .B0(n538), .CI(n1222), .CO(n535), .S0(n536)
         );
  HS65_LHS_XOR2X6 U2303 ( .A(n4694), .B(n2914), .Z(n1222) );
  HS65_LH_MX41X7 U2304 ( .D0(n4545), .S0(n1017), .D1(n4539), .S1(n4656), .D2(
        n4542), .S2(n4659), .D3(n4547), .S3(n4660), .Z(n2914) );
  HS65_LH_FA1X4 U2305 ( .A0(n523), .B0(n539), .CI(n1189), .CO(n520), .S0(n521)
         );
  HS65_LHS_XOR2X6 U2306 ( .A(n4697), .B(n2955), .Z(n1189) );
  HS65_LH_MX41X7 U2307 ( .D0(n4534), .S0(n1019), .D1(n4528), .S1(n4652), .D2(
        n4531), .S2(n4655), .D3(n4536), .S3(n4656), .Z(n2955) );
  HS65_LH_FA1X4 U2308 ( .A0(n567), .B0(n1320), .CI(n1352), .CO(n564), .S0(n565) );
  HS65_LHS_XOR2X6 U2309 ( .A(n19), .B(n2755), .Z(n1352) );
  HS65_LHS_XOR2X6 U2310 ( .A(n4686), .B(n2793), .Z(n1320) );
  HS65_LH_OAI21X3 U2311 ( .A(n4719), .B(n4587), .C(n2756), .Z(n2755) );
  HS65_LH_FA1X4 U2312 ( .A0(n506), .B0(n492), .CI(n1123), .CO(n489), .S0(n490)
         );
  HS65_LHS_XOR2X6 U2313 ( .A(n103), .B(n3037), .Z(n1123) );
  HS65_LH_MX41X7 U2314 ( .D0(n3019), .S0(n1023), .D1(n4507), .S1(n4644), .D2(
        n4511), .S2(n4647), .D3(n4516), .S3(n4648), .Z(n3037) );
  HS65_LH_FA1X4 U2315 ( .A0(n333), .B0(n339), .CI(n1142), .CO(n330), .S0(n331)
         );
  HS65_LHS_XOR2X6 U2316 ( .A(n91), .B(n3012), .Z(n1142) );
  HS65_LH_OAI21X3 U2317 ( .A(n4719), .B(n4524), .C(n3013), .Z(n3012) );
  HS65_LH_OAI22X6 U2318 ( .A(n4676), .B(n3014), .C(n4517), .D(n3014), .Z(n3013) );
  HS65_LH_FA1X4 U2319 ( .A0(n314), .B0(n318), .CI(n1107), .CO(n311), .S0(n312)
         );
  HS65_LHS_XOR2X6 U2320 ( .A(n103), .B(n3055), .Z(n1107) );
  HS65_LH_OAI21X3 U2321 ( .A(n4719), .B(n4513), .C(n3056), .Z(n3055) );
  HS65_LH_OAI22X6 U2322 ( .A(n4676), .B(n3057), .C(n4506), .D(n3057), .Z(n3056) );
  HS65_LH_FA1X4 U2323 ( .A0(n4710), .B0(n1058), .CI(n1090), .CO(n476), .S0(
        n477) );
  HS65_LH_MX41X7 U2324 ( .D0(n1028), .S0(n4491), .D1(n4638), .S1(n4607), .D2(
        n4636), .S2(n4603), .D3(n4634), .S3(n4609), .Z(n1058) );
  HS65_LHS_XOR2X6 U2325 ( .A(n4706), .B(n3078), .Z(n1090) );
  HS65_LH_MX41X7 U2326 ( .D0(n4501), .S0(n1025), .D1(n4495), .S1(n4640), .D2(
        n4498), .S2(n4643), .D3(n4503), .S3(n4644), .Z(n3078) );
  HS65_LH_FA1X4 U2327 ( .A0(n550), .B0(n534), .CI(n1286), .CO(n531), .S0(n532)
         );
  HS65_LHS_XOR2X6 U2328 ( .A(n43), .B(n2834), .Z(n1286) );
  HS65_LH_MX41X7 U2329 ( .D0(n2804), .S0(n1011), .D1(n4613), .S1(n4673), .D2(
        n4565), .S2(n4671), .D3(n4562), .S3(n4668), .Z(n2834) );
  HS65_LH_FA1X4 U2330 ( .A0(n519), .B0(n535), .CI(n1253), .CO(n516), .S0(n517)
         );
  HS65_LHS_XOR2X6 U2331 ( .A(n4691), .B(n2875), .Z(n1253) );
  HS65_LH_MX41X7 U2332 ( .D0(n4556), .S0(n1013), .D1(n4550), .S1(n4665), .D2(
        n4553), .S2(n4667), .D3(n4558), .S3(n4668), .Z(n2875) );
  HS65_LH_FA1X4 U2333 ( .A0(n502), .B0(n488), .CI(n1187), .CO(n485), .S0(n486)
         );
  HS65_LHS_XOR2X6 U2334 ( .A(n79), .B(n2957), .Z(n1187) );
  HS65_LH_MX41X7 U2335 ( .D0(n2933), .S0(n1017), .D1(n4529), .S1(n4656), .D2(
        n4533), .S2(n4659), .D3(n4538), .S3(n4660), .Z(n2957) );
  HS65_LH_FA1X4 U2336 ( .A0(n475), .B0(n489), .CI(n1154), .CO(n472), .S0(n473)
         );
  HS65_LHS_XOR2X6 U2337 ( .A(n4701), .B(n2998), .Z(n1154) );
  HS65_LH_MX41X7 U2338 ( .D0(n4523), .S0(n1019), .D1(n4525), .S1(n4657), .D2(
        n4517), .S2(n4653), .D3(n4520), .S3(n4654), .Z(n2998) );
  HS65_LH_FA1X4 U2339 ( .A0(n515), .B0(n531), .CI(n1317), .CO(n512), .S0(n513)
         );
  HS65_LHS_XOR2X6 U2340 ( .A(n31), .B(n2798), .Z(n1317) );
  HS65_LH_OAI21X3 U2341 ( .A(n4719), .B(n4576), .C(n2799), .Z(n2798) );
  HS65_LH_OAI22X6 U2342 ( .A(n4676), .B(n2800), .C(n4569), .D(n2800), .Z(n2799) );
  HS65_LH_FA1X4 U2343 ( .A0(n460), .B0(n447), .CI(n1088), .CO(n444), .S0(n445)
         );
  HS65_LHS_XOR2X6 U2344 ( .A(n4707), .B(n3080), .Z(n1088) );
  HS65_LH_MX41X7 U2345 ( .D0(n3062), .S0(n1023), .D1(n4496), .S1(n4644), .D2(
        n4499), .S2(n4647), .D3(n4504), .S3(n4648), .Z(n3080) );
  HS65_LH_FA1X4 U2346 ( .A0(n498), .B0(n484), .CI(n1251), .CO(n481), .S0(n482)
         );
  HS65_LHS_XOR2X6 U2347 ( .A(n4691), .B(n2877), .Z(n1251) );
  HS65_LH_MX41X7 U2348 ( .D0(n4556), .S0(n1011), .D1(n4550), .S1(n4668), .D2(
        n4553), .S2(n4671), .D3(n4558), .S3(n4672), .Z(n2877) );
  HS65_LH_FA1X4 U2349 ( .A0(n471), .B0(n485), .CI(n1218), .CO(n468), .S0(n469)
         );
  HS65_LHS_XOR2X6 U2350 ( .A(n4694), .B(n2918), .Z(n1218) );
  HS65_LH_MX41X7 U2351 ( .D0(n4545), .S0(n1013), .D1(n4539), .S1(n4664), .D2(
        n4542), .S2(n4667), .D3(n4547), .S3(n4668), .Z(n2918) );
  HS65_LH_FA1X4 U2352 ( .A0(n456), .B0(n443), .CI(n1152), .CO(n440), .S0(n441)
         );
  HS65_LHS_XOR2X6 U2353 ( .A(n4700), .B(n3000), .Z(n1152) );
  HS65_LH_MX41X7 U2354 ( .D0(n2976), .S0(n1017), .D1(n4527), .S1(n4661), .D2(
        n4518), .S2(n4657), .D3(n4522), .S3(n4658), .Z(n3000) );
  HS65_LH_FA1X4 U2355 ( .A0(n432), .B0(n444), .CI(n1119), .CO(n429), .S0(n430)
         );
  HS65_LHS_XOR2X6 U2356 ( .A(n4703), .B(n3041), .Z(n1119) );
  HS65_LH_MX41X7 U2357 ( .D0(n4512), .S0(n1019), .D1(n4506), .S1(n4653), .D2(
        n4509), .S2(n4655), .D3(n4514), .S3(n4656), .Z(n3041) );
  HS65_LH_FA1X4 U2358 ( .A0(n467), .B0(n481), .CI(n1282), .CO(n464), .S0(n465)
         );
  HS65_LHS_XOR2X6 U2359 ( .A(n43), .B(n2840), .Z(n1282) );
  HS65_LH_OAI21X3 U2360 ( .A(n4719), .B(n4568), .C(n2841), .Z(n2840) );
  HS65_LH_OAI22X6 U2361 ( .A(n4676), .B(n2842), .C(n4561), .D(n2842), .Z(n2841) );
  HS65_LH_FA1X4 U2362 ( .A0(n452), .B0(n439), .CI(n1216), .CO(n436), .S0(n437)
         );
  HS65_LHS_XOR2X6 U2363 ( .A(n4694), .B(n2920), .Z(n1216) );
  HS65_LH_MX41X7 U2364 ( .D0(n4545), .S0(n1011), .D1(n4539), .S1(n4668), .D2(
        n4542), .S2(n4671), .D3(n4547), .S3(n4672), .Z(n2920) );
  HS65_LH_FA1X4 U2365 ( .A0(n428), .B0(n440), .CI(n1183), .CO(n425), .S0(n426)
         );
  HS65_LHS_XOR2X6 U2366 ( .A(n4698), .B(n2961), .Z(n1183) );
  HS65_LH_MX41X7 U2367 ( .D0(n2933), .S0(n1013), .D1(n4529), .S1(n4664), .D2(
        n4532), .S2(n4667), .D3(n4537), .S3(n4668), .Z(n2961) );
  HS65_LH_FA1X4 U2368 ( .A0(n415), .B0(n405), .CI(n1117), .CO(n402), .S0(n403)
         );
  HS65_LHS_XOR2X6 U2369 ( .A(n4703), .B(n3043), .Z(n1117) );
  HS65_LH_MX41X7 U2370 ( .D0(n4512), .S0(n1017), .D1(n4506), .S1(n4657), .D2(
        n4509), .S2(n4659), .D3(n4514), .S3(n4660), .Z(n3043) );
  HS65_LH_FA1X4 U2371 ( .A0(n424), .B0(n436), .CI(n1247), .CO(n421), .S0(n422)
         );
  HS65_LHS_XOR2X6 U2372 ( .A(n55), .B(n2883), .Z(n1247) );
  HS65_LH_OAI21X3 U2373 ( .A(n4719), .B(n4557), .C(n2884), .Z(n2883) );
  HS65_LH_OAI22X6 U2374 ( .A(n4676), .B(n2885), .C(n4550), .D(n2885), .Z(n2884) );
  HS65_LH_FA1X4 U2375 ( .A0(n4711), .B0(n1053), .CI(n1084), .CO(n393), .S0(
        n394) );
  HS65_LH_MX41X7 U2376 ( .D0(n1022), .S0(n4491), .D1(n4646), .S1(n4610), .D2(
        n4648), .S2(n4602), .D3(n4650), .S3(n4606), .Z(n1053) );
  HS65_LHS_XOR2X6 U2377 ( .A(n4706), .B(n3084), .Z(n1084) );
  HS65_LH_MX41X7 U2378 ( .D0(n4501), .S0(n1019), .D1(n4495), .S1(n4653), .D2(
        n4498), .S2(n4655), .D3(n4503), .S3(n4656), .Z(n3084) );
  HS65_LH_FA1X4 U2379 ( .A0(n411), .B0(n401), .CI(n1181), .CO(n398), .S0(n399)
         );
  HS65_LHS_XOR2X6 U2380 ( .A(n79), .B(n2963), .Z(n1181) );
  HS65_LH_MX41X7 U2381 ( .D0(n2933), .S0(n1011), .D1(n4529), .S1(n4669), .D2(
        n4532), .S2(n4671), .D3(n4538), .S3(n4672), .Z(n2963) );
  HS65_LH_FA1X4 U2382 ( .A0(n392), .B0(n402), .CI(n1148), .CO(n389), .S0(n390)
         );
  HS65_LHS_XOR2X6 U2383 ( .A(n4700), .B(n3004), .Z(n1148) );
  HS65_LH_MX41X7 U2384 ( .D0(n4523), .S0(n1013), .D1(n4525), .S1(n4669), .D2(
        n4517), .S2(n4665), .D3(n4520), .S3(n4666), .Z(n3004) );
  HS65_LH_FA1X4 U2385 ( .A0(n381), .B0(n372), .CI(n1082), .CO(n369), .S0(n370)
         );
  HS65_LHS_XOR2X6 U2386 ( .A(n4707), .B(n3086), .Z(n1082) );
  HS65_LH_MX41X7 U2387 ( .D0(n4501), .S0(n1017), .D1(n4496), .S1(n4657), .D2(
        n4499), .S2(n4659), .D3(n4504), .S3(n4660), .Z(n3086) );
  HS65_LH_FA1X4 U2388 ( .A0(n388), .B0(n398), .CI(n1212), .CO(n385), .S0(n386)
         );
  HS65_LHS_XOR2X6 U2389 ( .A(n67), .B(n2926), .Z(n1212) );
  HS65_LH_OAI21X3 U2390 ( .A(n4719), .B(n4546), .C(n2927), .Z(n2926) );
  HS65_LH_OAI22X6 U2391 ( .A(n4676), .B(n2928), .C(n4539), .D(n2928), .Z(n2927) );
  HS65_LH_FA1X4 U2392 ( .A0(n377), .B0(n368), .CI(n1146), .CO(n365), .S0(n366)
         );
  HS65_LHS_XOR2X6 U2393 ( .A(n4700), .B(n3006), .Z(n1146) );
  HS65_LH_MX41X7 U2394 ( .D0(n4523), .S0(n1011), .D1(n4525), .S1(n4673), .D2(
        n4517), .S2(n4669), .D3(n4520), .S3(n4670), .Z(n3006) );
  HS65_LH_FA1X4 U2395 ( .A0(n361), .B0(n369), .CI(n1113), .CO(n358), .S0(n359)
         );
  HS65_LHS_XOR2X6 U2396 ( .A(n4703), .B(n3047), .Z(n1113) );
  HS65_LH_MX41X7 U2397 ( .D0(n4512), .S0(n1013), .D1(n4506), .S1(n4665), .D2(
        n4509), .S2(n4667), .D3(n4514), .S3(n4668), .Z(n3047) );
  HS65_LH_FA1X4 U2398 ( .A0(n357), .B0(n365), .CI(n1177), .CO(n354), .S0(n355)
         );
  HS65_LHS_XOR2X6 U2399 ( .A(n4697), .B(n2969), .Z(n1177) );
  HS65_LH_OAI21X3 U2400 ( .A(n4719), .B(n4535), .C(n2970), .Z(n2969) );
  HS65_LH_OAI22X6 U2401 ( .A(n4676), .B(n2971), .C(n4528), .D(n2971), .Z(n2970) );
  HS65_LH_FA1X4 U2402 ( .A0(n348), .B0(n342), .CI(n1111), .CO(n339), .S0(n340)
         );
  HS65_LHS_XOR2X6 U2403 ( .A(n4703), .B(n3049), .Z(n1111) );
  HS65_LH_MX41X7 U2404 ( .D0(n4512), .S0(n1011), .D1(n4506), .S1(n4669), .D2(
        n4509), .S2(n4671), .D3(n4514), .S3(n4672), .Z(n3049) );
  HS65_LH_FA1X4 U2405 ( .A0(n4712), .B0(n1048), .CI(n1078), .CO(n334), .S0(
        n335) );
  HS65_LH_MX41X7 U2406 ( .D0(n1016), .S0(n4491), .D1(n4658), .S1(n4610), .D2(
        n4660), .S2(n4602), .D3(n4662), .S3(n4606), .Z(n1048) );
  HS65_LHS_XOR2X6 U2407 ( .A(n4706), .B(n3090), .Z(n1078) );
  HS65_LH_MX41X7 U2408 ( .D0(n4501), .S0(n1013), .D1(n4495), .S1(n4665), .D2(
        n4498), .S2(n4667), .D3(n4503), .S3(n4668), .Z(n3090) );
  HS65_LH_FA1X4 U2409 ( .A0(n326), .B0(n321), .CI(n1076), .CO(n318), .S0(n319)
         );
  HS65_LHS_XOR2X6 U2410 ( .A(n4707), .B(n3092), .Z(n1076) );
  HS65_LH_MX41X7 U2411 ( .D0(n4501), .S0(n1011), .D1(n4496), .S1(n4668), .D2(
        n4499), .S2(n4671), .D3(n4504), .S3(n4672), .Z(n3092) );
  HS65_LH_FA1X4 U2412 ( .A0(n4716), .B0(n1043), .CI(n1072), .CO(n299), .S0(
        n300) );
  HS65_LH_MX41X7 U2413 ( .D0(n1010), .S0(n4491), .D1(n4670), .S1(n4610), .D2(
        n4672), .S2(n4603), .D3(n4674), .S3(n4607), .Z(n1043) );
  HS65_LHS_XOR2X6 U2414 ( .A(n4707), .B(n3098), .Z(n1072) );
  HS65_LH_OAI21X3 U2415 ( .A(n4719), .B(n4502), .C(n3099), .Z(n3098) );
  HS65_LH_FA1X4 U2416 ( .A0(n293), .B0(n292), .CI(n228), .CO(n227), .S0(
        product[62]) );
  HS65_LH_HA1X4 U2417 ( .A0(n4680), .B0(n1419), .CO(n289), .S0(product[0]) );
  HS65_LHS_XOR2X6 U2418 ( .A(n7), .B(n2676), .Z(n1419) );
  HS65_LH_AO22X9 U2419 ( .A(n4616), .B(n4600), .C(n4493), .D(n4616), .Z(n2676)
         );
  HS65_LH_HA1X4 U2420 ( .A0(n1418), .B0(n289), .CO(n288), .S0(product[1]) );
  HS65_LHS_XOR2X6 U2421 ( .A(n7), .B(n2678), .Z(n1418) );
  HS65_LH_AO222X4 U2422 ( .A(n4617), .B(n4596), .C(n4598), .D(n4619), .E(n4493), .F(n1038), .Z(n2678) );
  HS65_LH_IVX9 U2423 ( .A(n4687), .Z(n4685) );
  HS65_LH_IVX9 U2424 ( .A(n4693), .Z(n4692) );
  HS65_LH_IVX9 U2425 ( .A(n4687), .Z(n4686) );
  HS65_LH_IVX9 U2426 ( .A(n4693), .Z(n4691) );
  HS65_LH_IVX9 U2427 ( .A(n4696), .Z(n4695) );
  HS65_LH_IVX9 U2428 ( .A(n4696), .Z(n4694) );
  HS65_LH_IVX9 U2429 ( .A(n4708), .Z(n4706) );
  HS65_LH_IVX9 U2430 ( .A(n4708), .Z(n4707) );
  HS65_LH_IVX9 U2431 ( .A(n4699), .Z(n4697) );
  HS65_LH_IVX9 U2432 ( .A(n4699), .Z(n4698) );
  HS65_LH_IVX9 U2433 ( .A(n4690), .Z(n4688) );
  HS65_LH_IVX9 U2434 ( .A(n4690), .Z(n4689) );
  HS65_LH_IVX9 U2435 ( .A(n4705), .Z(n4704) );
  HS65_LH_IVX9 U2436 ( .A(n4705), .Z(n4703) );
  HS65_LH_IVX9 U2437 ( .A(n4702), .Z(n4700) );
  HS65_LH_IVX9 U2438 ( .A(n4702), .Z(n4701) );
  HS65_LH_MX41X7 U2439 ( .D0(n1025), .S0(n4491), .D1(n4644), .S1(n4607), .D2(
        n4642), .S2(n4603), .D3(n4640), .S3(n4609), .Z(n419) );
  HS65_LH_MX41X7 U2440 ( .D0(n1019), .S0(n4491), .D1(n4652), .S1(n4610), .D2(
        n4654), .S2(n4603), .D3(n4656), .S3(n4607), .Z(n352) );
  HS65_LH_MX41X7 U2441 ( .D0(n1013), .S0(n4490), .D1(n4664), .S1(n4610), .D2(
        n4666), .S2(n4602), .D3(n4668), .S3(n4606), .Z(n309) );
  HS65_LH_IVX9 U2442 ( .A(n4684), .Z(n4683) );
  HS65_LH_IVX9 U2443 ( .A(n19), .Z(n4684) );
  HS65_LH_HA1X4 U2444 ( .A0(n1417), .B0(n288), .CO(n287), .S0(product[2]) );
  HS65_LHS_XOR2X6 U2445 ( .A(n4680), .B(n2680), .Z(n1417) );
  HS65_LH_MX41X7 U2446 ( .D0(n1037), .S0(n4493), .D1(n4591), .S1(n4616), .D2(
        n4594), .S2(n4619), .D3(n4620), .S3(n4598), .Z(n2680) );
  HS65_LH_FA1X4 U2447 ( .A0(n1416), .B0(n941), .CI(n287), .CO(n286), .S0(
        product[3]) );
  HS65_LHS_XOR2X6 U2448 ( .A(n4681), .B(n2682), .Z(n1416) );
  HS65_LH_MX41X7 U2449 ( .D0(n1036), .S0(n4493), .D1(n4591), .S1(n4618), .D2(
        n4620), .S2(n4595), .D3(n4622), .S3(n4599), .Z(n2682) );
  HS65_LH_FA1X4 U2450 ( .A0(n1415), .B0(n939), .CI(n286), .CO(n285), .S0(
        product[4]) );
  HS65_LHS_XOR2X6 U2451 ( .A(n4681), .B(n2683), .Z(n1415) );
  HS65_LH_MX41X7 U2452 ( .D0(n1035), .S0(n4493), .D1(n4591), .S1(n4621), .D2(
        n4622), .S2(n4595), .D3(n4624), .S3(n4599), .Z(n2683) );
  HS65_LH_FA1X4 U2453 ( .A0(n1414), .B0(n937), .CI(n285), .CO(n284), .S0(
        product[5]) );
  HS65_LHS_XOR2X6 U2454 ( .A(n7), .B(n2684), .Z(n1414) );
  HS65_LH_MX41X7 U2455 ( .D0(n1034), .S0(n4494), .D1(n4622), .S1(n4592), .D2(
        n4624), .S2(n4596), .D3(n4626), .S3(n4600), .Z(n2684) );
  HS65_LH_FA1X4 U2456 ( .A0(n1413), .B0(n933), .CI(n284), .CO(n283), .S0(
        product[6]) );
  HS65_LHS_XOR2X6 U2457 ( .A(n4681), .B(n2685), .Z(n1413) );
  HS65_LH_MX41X7 U2458 ( .D0(n1033), .S0(n4493), .D1(n4624), .S1(n4592), .D2(
        n4626), .S2(n4595), .D3(n4628), .S3(n4599), .Z(n2685) );
  HS65_LH_FA1X4 U2459 ( .A0(n1380), .B0(n931), .CI(n932), .CO(n928), .S0(n929)
         );
  HS65_LHS_XOR2X6 U2460 ( .A(n4683), .B(n2725), .Z(n1380) );
  HS65_LH_MX41X7 U2461 ( .D0(n2719), .S0(n1035), .D1(n4581), .S1(n4621), .D2(
        n4584), .S2(n4623), .D3(n4590), .S3(n4624), .Z(n2725) );
  HS65_LH_FA1X4 U2462 ( .A0(n1412), .B0(n929), .CI(n283), .CO(n282), .S0(
        product[7]) );
  HS65_LHS_XOR2X6 U2463 ( .A(n4681), .B(n2686), .Z(n1412) );
  HS65_LH_MX41X7 U2464 ( .D0(n1032), .S0(n4493), .D1(n4626), .S1(n4592), .D2(
        n4628), .S2(n4595), .D3(n4630), .S3(n4599), .Z(n2686) );
  HS65_LH_FA1X4 U2465 ( .A0(n1379), .B0(n927), .CI(n928), .CO(n924), .S0(n925)
         );
  HS65_LHS_XOR2X6 U2466 ( .A(n4683), .B(n2726), .Z(n1379) );
  HS65_LH_MX41X7 U2467 ( .D0(n2719), .S0(n1034), .D1(n4580), .S1(n4622), .D2(
        n4585), .S2(n4625), .D3(n4590), .S3(n4626), .Z(n2726) );
  HS65_LH_FA1X4 U2468 ( .A0(n1411), .B0(n925), .CI(n282), .CO(n281), .S0(
        product[8]) );
  HS65_LHS_XOR2X6 U2469 ( .A(n4680), .B(n2687), .Z(n1411) );
  HS65_LH_MX41X7 U2470 ( .D0(n1031), .S0(n4493), .D1(n4628), .S1(n4592), .D2(
        n4630), .S2(n4595), .D3(n4632), .S3(n4599), .Z(n2687) );
  HS65_LH_FA1X4 U2471 ( .A0(n1345), .B0(n917), .CI(n920), .CO(n914), .S0(n915)
         );
  HS65_LHS_XOR2X6 U2472 ( .A(n4685), .B(n2768), .Z(n1345) );
  HS65_LH_MX41X7 U2473 ( .D0(n2762), .S0(n1035), .D1(n4570), .S1(n4621), .D2(
        n4573), .S2(n4623), .D3(n4579), .S3(n4624), .Z(n2768) );
  HS65_LH_FA1X4 U2474 ( .A0(n1378), .B0(n921), .CI(n924), .CO(n918), .S0(n919)
         );
  HS65_LHS_XOR2X6 U2475 ( .A(n4683), .B(n2727), .Z(n1378) );
  HS65_LH_MX41X7 U2476 ( .D0(n4586), .S0(n1033), .D1(n4580), .S1(n4624), .D2(
        n4583), .S2(n4627), .D3(n4588), .S3(n4628), .Z(n2727) );
  HS65_LH_FA1X4 U2477 ( .A0(n1410), .B0(n919), .CI(n281), .CO(n280), .S0(
        product[9]) );
  HS65_LHS_XOR2X6 U2478 ( .A(n4680), .B(n2688), .Z(n1410) );
  HS65_LH_MX41X7 U2479 ( .D0(n1030), .S0(n4493), .D1(n4630), .S1(n4591), .D2(
        n4632), .S2(n4595), .D3(n4634), .S3(n4599), .Z(n2688) );
  HS65_LH_FA1X4 U2480 ( .A0(n1344), .B0(n911), .CI(n914), .CO(n908), .S0(n909)
         );
  HS65_LHS_XOR2X6 U2481 ( .A(n4686), .B(n2769), .Z(n1344) );
  HS65_LH_MX41X7 U2482 ( .D0(n2762), .S0(n1034), .D1(n4569), .S1(n4623), .D2(
        n4574), .S2(n4625), .D3(n4579), .S3(n4626), .Z(n2769) );
  HS65_LH_FA1X4 U2483 ( .A0(n1377), .B0(n915), .CI(n918), .CO(n912), .S0(n913)
         );
  HS65_LHS_XOR2X6 U2484 ( .A(n19), .B(n2728), .Z(n1377) );
  HS65_LH_MX41X7 U2485 ( .D0(n4586), .S0(n1032), .D1(n4580), .S1(n4627), .D2(
        n4583), .S2(n4629), .D3(n4588), .S3(n4630), .Z(n2728) );
  HS65_LH_FA1X4 U2486 ( .A0(n1409), .B0(n913), .CI(n280), .CO(n279), .S0(
        product[10]) );
  HS65_LHS_XOR2X6 U2487 ( .A(n4680), .B(n2689), .Z(n1409) );
  HS65_LH_MX41X7 U2488 ( .D0(n1029), .S0(n4493), .D1(n4632), .S1(n4592), .D2(
        n4634), .S2(n4595), .D3(n4636), .S3(n4599), .Z(n2689) );
  HS65_LH_FA1X4 U2489 ( .A0(n1310), .B0(n897), .CI(n902), .CO(n894), .S0(n895)
         );
  HS65_LHS_XOR2X6 U2490 ( .A(n4688), .B(n2810), .Z(n1310) );
  HS65_LH_MX41X7 U2491 ( .D0(n2804), .S0(n1035), .D1(n4612), .S1(n4624), .D2(
        n4565), .S2(n4623), .D3(n4562), .S3(n4620), .Z(n2810) );
  HS65_LH_FA1X4 U2492 ( .A0(n1343), .B0(n903), .CI(n908), .CO(n900), .S0(n901)
         );
  HS65_LHS_XOR2X6 U2493 ( .A(n4685), .B(n2770), .Z(n1343) );
  HS65_LH_MX41X7 U2494 ( .D0(n4575), .S0(n1033), .D1(n4569), .S1(n4624), .D2(
        n4572), .S2(n4627), .D3(n4577), .S3(n4628), .Z(n2770) );
  HS65_LH_FA1X4 U2495 ( .A0(n1376), .B0(n909), .CI(n912), .CO(n906), .S0(n907)
         );
  HS65_LHS_XOR2X6 U2496 ( .A(n4683), .B(n2729), .Z(n1376) );
  HS65_LH_MX41X7 U2497 ( .D0(n4586), .S0(n1031), .D1(n4580), .S1(n4629), .D2(
        n4583), .S2(n4631), .D3(n4588), .S3(n4632), .Z(n2729) );
  HS65_LH_FA1X4 U2498 ( .A0(n1408), .B0(n907), .CI(n279), .CO(n278), .S0(
        product[11]) );
  HS65_LHS_XOR2X6 U2499 ( .A(n4680), .B(n2690), .Z(n1408) );
  HS65_LH_MX41X7 U2500 ( .D0(n1028), .S0(n4493), .D1(n4634), .S1(n4592), .D2(
        n4636), .S2(n4595), .D3(n4638), .S3(n4599), .Z(n2690) );
  HS65_LH_FA1X4 U2501 ( .A0(n1309), .B0(n889), .CI(n894), .CO(n886), .S0(n887)
         );
  HS65_LHS_XOR2X6 U2502 ( .A(n4689), .B(n2811), .Z(n1309) );
  HS65_LH_MX41X7 U2503 ( .D0(n2804), .S0(n1034), .D1(n4613), .S1(n4626), .D2(
        n4566), .S2(n4625), .D3(n4561), .S3(n4622), .Z(n2811) );
  HS65_LH_FA1X4 U2504 ( .A0(n1342), .B0(n895), .CI(n900), .CO(n892), .S0(n893)
         );
  HS65_LHS_XOR2X6 U2505 ( .A(n4685), .B(n2771), .Z(n1342) );
  HS65_LH_MX41X7 U2506 ( .D0(n4575), .S0(n1032), .D1(n4569), .S1(n4627), .D2(
        n4572), .S2(n4629), .D3(n4577), .S3(n4630), .Z(n2771) );
  HS65_LH_FA1X4 U2507 ( .A0(n1375), .B0(n901), .CI(n906), .CO(n898), .S0(n899)
         );
  HS65_LHS_XOR2X6 U2508 ( .A(n19), .B(n2730), .Z(n1375) );
  HS65_LH_MX41X7 U2509 ( .D0(n4586), .S0(n1030), .D1(n4580), .S1(n4631), .D2(
        n4583), .S2(n4633), .D3(n4588), .S3(n4634), .Z(n2730) );
  HS65_LH_FA1X4 U2510 ( .A0(n1407), .B0(n899), .CI(n278), .CO(n277), .S0(
        product[12]) );
  HS65_LHS_XOR2X6 U2511 ( .A(n4681), .B(n2691), .Z(n1407) );
  HS65_LH_MX41X7 U2512 ( .D0(n1027), .S0(n4494), .D1(n4636), .S1(n4592), .D2(
        n4638), .S2(n4595), .D3(n4598), .S3(n4640), .Z(n2691) );
  HS65_LH_FA1X4 U2513 ( .A0(n1275), .B0(n871), .CI(n878), .CO(n868), .S0(n869)
         );
  HS65_LHS_XOR2X6 U2514 ( .A(n4692), .B(n2853), .Z(n1275) );
  HS65_LH_MX41X7 U2515 ( .D0(n2847), .S0(n1035), .D1(n4551), .S1(n4621), .D2(
        n4554), .S2(n4623), .D3(n4560), .S3(n4624), .Z(n2853) );
  HS65_LH_FA1X4 U2516 ( .A0(n1308), .B0(n879), .CI(n886), .CO(n876), .S0(n877)
         );
  HS65_LHS_XOR2X6 U2517 ( .A(n4688), .B(n2812), .Z(n1308) );
  HS65_LH_MX41X7 U2518 ( .D0(n4567), .S0(n1033), .D1(n4611), .S1(n4629), .D2(
        n4564), .S2(n4627), .D3(n4561), .S3(n4624), .Z(n2812) );
  HS65_LH_FA1X4 U2519 ( .A0(n1341), .B0(n887), .CI(n892), .CO(n884), .S0(n885)
         );
  HS65_LHS_XOR2X6 U2520 ( .A(n4685), .B(n2772), .Z(n1341) );
  HS65_LH_MX41X7 U2521 ( .D0(n4575), .S0(n1031), .D1(n4569), .S1(n4629), .D2(
        n4572), .S2(n4631), .D3(n4577), .S3(n4632), .Z(n2772) );
  HS65_LH_FA1X4 U2522 ( .A0(n1374), .B0(n893), .CI(n898), .CO(n890), .S0(n891)
         );
  HS65_LHS_XOR2X6 U2523 ( .A(n4683), .B(n2731), .Z(n1374) );
  HS65_LH_MX41X7 U2524 ( .D0(n4586), .S0(n1029), .D1(n4580), .S1(n4633), .D2(
        n4583), .S2(n4635), .D3(n4588), .S3(n4636), .Z(n2731) );
  HS65_LH_FA1X4 U2525 ( .A0(n1406), .B0(n891), .CI(n277), .CO(n276), .S0(
        product[13]) );
  HS65_LHS_XOR2X6 U2526 ( .A(n4680), .B(n2692), .Z(n1406) );
  HS65_LH_MX41X7 U2527 ( .D0(n1026), .S0(n4493), .D1(n4638), .S1(n4591), .D2(
        n4594), .S2(n4641), .D3(n4598), .S3(n4642), .Z(n2692) );
  HS65_LH_FA1X4 U2528 ( .A0(n1274), .B0(n861), .CI(n868), .CO(n858), .S0(n859)
         );
  HS65_LHS_XOR2X6 U2529 ( .A(n4691), .B(n2854), .Z(n1274) );
  HS65_LH_MX41X7 U2530 ( .D0(n2847), .S0(n1034), .D1(n4550), .S1(n4623), .D2(
        n4555), .S2(n4625), .D3(n4560), .S3(n4626), .Z(n2854) );
  HS65_LH_FA1X4 U2531 ( .A0(n1307), .B0(n869), .CI(n876), .CO(n866), .S0(n867)
         );
  HS65_LHS_XOR2X6 U2532 ( .A(n4688), .B(n2813), .Z(n1307) );
  HS65_LH_MX41X7 U2533 ( .D0(n4567), .S0(n1032), .D1(n4611), .S1(n4631), .D2(
        n4564), .S2(n4629), .D3(n4561), .S3(n4626), .Z(n2813) );
  HS65_LH_FA1X4 U2534 ( .A0(n1340), .B0(n877), .CI(n884), .CO(n874), .S0(n875)
         );
  HS65_LHS_XOR2X6 U2535 ( .A(n4685), .B(n2773), .Z(n1340) );
  HS65_LH_MX41X7 U2536 ( .D0(n4575), .S0(n1030), .D1(n4569), .S1(n4631), .D2(
        n4572), .S2(n4633), .D3(n4577), .S3(n4634), .Z(n2773) );
  HS65_LH_FA1X4 U2537 ( .A0(n1373), .B0(n885), .CI(n890), .CO(n882), .S0(n883)
         );
  HS65_LHS_XOR2X6 U2538 ( .A(n4683), .B(n2732), .Z(n1373) );
  HS65_LH_MX41X7 U2539 ( .D0(n4586), .S0(n1028), .D1(n4580), .S1(n4635), .D2(
        n4583), .S2(n4637), .D3(n4588), .S3(n4638), .Z(n2732) );
  HS65_LH_FA1X4 U2540 ( .A0(n1405), .B0(n883), .CI(n276), .CO(n275), .S0(
        product[14]) );
  HS65_LHS_XOR2X6 U2541 ( .A(n4681), .B(n2693), .Z(n1405) );
  HS65_LH_MX41X7 U2542 ( .D0(n4493), .S0(n1025), .D1(n4591), .S1(n4641), .D2(
        n4594), .S2(n4643), .D3(n4598), .S3(n4644), .Z(n2693) );
  HS65_LH_FA1X4 U2543 ( .A0(n1240), .B0(n839), .CI(n848), .CO(n836), .S0(n837)
         );
  HS65_LHS_XOR2X6 U2544 ( .A(n67), .B(n2896), .Z(n1240) );
  HS65_LH_MX41X7 U2545 ( .D0(n2890), .S0(n1035), .D1(n4540), .S1(n4621), .D2(
        n4543), .S2(n4623), .D3(n4549), .S3(n4624), .Z(n2896) );
  HS65_LH_FA1X4 U2546 ( .A0(n1273), .B0(n849), .CI(n858), .CO(n846), .S0(n847)
         );
  HS65_LHS_XOR2X6 U2547 ( .A(n4692), .B(n2855), .Z(n1273) );
  HS65_LH_MX41X7 U2548 ( .D0(n4556), .S0(n1033), .D1(n4551), .S1(n4625), .D2(
        n4554), .S2(n4627), .D3(n4559), .S3(n4628), .Z(n2855) );
  HS65_LH_FA1X4 U2549 ( .A0(n1306), .B0(n859), .CI(n866), .CO(n856), .S0(n857)
         );
  HS65_LHS_XOR2X6 U2550 ( .A(n4689), .B(n2814), .Z(n1306) );
  HS65_LH_MX41X7 U2551 ( .D0(n4567), .S0(n1031), .D1(n4611), .S1(n4633), .D2(
        n4564), .S2(n4631), .D3(n4561), .S3(n4628), .Z(n2814) );
  HS65_LH_FA1X4 U2552 ( .A0(n1339), .B0(n867), .CI(n874), .CO(n864), .S0(n865)
         );
  HS65_LHS_XOR2X6 U2553 ( .A(n4686), .B(n2774), .Z(n1339) );
  HS65_LH_MX41X7 U2554 ( .D0(n4575), .S0(n1029), .D1(n4569), .S1(n4633), .D2(
        n4572), .S2(n4635), .D3(n4577), .S3(n4636), .Z(n2774) );
  HS65_LH_FA1X4 U2555 ( .A0(n1372), .B0(n875), .CI(n882), .CO(n872), .S0(n873)
         );
  HS65_LHS_XOR2X6 U2556 ( .A(n4683), .B(n2733), .Z(n1372) );
  HS65_LH_MX41X7 U2557 ( .D0(n2719), .S0(n1027), .D1(n4581), .S1(n4637), .D2(
        n4584), .S2(n4639), .D3(n4590), .S3(n4640), .Z(n2733) );
  HS65_LH_FA1X4 U2558 ( .A0(n1404), .B0(n873), .CI(n275), .CO(n274), .S0(
        product[15]) );
  HS65_LHS_XOR2X6 U2559 ( .A(n4681), .B(n2694), .Z(n1404) );
  HS65_LH_MX41X7 U2560 ( .D0(n1024), .S0(n4494), .D1(n4591), .S1(n4643), .D2(
        n4594), .S2(n4645), .D3(n4646), .S3(n4599), .Z(n2694) );
  HS65_LH_FA1X4 U2561 ( .A0(n1239), .B0(n827), .CI(n836), .CO(n824), .S0(n825)
         );
  HS65_LHS_XOR2X6 U2562 ( .A(n4695), .B(n2897), .Z(n1239) );
  HS65_LH_MX41X7 U2563 ( .D0(n2890), .S0(n1034), .D1(n4539), .S1(n4623), .D2(
        n4544), .S2(n4625), .D3(n4549), .S3(n4626), .Z(n2897) );
  HS65_LH_FA1X4 U2564 ( .A0(n1272), .B0(n837), .CI(n846), .CO(n834), .S0(n835)
         );
  HS65_LHS_XOR2X6 U2565 ( .A(n4692), .B(n2856), .Z(n1272) );
  HS65_LH_MX41X7 U2566 ( .D0(n4556), .S0(n1032), .D1(n4550), .S1(n4627), .D2(
        n4554), .S2(n4629), .D3(n4559), .S3(n4630), .Z(n2856) );
  HS65_LH_FA1X4 U2567 ( .A0(n1305), .B0(n847), .CI(n856), .CO(n844), .S0(n845)
         );
  HS65_LHS_XOR2X6 U2568 ( .A(n4688), .B(n2815), .Z(n1305) );
  HS65_LH_MX41X7 U2569 ( .D0(n4567), .S0(n1030), .D1(n4611), .S1(n4635), .D2(
        n4564), .S2(n4633), .D3(n4561), .S3(n4630), .Z(n2815) );
  HS65_LH_FA1X4 U2570 ( .A0(n1338), .B0(n857), .CI(n864), .CO(n854), .S0(n855)
         );
  HS65_LHS_XOR2X6 U2571 ( .A(n4685), .B(n2775), .Z(n1338) );
  HS65_LH_MX41X7 U2572 ( .D0(n4575), .S0(n1028), .D1(n4569), .S1(n4635), .D2(
        n4572), .S2(n4637), .D3(n4577), .S3(n4638), .Z(n2775) );
  HS65_LH_FA1X4 U2573 ( .A0(n1371), .B0(n865), .CI(n872), .CO(n862), .S0(n863)
         );
  HS65_LHS_XOR2X6 U2574 ( .A(n4683), .B(n2734), .Z(n1371) );
  HS65_LH_MX41X7 U2575 ( .D0(n2719), .S0(n1026), .D1(n4581), .S1(n4638), .D2(
        n4584), .S2(n4641), .D3(n4589), .S3(n4642), .Z(n2734) );
  HS65_LH_FA1X4 U2576 ( .A0(n1403), .B0(n863), .CI(n274), .CO(n273), .S0(
        product[16]) );
  HS65_LHS_XOR2X6 U2577 ( .A(n4681), .B(n2695), .Z(n1403) );
  HS65_LH_MX41X7 U2578 ( .D0(n1023), .S0(n4493), .D1(n4591), .S1(n4645), .D2(
        n4646), .S2(n4595), .D3(n4648), .S3(n4599), .Z(n2695) );
  HS65_LH_FA1X4 U2579 ( .A0(n1205), .B0(n801), .CI(n812), .CO(n798), .S0(n799)
         );
  HS65_LHS_XOR2X6 U2580 ( .A(n4698), .B(n2939), .Z(n1205) );
  HS65_LH_MX41X7 U2581 ( .D0(n2933), .S0(n1035), .D1(n4529), .S1(n4620), .D2(
        n4532), .S2(n4623), .D3(n4537), .S3(n4624), .Z(n2939) );
  HS65_LH_FA1X4 U2582 ( .A0(n1238), .B0(n813), .CI(n824), .CO(n810), .S0(n811)
         );
  HS65_LHS_XOR2X6 U2583 ( .A(n4695), .B(n2898), .Z(n1238) );
  HS65_LH_MX41X7 U2584 ( .D0(n2890), .S0(n1033), .D1(n4540), .S1(n4625), .D2(
        n4543), .S2(n4627), .D3(n4548), .S3(n4628), .Z(n2898) );
  HS65_LH_FA1X4 U2585 ( .A0(n1271), .B0(n825), .CI(n834), .CO(n822), .S0(n823)
         );
  HS65_LHS_XOR2X6 U2586 ( .A(n4692), .B(n2857), .Z(n1271) );
  HS65_LH_MX41X7 U2587 ( .D0(n4556), .S0(n1031), .D1(n4550), .S1(n4628), .D2(
        n4553), .S2(n4631), .D3(n4559), .S3(n4632), .Z(n2857) );
  HS65_LH_FA1X4 U2588 ( .A0(n1304), .B0(n835), .CI(n844), .CO(n832), .S0(n833)
         );
  HS65_LHS_XOR2X6 U2589 ( .A(n4688), .B(n2816), .Z(n1304) );
  HS65_LH_MX41X7 U2590 ( .D0(n4567), .S0(n1029), .D1(n4611), .S1(n4637), .D2(
        n4564), .S2(n4635), .D3(n4561), .S3(n4632), .Z(n2816) );
  HS65_LH_FA1X4 U2591 ( .A0(n1337), .B0(n845), .CI(n854), .CO(n842), .S0(n843)
         );
  HS65_LHS_XOR2X6 U2592 ( .A(n4686), .B(n2776), .Z(n1337) );
  HS65_LH_MX41X7 U2593 ( .D0(n2762), .S0(n1027), .D1(n4570), .S1(n4637), .D2(
        n4573), .S2(n4639), .D3(n4578), .S3(n4640), .Z(n2776) );
  HS65_LH_FA1X4 U2594 ( .A0(n1370), .B0(n855), .CI(n862), .CO(n852), .S0(n853)
         );
  HS65_LHS_XOR2X6 U2595 ( .A(n4683), .B(n2735), .Z(n1370) );
  HS65_LH_MX41X7 U2596 ( .D0(n2719), .S0(n1025), .D1(n4581), .S1(n4641), .D2(
        n4584), .S2(n4643), .D3(n4589), .S3(n4644), .Z(n2735) );
  HS65_LH_FA1X4 U2597 ( .A0(n1402), .B0(n853), .CI(n273), .CO(n272), .S0(
        product[17]) );
  HS65_LHS_XOR2X6 U2598 ( .A(n4680), .B(n2696), .Z(n1402) );
  HS65_LH_MX41X7 U2599 ( .D0(n1022), .S0(n4493), .D1(n4646), .S1(n4592), .D2(
        n4648), .S2(n4595), .D3(n4650), .S3(n4598), .Z(n2696) );
  HS65_LH_FA1X4 U2600 ( .A0(n1237), .B0(n799), .CI(n810), .CO(n796), .S0(n797)
         );
  HS65_LHS_XOR2X6 U2601 ( .A(n4695), .B(n2899), .Z(n1237) );
  HS65_LH_MX41X7 U2602 ( .D0(n4545), .S0(n1032), .D1(n4540), .S1(n4627), .D2(
        n4543), .S2(n4629), .D3(n4548), .S3(n4630), .Z(n2899) );
  HS65_LH_FA1X4 U2603 ( .A0(n1270), .B0(n811), .CI(n822), .CO(n808), .S0(n809)
         );
  HS65_LHS_XOR2X6 U2604 ( .A(n4692), .B(n2858), .Z(n1270) );
  HS65_LH_MX41X7 U2605 ( .D0(n4556), .S0(n1030), .D1(n4550), .S1(n4631), .D2(
        n4553), .S2(n4633), .D3(n4558), .S3(n4634), .Z(n2858) );
  HS65_LH_FA1X4 U2606 ( .A0(n1303), .B0(n823), .CI(n832), .CO(n820), .S0(n821)
         );
  HS65_LHS_XOR2X6 U2607 ( .A(n4688), .B(n2817), .Z(n1303) );
  HS65_LH_MX41X7 U2608 ( .D0(n4567), .S0(n1028), .D1(n4611), .S1(n4638), .D2(
        n4564), .S2(n4637), .D3(n4561), .S3(n4634), .Z(n2817) );
  HS65_LH_FA1X4 U2609 ( .A0(n1336), .B0(n833), .CI(n842), .CO(n830), .S0(n831)
         );
  HS65_LHS_XOR2X6 U2610 ( .A(n4686), .B(n2777), .Z(n1336) );
  HS65_LH_MX41X7 U2611 ( .D0(n2762), .S0(n1026), .D1(n4570), .S1(n4639), .D2(
        n4573), .S2(n4641), .D3(n4578), .S3(n4642), .Z(n2777) );
  HS65_LH_FA1X4 U2612 ( .A0(n1369), .B0(n843), .CI(n852), .CO(n840), .S0(n841)
         );
  HS65_LHS_XOR2X6 U2613 ( .A(n19), .B(n2736), .Z(n1369) );
  HS65_LH_MX41X7 U2614 ( .D0(n4586), .S0(n1024), .D1(n4580), .S1(n4643), .D2(
        n4583), .S2(n4645), .D3(n4588), .S3(n4646), .Z(n2736) );
  HS65_LH_FA1X4 U2615 ( .A0(n1401), .B0(n841), .CI(n272), .CO(n271), .S0(
        product[18]) );
  HS65_LHS_XOR2X6 U2616 ( .A(n4680), .B(n2697), .Z(n1401) );
  HS65_LH_MX41X7 U2617 ( .D0(n1021), .S0(n4493), .D1(n4648), .S1(n4591), .D2(
        n4650), .S2(n4594), .D3(n4598), .S3(n4652), .Z(n2697) );
  HS65_LH_FA1X4 U2618 ( .A0(n1170), .B0(n757), .CI(n770), .CO(n754), .S0(n755)
         );
  HS65_LHS_XOR2X6 U2619 ( .A(n4701), .B(n2982), .Z(n1170) );
  HS65_LH_MX41X7 U2620 ( .D0(n2976), .S0(n1035), .D1(n4527), .S1(n4625), .D2(
        n4518), .S2(n4621), .D3(n4521), .S3(n4622), .Z(n2982) );
  HS65_LH_FA1X4 U2621 ( .A0(n1203), .B0(n771), .CI(n784), .CO(n768), .S0(n769)
         );
  HS65_LHS_XOR2X6 U2622 ( .A(n4698), .B(n2941), .Z(n1203) );
  HS65_LH_MX41X7 U2623 ( .D0(n4534), .S0(n1033), .D1(n4529), .S1(n4625), .D2(
        n4532), .S2(n4627), .D3(n4537), .S3(n4628), .Z(n2941) );
  HS65_LH_FA1X4 U2624 ( .A0(n1236), .B0(n785), .CI(n796), .CO(n782), .S0(n783)
         );
  HS65_LHS_XOR2X6 U2625 ( .A(n4695), .B(n2900), .Z(n1236) );
  HS65_LH_MX41X7 U2626 ( .D0(n4545), .S0(n1031), .D1(n4540), .S1(n4628), .D2(
        n4543), .S2(n4631), .D3(n4548), .S3(n4632), .Z(n2900) );
  HS65_LH_FA1X4 U2627 ( .A0(n1269), .B0(n797), .CI(n808), .CO(n794), .S0(n795)
         );
  HS65_LHS_XOR2X6 U2628 ( .A(n4691), .B(n2859), .Z(n1269) );
  HS65_LH_MX41X7 U2629 ( .D0(n4556), .S0(n1029), .D1(n4550), .S1(n4633), .D2(
        n4553), .S2(n4635), .D3(n4558), .S3(n4636), .Z(n2859) );
  HS65_LH_FA1X4 U2630 ( .A0(n1302), .B0(n809), .CI(n820), .CO(n806), .S0(n807)
         );
  HS65_LHS_XOR2X6 U2631 ( .A(n4689), .B(n2818), .Z(n1302) );
  HS65_LH_MX41X7 U2632 ( .D0(n2804), .S0(n1027), .D1(n4612), .S1(n4640), .D2(
        n4565), .S2(n4639), .D3(n4562), .S3(n4636), .Z(n2818) );
  HS65_LH_FA1X4 U2633 ( .A0(n1335), .B0(n821), .CI(n830), .CO(n818), .S0(n819)
         );
  HS65_LHS_XOR2X6 U2634 ( .A(n4686), .B(n2778), .Z(n1335) );
  HS65_LH_MX41X7 U2635 ( .D0(n2762), .S0(n1025), .D1(n4570), .S1(n4641), .D2(
        n4573), .S2(n4643), .D3(n4578), .S3(n4644), .Z(n2778) );
  HS65_LH_FA1X4 U2636 ( .A0(n1368), .B0(n831), .CI(n840), .CO(n828), .S0(n829)
         );
  HS65_LHS_XOR2X6 U2637 ( .A(n4683), .B(n2737), .Z(n1368) );
  HS65_LH_MX41X7 U2638 ( .D0(n2719), .S0(n1023), .D1(n4581), .S1(n4645), .D2(
        n4584), .S2(n4647), .D3(n4589), .S3(n4648), .Z(n2737) );
  HS65_LH_FA1X4 U2639 ( .A0(n1400), .B0(n829), .CI(n271), .CO(n270), .S0(
        product[19]) );
  HS65_LHS_XOR2X6 U2640 ( .A(n7), .B(n2698), .Z(n1400) );
  HS65_LH_MX41X7 U2641 ( .D0(n1020), .S0(n4494), .D1(n4650), .S1(n4592), .D2(
        n4594), .S2(n4653), .D3(n4598), .S3(n4654), .Z(n2698) );
  HS65_LH_FA1X4 U2642 ( .A0(n1169), .B0(n741), .CI(n754), .CO(n738), .S0(n739)
         );
  HS65_LHS_XOR2X6 U2643 ( .A(n91), .B(n2983), .Z(n1169) );
  HS65_LH_MX41X7 U2644 ( .D0(n2976), .S0(n1034), .D1(n4527), .S1(n4627), .D2(
        n4517), .S2(n4623), .D3(n4522), .S3(n4624), .Z(n2983) );
  HS65_LH_FA1X4 U2645 ( .A0(n1202), .B0(n755), .CI(n768), .CO(n752), .S0(n753)
         );
  HS65_LHS_XOR2X6 U2646 ( .A(n4698), .B(n2942), .Z(n1202) );
  HS65_LH_MX41X7 U2647 ( .D0(n4534), .S0(n1032), .D1(n4528), .S1(n4626), .D2(
        n4532), .S2(n4629), .D3(n4537), .S3(n4630), .Z(n2942) );
  HS65_LH_FA1X4 U2648 ( .A0(n1235), .B0(n769), .CI(n782), .CO(n766), .S0(n767)
         );
  HS65_LHS_XOR2X6 U2649 ( .A(n4695), .B(n2901), .Z(n1235) );
  HS65_LH_MX41X7 U2650 ( .D0(n4545), .S0(n1030), .D1(n4540), .S1(n4631), .D2(
        n4543), .S2(n4633), .D3(n4548), .S3(n4634), .Z(n2901) );
  HS65_LH_FA1X4 U2651 ( .A0(n1268), .B0(n783), .CI(n794), .CO(n780), .S0(n781)
         );
  HS65_LHS_XOR2X6 U2652 ( .A(n4691), .B(n2860), .Z(n1268) );
  HS65_LH_MX41X7 U2653 ( .D0(n4556), .S0(n1028), .D1(n4550), .S1(n4635), .D2(
        n4553), .S2(n4637), .D3(n4558), .S3(n4638), .Z(n2860) );
  HS65_LH_FA1X4 U2654 ( .A0(n1301), .B0(n795), .CI(n806), .CO(n792), .S0(n793)
         );
  HS65_LHS_XOR2X6 U2655 ( .A(n4689), .B(n2819), .Z(n1301) );
  HS65_LH_MX41X7 U2656 ( .D0(n2804), .S0(n1026), .D1(n4612), .S1(n4642), .D2(
        n4565), .S2(n4641), .D3(n4562), .S3(n4638), .Z(n2819) );
  HS65_LH_FA1X4 U2657 ( .A0(n1334), .B0(n807), .CI(n818), .CO(n804), .S0(n805)
         );
  HS65_LHS_XOR2X6 U2658 ( .A(n4685), .B(n2779), .Z(n1334) );
  HS65_LH_MX41X7 U2659 ( .D0(n4575), .S0(n1024), .D1(n4569), .S1(n4643), .D2(
        n4572), .S2(n4645), .D3(n4577), .S3(n4646), .Z(n2779) );
  HS65_LH_FA1X4 U2660 ( .A0(n1367), .B0(n819), .CI(n828), .CO(n816), .S0(n817)
         );
  HS65_LHS_XOR2X6 U2661 ( .A(n4683), .B(n2738), .Z(n1367) );
  HS65_LH_MX41X7 U2662 ( .D0(n2719), .S0(n1022), .D1(n4581), .S1(n4646), .D2(
        n4584), .S2(n4649), .D3(n4589), .S3(n4650), .Z(n2738) );
  HS65_LH_FA1X4 U2663 ( .A0(n1399), .B0(n817), .CI(n270), .CO(n269), .S0(
        product[20]) );
  HS65_LHS_XOR2X6 U2664 ( .A(n7), .B(n2699), .Z(n1399) );
  HS65_LH_MX41X7 U2665 ( .D0(n4493), .S0(n1019), .D1(n4591), .S1(n4653), .D2(
        n4594), .S2(n4655), .D3(n4598), .S3(n4656), .Z(n2699) );
  HS65_LH_FA1X4 U2666 ( .A0(n1135), .B0(n707), .CI(n722), .CO(n704), .S0(n705)
         );
  HS65_LHS_XOR2X6 U2667 ( .A(n103), .B(n3025), .Z(n1135) );
  HS65_LH_MX41X7 U2668 ( .D0(n3019), .S0(n1035), .D1(n4507), .S1(n4621), .D2(
        n4510), .S2(n4623), .D3(n4516), .S3(n4624), .Z(n3025) );
  HS65_LH_FA1X4 U2669 ( .A0(n1168), .B0(n723), .CI(n738), .CO(n720), .S0(n721)
         );
  HS65_LHS_XOR2X6 U2670 ( .A(n4701), .B(n2984), .Z(n1168) );
  HS65_LH_MX41X7 U2671 ( .D0(n4523), .S0(n1033), .D1(n4526), .S1(n4628), .D2(
        n4518), .S2(n4625), .D3(n4521), .S3(n4626), .Z(n2984) );
  HS65_LH_FA1X4 U2672 ( .A0(n1201), .B0(n739), .CI(n752), .CO(n736), .S0(n737)
         );
  HS65_LHS_XOR2X6 U2673 ( .A(n4698), .B(n2943), .Z(n1201) );
  HS65_LH_MX41X7 U2674 ( .D0(n4534), .S0(n1031), .D1(n4528), .S1(n4629), .D2(
        n4531), .S2(n4631), .D3(n4537), .S3(n4632), .Z(n2943) );
  HS65_LH_FA1X4 U2675 ( .A0(n1234), .B0(n753), .CI(n766), .CO(n750), .S0(n751)
         );
  HS65_LHS_XOR2X6 U2676 ( .A(n4695), .B(n2902), .Z(n1234) );
  HS65_LH_MX41X7 U2677 ( .D0(n4545), .S0(n1029), .D1(n4539), .S1(n4633), .D2(
        n4543), .S2(n4635), .D3(n4548), .S3(n4636), .Z(n2902) );
  HS65_LH_FA1X4 U2678 ( .A0(n1267), .B0(n767), .CI(n780), .CO(n764), .S0(n765)
         );
  HS65_LHS_XOR2X6 U2679 ( .A(n4692), .B(n2861), .Z(n1267) );
  HS65_LH_MX41X7 U2680 ( .D0(n2847), .S0(n1027), .D1(n4551), .S1(n4637), .D2(
        n4554), .S2(n4639), .D3(n4559), .S3(n4640), .Z(n2861) );
  HS65_LH_FA1X4 U2681 ( .A0(n1300), .B0(n781), .CI(n792), .CO(n778), .S0(n779)
         );
  HS65_LHS_XOR2X6 U2682 ( .A(n4689), .B(n2820), .Z(n1300) );
  HS65_LH_MX41X7 U2683 ( .D0(n2804), .S0(n1025), .D1(n4612), .S1(n4644), .D2(
        n4565), .S2(n4643), .D3(n4562), .S3(n4640), .Z(n2820) );
  HS65_LH_FA1X4 U2684 ( .A0(n1333), .B0(n793), .CI(n804), .CO(n790), .S0(n791)
         );
  HS65_LHS_XOR2X6 U2685 ( .A(n4686), .B(n2780), .Z(n1333) );
  HS65_LH_MX41X7 U2686 ( .D0(n2762), .S0(n1023), .D1(n4570), .S1(n4645), .D2(
        n4573), .S2(n4647), .D3(n4578), .S3(n4648), .Z(n2780) );
  HS65_LH_FA1X4 U2687 ( .A0(n1366), .B0(n805), .CI(n816), .CO(n802), .S0(n803)
         );
  HS65_LHS_XOR2X6 U2688 ( .A(n4683), .B(n2739), .Z(n1366) );
  HS65_LH_MX41X7 U2689 ( .D0(n2719), .S0(n1021), .D1(n4581), .S1(n4649), .D2(
        n4584), .S2(n4651), .D3(n4589), .S3(n4652), .Z(n2739) );
  HS65_LH_FA1X4 U2690 ( .A0(n1398), .B0(n803), .CI(n269), .CO(n268), .S0(
        product[21]) );
  HS65_LHS_XOR2X6 U2691 ( .A(n4681), .B(n2700), .Z(n1398) );
  HS65_LH_MX41X7 U2692 ( .D0(n1018), .S0(n4494), .D1(n4591), .S1(n4655), .D2(
        n4594), .S2(n4657), .D3(n4658), .S3(n4599), .Z(n2700) );
  HS65_LH_FA1X4 U2693 ( .A0(n1101), .B0(n1069), .CI(n688), .CO(n670), .S0(n671) );
  HS65_LH_AO22X9 U2694 ( .A(n4606), .B(n4617), .C(n4490), .D(n4617), .Z(n1069)
         );
  HS65_LHS_XOR2X6 U2695 ( .A(n115), .B(n3067), .Z(n1101) );
  HS65_LH_MX41X7 U2696 ( .D0(n3062), .S0(n1036), .D1(n4496), .S1(n4618), .D2(
        n4500), .S2(n4621), .D3(n4505), .S3(n4622), .Z(n3067) );
  HS65_LH_FA1X4 U2697 ( .A0(n1134), .B0(n689), .CI(n704), .CO(n686), .S0(n687)
         );
  HS65_LHS_XOR2X6 U2698 ( .A(n4704), .B(n3026), .Z(n1134) );
  HS65_LH_MX41X7 U2699 ( .D0(n3019), .S0(n1034), .D1(n4506), .S1(n4623), .D2(
        n4511), .S2(n4625), .D3(n4516), .S3(n4626), .Z(n3026) );
  HS65_LH_FA1X4 U2700 ( .A0(n1167), .B0(n705), .CI(n720), .CO(n702), .S0(n703)
         );
  HS65_LHS_XOR2X6 U2701 ( .A(n4701), .B(n2985), .Z(n1167) );
  HS65_LH_MX41X7 U2702 ( .D0(n4523), .S0(n1032), .D1(n4526), .S1(n4631), .D2(
        n4518), .S2(n4627), .D3(n4521), .S3(n4628), .Z(n2985) );
  HS65_LH_FA1X4 U2703 ( .A0(n1200), .B0(n721), .CI(n736), .CO(n718), .S0(n719)
         );
  HS65_LHS_XOR2X6 U2704 ( .A(n4697), .B(n2944), .Z(n1200) );
  HS65_LH_MX41X7 U2705 ( .D0(n4534), .S0(n1030), .D1(n4528), .S1(n4630), .D2(
        n4531), .S2(n4633), .D3(n4537), .S3(n4634), .Z(n2944) );
  HS65_LH_FA1X4 U2706 ( .A0(n1233), .B0(n737), .CI(n750), .CO(n734), .S0(n735)
         );
  HS65_LHS_XOR2X6 U2707 ( .A(n4695), .B(n2903), .Z(n1233) );
  HS65_LH_MX41X7 U2708 ( .D0(n4545), .S0(n1028), .D1(n4539), .S1(n4635), .D2(
        n4542), .S2(n4637), .D3(n4548), .S3(n4638), .Z(n2903) );
  HS65_LH_FA1X4 U2709 ( .A0(n1266), .B0(n751), .CI(n764), .CO(n748), .S0(n749)
         );
  HS65_LHS_XOR2X6 U2710 ( .A(n4692), .B(n2862), .Z(n1266) );
  HS65_LH_MX41X7 U2711 ( .D0(n2847), .S0(n1026), .D1(n4551), .S1(n4639), .D2(
        n4554), .S2(n4641), .D3(n4559), .S3(n4642), .Z(n2862) );
  HS65_LH_FA1X4 U2712 ( .A0(n1299), .B0(n765), .CI(n778), .CO(n762), .S0(n763)
         );
  HS65_LHS_XOR2X6 U2713 ( .A(n4689), .B(n2821), .Z(n1299) );
  HS65_LH_MX41X7 U2714 ( .D0(n4567), .S0(n1024), .D1(n4566), .S1(n4645), .D2(
        n4611), .S2(n4647), .D3(n4561), .S3(n4642), .Z(n2821) );
  HS65_LH_FA1X4 U2715 ( .A0(n1332), .B0(n779), .CI(n790), .CO(n776), .S0(n777)
         );
  HS65_LHS_XOR2X6 U2716 ( .A(n4686), .B(n2781), .Z(n1332) );
  HS65_LH_MX41X7 U2717 ( .D0(n2762), .S0(n1022), .D1(n4570), .S1(n4647), .D2(
        n4573), .S2(n4649), .D3(n4578), .S3(n4650), .Z(n2781) );
  HS65_LH_FA1X4 U2718 ( .A0(n1365), .B0(n791), .CI(n802), .CO(n788), .S0(n789)
         );
  HS65_LHS_XOR2X6 U2719 ( .A(n4683), .B(n2740), .Z(n1365) );
  HS65_LH_MX41X7 U2720 ( .D0(n2719), .S0(n1020), .D1(n4581), .S1(n4651), .D2(
        n4584), .S2(n4653), .D3(n4589), .S3(n4654), .Z(n2740) );
  HS65_LH_FA1X4 U2721 ( .A0(n1397), .B0(n789), .CI(n268), .CO(n267), .S0(
        product[22]) );
  HS65_LHS_XOR2X6 U2722 ( .A(n7), .B(n2701), .Z(n1397) );
  HS65_LH_MX41X7 U2723 ( .D0(n1017), .S0(n4494), .D1(n4591), .S1(n4656), .D2(
        n4658), .S2(n4596), .D3(n4660), .S3(n4600), .Z(n2701) );
  HS65_LH_FA1X4 U2724 ( .A0(n1100), .B0(n1068), .CI(n670), .CO(n652), .S0(n653) );
  HS65_LH_AO222X4 U2725 ( .A(n4608), .B(n4619), .C(n4602), .D(n4617), .E(n4490), .F(n1038), .Z(n1068) );
  HS65_LHS_XOR2X6 U2726 ( .A(n4706), .B(n3068), .Z(n1100) );
  HS65_LH_MX41X7 U2727 ( .D0(n3062), .S0(n1035), .D1(n4496), .S1(n4620), .D2(
        n4499), .S2(n4623), .D3(n4505), .S3(n4624), .Z(n3068) );
  HS65_LH_FA1X4 U2728 ( .A0(n1133), .B0(n671), .CI(n686), .CO(n668), .S0(n669)
         );
  HS65_LHS_XOR2X6 U2729 ( .A(n4704), .B(n3027), .Z(n1133) );
  HS65_LH_MX41X7 U2730 ( .D0(n3019), .S0(n1033), .D1(n4507), .S1(n4625), .D2(
        n4510), .S2(n4627), .D3(n4515), .S3(n4628), .Z(n3027) );
  HS65_LH_FA1X4 U2731 ( .A0(n1166), .B0(n687), .CI(n702), .CO(n684), .S0(n685)
         );
  HS65_LHS_XOR2X6 U2732 ( .A(n4701), .B(n2986), .Z(n1166) );
  HS65_LH_MX41X7 U2733 ( .D0(n4523), .S0(n1031), .D1(n4526), .S1(n4633), .D2(
        n4517), .S2(n4629), .D3(n4521), .S3(n4630), .Z(n2986) );
  HS65_LH_FA1X4 U2734 ( .A0(n1199), .B0(n703), .CI(n718), .CO(n700), .S0(n701)
         );
  HS65_LHS_XOR2X6 U2735 ( .A(n4697), .B(n2945), .Z(n1199) );
  HS65_LH_MX41X7 U2736 ( .D0(n4534), .S0(n1029), .D1(n4528), .S1(n4632), .D2(
        n4531), .S2(n4635), .D3(n4536), .S3(n4636), .Z(n2945) );
  HS65_LH_FA1X4 U2737 ( .A0(n1232), .B0(n719), .CI(n734), .CO(n716), .S0(n717)
         );
  HS65_LHS_XOR2X6 U2738 ( .A(n4694), .B(n2904), .Z(n1232) );
  HS65_LH_MX41X7 U2739 ( .D0(n2890), .S0(n1027), .D1(n4540), .S1(n4637), .D2(
        n4543), .S2(n4639), .D3(n4549), .S3(n4640), .Z(n2904) );
  HS65_LH_FA1X4 U2740 ( .A0(n1265), .B0(n735), .CI(n748), .CO(n732), .S0(n733)
         );
  HS65_LHS_XOR2X6 U2741 ( .A(n4692), .B(n2863), .Z(n1265) );
  HS65_LH_MX41X7 U2742 ( .D0(n2847), .S0(n1025), .D1(n4551), .S1(n4641), .D2(
        n4554), .S2(n4643), .D3(n4559), .S3(n4644), .Z(n2863) );
  HS65_LH_FA1X4 U2743 ( .A0(n1298), .B0(n749), .CI(n762), .CO(n746), .S0(n747)
         );
  HS65_LHS_XOR2X6 U2744 ( .A(n4688), .B(n2822), .Z(n1298) );
  HS65_LH_MX41X7 U2745 ( .D0(n4567), .S0(n1023), .D1(n4566), .S1(n4646), .D2(
        n4611), .S2(n4649), .D3(n4561), .S3(n4644), .Z(n2822) );
  HS65_LH_FA1X4 U2746 ( .A0(n1331), .B0(n763), .CI(n776), .CO(n760), .S0(n761)
         );
  HS65_LHS_XOR2X6 U2747 ( .A(n4686), .B(n2782), .Z(n1331) );
  HS65_LH_MX41X7 U2748 ( .D0(n4575), .S0(n1021), .D1(n4570), .S1(n4649), .D2(
        n4573), .S2(n4651), .D3(n4578), .S3(n4652), .Z(n2782) );
  HS65_LH_FA1X4 U2749 ( .A0(n1364), .B0(n777), .CI(n788), .CO(n774), .S0(n775)
         );
  HS65_LHS_XOR2X6 U2750 ( .A(n4683), .B(n2741), .Z(n1364) );
  HS65_LH_MX41X7 U2751 ( .D0(n4586), .S0(n1019), .D1(n4581), .S1(n4652), .D2(
        n4584), .S2(n4655), .D3(n4589), .S3(n4656), .Z(n2741) );
  HS65_LH_FA1X4 U2752 ( .A0(n1396), .B0(n775), .CI(n267), .CO(n266), .S0(
        product[23]) );
  HS65_LHS_XOR2X6 U2753 ( .A(n7), .B(n2702), .Z(n1396) );
  HS65_LH_MX41X7 U2754 ( .D0(n1016), .S0(n4494), .D1(n4658), .S1(n4592), .D2(
        n4660), .S2(n4596), .D3(n4662), .S3(n4600), .Z(n2702) );
  HS65_LH_FA1X4 U2755 ( .A0(n1099), .B0(n1067), .CI(n652), .CO(n634), .S0(n635) );
  HS65_LH_MX41X7 U2756 ( .D0(n1037), .S0(n4492), .D1(n4620), .S1(n4608), .D2(
        n4618), .S2(n4604), .D3(n4616), .S3(n4609), .Z(n1067) );
  HS65_LHS_XOR2X6 U2757 ( .A(n4707), .B(n3069), .Z(n1099) );
  HS65_LH_MX41X7 U2758 ( .D0(n3062), .S0(n1034), .D1(n4496), .S1(n4622), .D2(
        n4499), .S2(n4625), .D3(n4505), .S3(n4626), .Z(n3069) );
  HS65_LH_FA1X4 U2759 ( .A0(n1132), .B0(n653), .CI(n668), .CO(n650), .S0(n651)
         );
  HS65_LHS_XOR2X6 U2760 ( .A(n4704), .B(n3028), .Z(n1132) );
  HS65_LH_MX41X7 U2761 ( .D0(n3019), .S0(n1032), .D1(n4507), .S1(n4626), .D2(
        n4510), .S2(n4629), .D3(n4515), .S3(n4630), .Z(n3028) );
  HS65_LH_FA1X4 U2762 ( .A0(n1165), .B0(n669), .CI(n684), .CO(n666), .S0(n667)
         );
  HS65_LHS_XOR2X6 U2763 ( .A(n4701), .B(n2987), .Z(n1165) );
  HS65_LH_MX41X7 U2764 ( .D0(n4523), .S0(n1030), .D1(n4526), .S1(n4634), .D2(
        n4517), .S2(n4631), .D3(n4521), .S3(n4632), .Z(n2987) );
  HS65_LH_FA1X4 U2765 ( .A0(n1198), .B0(n685), .CI(n700), .CO(n682), .S0(n683)
         );
  HS65_LHS_XOR2X6 U2766 ( .A(n4697), .B(n2946), .Z(n1198) );
  HS65_LH_MX41X7 U2767 ( .D0(n4534), .S0(n1028), .D1(n4528), .S1(n4634), .D2(
        n4531), .S2(n4637), .D3(n4536), .S3(n4638), .Z(n2946) );
  HS65_LH_FA1X4 U2768 ( .A0(n1231), .B0(n701), .CI(n716), .CO(n698), .S0(n699)
         );
  HS65_LHS_XOR2X6 U2769 ( .A(n4695), .B(n2905), .Z(n1231) );
  HS65_LH_MX41X7 U2770 ( .D0(n2890), .S0(n1026), .D1(n4540), .S1(n4638), .D2(
        n4543), .S2(n4641), .D3(n4548), .S3(n4642), .Z(n2905) );
  HS65_LH_FA1X4 U2771 ( .A0(n1264), .B0(n717), .CI(n732), .CO(n714), .S0(n715)
         );
  HS65_LHS_XOR2X6 U2772 ( .A(n4692), .B(n2864), .Z(n1264) );
  HS65_LH_MX41X7 U2773 ( .D0(n4556), .S0(n1024), .D1(n4550), .S1(n4643), .D2(
        n4553), .S2(n4645), .D3(n4558), .S3(n4646), .Z(n2864) );
  HS65_LH_FA1X4 U2774 ( .A0(n1297), .B0(n733), .CI(n746), .CO(n730), .S0(n731)
         );
  HS65_LHS_XOR2X6 U2775 ( .A(n4688), .B(n2823), .Z(n1297) );
  HS65_LH_MX41X7 U2776 ( .D0(n4567), .S0(n1022), .D1(n4611), .S1(n4651), .D2(
        n4564), .S2(n4649), .D3(n4561), .S3(n4646), .Z(n2823) );
  HS65_LH_FA1X4 U2777 ( .A0(n1330), .B0(n747), .CI(n760), .CO(n744), .S0(n745)
         );
  HS65_LHS_XOR2X6 U2778 ( .A(n4686), .B(n2783), .Z(n1330) );
  HS65_LH_MX41X7 U2779 ( .D0(n4575), .S0(n1020), .D1(n4570), .S1(n4651), .D2(
        n4573), .S2(n4653), .D3(n4578), .S3(n4654), .Z(n2783) );
  HS65_LH_FA1X4 U2780 ( .A0(n1363), .B0(n761), .CI(n774), .CO(n758), .S0(n759)
         );
  HS65_LHS_XOR2X6 U2781 ( .A(n4683), .B(n2742), .Z(n1363) );
  HS65_LH_MX41X7 U2782 ( .D0(n4586), .S0(n1018), .D1(n4580), .S1(n4654), .D2(
        n4583), .S2(n4657), .D3(n4588), .S3(n4658), .Z(n2742) );
  HS65_LH_FA1X4 U2783 ( .A0(n1395), .B0(n759), .CI(n266), .CO(n265), .S0(
        product[24]) );
  HS65_LHS_XOR2X6 U2784 ( .A(n4681), .B(n2703), .Z(n1395) );
  HS65_LH_MX41X7 U2785 ( .D0(n1015), .S0(n4494), .D1(n4660), .S1(n4592), .D2(
        n4662), .S2(n4596), .D3(n4598), .S3(n4664), .Z(n2703) );
  HS65_LH_FA1X4 U2786 ( .A0(n1131), .B0(n635), .CI(n650), .CO(n632), .S0(n633)
         );
  HS65_LHS_XOR2X6 U2787 ( .A(n4704), .B(n3029), .Z(n1131) );
  HS65_LH_MX41X7 U2788 ( .D0(n3019), .S0(n1031), .D1(n4507), .S1(n4629), .D2(
        n4510), .S2(n4631), .D3(n4515), .S3(n4632), .Z(n3029) );
  HS65_LH_FA1X4 U2789 ( .A0(n1164), .B0(n651), .CI(n666), .CO(n648), .S0(n649)
         );
  HS65_LHS_XOR2X6 U2790 ( .A(n4701), .B(n2988), .Z(n1164) );
  HS65_LH_MX41X7 U2791 ( .D0(n4523), .S0(n1029), .D1(n4526), .S1(n4636), .D2(
        n4517), .S2(n4633), .D3(n4520), .S3(n4634), .Z(n2988) );
  HS65_LH_FA1X4 U2792 ( .A0(n1197), .B0(n667), .CI(n682), .CO(n664), .S0(n665)
         );
  HS65_LHS_XOR2X6 U2793 ( .A(n4698), .B(n2947), .Z(n1197) );
  HS65_LH_MX41X7 U2794 ( .D0(n2933), .S0(n1027), .D1(n4529), .S1(n4636), .D2(
        n4532), .S2(n4639), .D3(n4537), .S3(n4640), .Z(n2947) );
  HS65_LH_FA1X4 U2795 ( .A0(n1230), .B0(n683), .CI(n698), .CO(n680), .S0(n681)
         );
  HS65_LHS_XOR2X6 U2796 ( .A(n4695), .B(n2906), .Z(n1230) );
  HS65_LH_MX41X7 U2797 ( .D0(n2890), .S0(n1025), .D1(n4540), .S1(n4641), .D2(
        n4543), .S2(n4643), .D3(n4548), .S3(n4644), .Z(n2906) );
  HS65_LH_FA1X4 U2798 ( .A0(n1263), .B0(n699), .CI(n714), .CO(n696), .S0(n697)
         );
  HS65_LHS_XOR2X6 U2799 ( .A(n4692), .B(n2865), .Z(n1263) );
  HS65_LH_MX41X7 U2800 ( .D0(n2847), .S0(n1023), .D1(n4551), .S1(n4645), .D2(
        n4554), .S2(n4647), .D3(n4559), .S3(n4648), .Z(n2865) );
  HS65_LH_FA1X4 U2801 ( .A0(n1296), .B0(n715), .CI(n730), .CO(n712), .S0(n713)
         );
  HS65_LHS_XOR2X6 U2802 ( .A(n4689), .B(n2824), .Z(n1296) );
  HS65_LH_MX41X7 U2803 ( .D0(n2804), .S0(n1021), .D1(n4612), .S1(n4653), .D2(
        n4565), .S2(n4651), .D3(n4562), .S3(n4648), .Z(n2824) );
  HS65_LH_FA1X4 U2804 ( .A0(n1329), .B0(n731), .CI(n744), .CO(n728), .S0(n729)
         );
  HS65_LHS_XOR2X6 U2805 ( .A(n4686), .B(n2784), .Z(n1329) );
  HS65_LH_MX41X7 U2806 ( .D0(n4575), .S0(n1019), .D1(n4570), .S1(n4652), .D2(
        n4573), .S2(n4655), .D3(n4578), .S3(n4656), .Z(n2784) );
  HS65_LH_FA1X4 U2807 ( .A0(n1362), .B0(n745), .CI(n758), .CO(n742), .S0(n743)
         );
  HS65_LHS_XOR2X6 U2808 ( .A(n4683), .B(n2743), .Z(n1362) );
  HS65_LH_MX41X7 U2809 ( .D0(n4586), .S0(n1017), .D1(n4581), .S1(n4656), .D2(
        n4584), .S2(n4659), .D3(n4589), .S3(n4660), .Z(n2743) );
  HS65_LH_FA1X4 U2810 ( .A0(n1394), .B0(n743), .CI(n265), .CO(n264), .S0(
        product[25]) );
  HS65_LHS_XOR2X6 U2811 ( .A(n7), .B(n2704), .Z(n1394) );
  HS65_LH_MX41X7 U2812 ( .D0(n1014), .S0(n4494), .D1(n4662), .S1(n4592), .D2(
        n4594), .S2(n4665), .D3(n4598), .S3(n4666), .Z(n2704) );
  HS65_LH_FA1X4 U2813 ( .A0(n1163), .B0(n633), .CI(n648), .CO(n630), .S0(n631)
         );
  HS65_LHS_XOR2X6 U2814 ( .A(n4701), .B(n2989), .Z(n1163) );
  HS65_LH_MX41X7 U2815 ( .D0(n2976), .S0(n1028), .D1(n4526), .S1(n4639), .D2(
        n4518), .S2(n4635), .D3(n4521), .S3(n4636), .Z(n2989) );
  HS65_LH_FA1X4 U2816 ( .A0(n1196), .B0(n649), .CI(n664), .CO(n646), .S0(n647)
         );
  HS65_LHS_XOR2X6 U2817 ( .A(n4698), .B(n2948), .Z(n1196) );
  HS65_LH_MX41X7 U2818 ( .D0(n2933), .S0(n1026), .D1(n4529), .S1(n4639), .D2(
        n4532), .S2(n4641), .D3(n4537), .S3(n4642), .Z(n2948) );
  HS65_LH_FA1X4 U2819 ( .A0(n1229), .B0(n665), .CI(n680), .CO(n662), .S0(n663)
         );
  HS65_LHS_XOR2X6 U2820 ( .A(n4694), .B(n2907), .Z(n1229) );
  HS65_LH_MX41X7 U2821 ( .D0(n4545), .S0(n1024), .D1(n4539), .S1(n4643), .D2(
        n4542), .S2(n4645), .D3(n4547), .S3(n4646), .Z(n2907) );
  HS65_LH_FA1X4 U2822 ( .A0(n1262), .B0(n681), .CI(n696), .CO(n678), .S0(n679)
         );
  HS65_LHS_XOR2X6 U2823 ( .A(n4692), .B(n2866), .Z(n1262) );
  HS65_LH_MX41X7 U2824 ( .D0(n2847), .S0(n1022), .D1(n4551), .S1(n4647), .D2(
        n4554), .S2(n4649), .D3(n4559), .S3(n4650), .Z(n2866) );
  HS65_LH_FA1X4 U2825 ( .A0(n1295), .B0(n697), .CI(n712), .CO(n694), .S0(n695)
         );
  HS65_LHS_XOR2X6 U2826 ( .A(n4689), .B(n2825), .Z(n1295) );
  HS65_LH_MX41X7 U2827 ( .D0(n2804), .S0(n1020), .D1(n4612), .S1(n4654), .D2(
        n4565), .S2(n4653), .D3(n4562), .S3(n4650), .Z(n2825) );
  HS65_LH_FA1X4 U2828 ( .A0(n1328), .B0(n713), .CI(n728), .CO(n710), .S0(n711)
         );
  HS65_LHS_XOR2X6 U2829 ( .A(n4685), .B(n2785), .Z(n1328) );
  HS65_LH_MX41X7 U2830 ( .D0(n4575), .S0(n1018), .D1(n4569), .S1(n4655), .D2(
        n4572), .S2(n4657), .D3(n4577), .S3(n4658), .Z(n2785) );
  HS65_LH_FA1X4 U2831 ( .A0(n1361), .B0(n729), .CI(n742), .CO(n726), .S0(n727)
         );
  HS65_LHS_XOR2X6 U2832 ( .A(n4683), .B(n2744), .Z(n1361) );
  HS65_LH_MX41X7 U2833 ( .D0(n4586), .S0(n1016), .D1(n4581), .S1(n4659), .D2(
        n4584), .S2(n4661), .D3(n4589), .S3(n4662), .Z(n2744) );
  HS65_LH_FA1X4 U2834 ( .A0(n1393), .B0(n727), .CI(n264), .CO(n263), .S0(
        product[26]) );
  HS65_LHS_XOR2X6 U2835 ( .A(n4680), .B(n2705), .Z(n1393) );
  HS65_LH_MX41X7 U2836 ( .D0(n4493), .S0(n1013), .D1(n4591), .S1(n4665), .D2(
        n4594), .S2(n4667), .D3(n4598), .S3(n4668), .Z(n2705) );
  HS65_LH_FA1X4 U2837 ( .A0(n1195), .B0(n631), .CI(n646), .CO(n628), .S0(n629)
         );
  HS65_LHS_XOR2X6 U2838 ( .A(n4698), .B(n2949), .Z(n1195) );
  HS65_LH_MX41X7 U2839 ( .D0(n4534), .S0(n1025), .D1(n4529), .S1(n4640), .D2(
        n4532), .S2(n4643), .D3(n4537), .S3(n4644), .Z(n2949) );
  HS65_LH_FA1X4 U2840 ( .A0(n1228), .B0(n647), .CI(n662), .CO(n644), .S0(n645)
         );
  HS65_LHS_XOR2X6 U2841 ( .A(n4695), .B(n2908), .Z(n1228) );
  HS65_LH_MX41X7 U2842 ( .D0(n2890), .S0(n1023), .D1(n4540), .S1(n4645), .D2(
        n4543), .S2(n4647), .D3(n4548), .S3(n4648), .Z(n2908) );
  HS65_LH_FA1X4 U2843 ( .A0(n1261), .B0(n663), .CI(n678), .CO(n660), .S0(n661)
         );
  HS65_LHS_XOR2X6 U2844 ( .A(n4692), .B(n2867), .Z(n1261) );
  HS65_LH_MX41X7 U2845 ( .D0(n2847), .S0(n1021), .D1(n4551), .S1(n4649), .D2(
        n4554), .S2(n4651), .D3(n4559), .S3(n4652), .Z(n2867) );
  HS65_LH_FA1X4 U2846 ( .A0(n1294), .B0(n679), .CI(n694), .CO(n676), .S0(n677)
         );
  HS65_LHS_XOR2X6 U2847 ( .A(n4689), .B(n2826), .Z(n1294) );
  HS65_LH_MX41X7 U2848 ( .D0(n2804), .S0(n1019), .D1(n4612), .S1(n4657), .D2(
        n4565), .S2(n4655), .D3(n4562), .S3(n4652), .Z(n2826) );
  HS65_LH_FA1X4 U2849 ( .A0(n1327), .B0(n695), .CI(n710), .CO(n692), .S0(n693)
         );
  HS65_LHS_XOR2X6 U2850 ( .A(n4686), .B(n2786), .Z(n1327) );
  HS65_LH_MX41X7 U2851 ( .D0(n4575), .S0(n1017), .D1(n4569), .S1(n4657), .D2(
        n4573), .S2(n4659), .D3(n4578), .S3(n4660), .Z(n2786) );
  HS65_LH_FA1X4 U2852 ( .A0(n1360), .B0(n711), .CI(n726), .CO(n708), .S0(n709)
         );
  HS65_LHS_XOR2X6 U2853 ( .A(n19), .B(n2745), .Z(n1360) );
  HS65_LH_MX41X7 U2854 ( .D0(n4586), .S0(n1015), .D1(n4580), .S1(n4661), .D2(
        n4583), .S2(n4663), .D3(n4588), .S3(n4664), .Z(n2745) );
  HS65_LH_FA1X4 U2855 ( .A0(n1392), .B0(n709), .CI(n263), .CO(n262), .S0(
        product[27]) );
  HS65_LHS_XOR2X6 U2856 ( .A(n4681), .B(n2706), .Z(n1392) );
  HS65_LH_MX41X7 U2857 ( .D0(n1012), .S0(n4494), .D1(n4591), .S1(n4667), .D2(
        n4594), .S2(n4669), .D3(n4670), .S3(n4600), .Z(n2706) );
  HS65_LH_FA1X4 U2858 ( .A0(n1227), .B0(n629), .CI(n644), .CO(n626), .S0(n627)
         );
  HS65_LHS_XOR2X6 U2859 ( .A(n4695), .B(n2909), .Z(n1227) );
  HS65_LH_MX41X7 U2860 ( .D0(n2890), .S0(n1022), .D1(n4540), .S1(n4646), .D2(
        n4543), .S2(n4649), .D3(n4548), .S3(n4650), .Z(n2909) );
  HS65_LH_FA1X4 U2861 ( .A0(n1260), .B0(n645), .CI(n660), .CO(n642), .S0(n643)
         );
  HS65_LHS_XOR2X6 U2862 ( .A(n4692), .B(n2868), .Z(n1260) );
  HS65_LH_MX41X7 U2863 ( .D0(n4556), .S0(n1020), .D1(n4551), .S1(n4651), .D2(
        n4554), .S2(n4653), .D3(n4559), .S3(n4654), .Z(n2868) );
  HS65_LH_FA1X4 U2864 ( .A0(n1293), .B0(n661), .CI(n676), .CO(n658), .S0(n659)
         );
  HS65_LHS_XOR2X6 U2865 ( .A(n4689), .B(n2827), .Z(n1293) );
  HS65_LH_MX41X7 U2866 ( .D0(n4567), .S0(n1018), .D1(n4612), .S1(n4658), .D2(
        n4565), .S2(n4657), .D3(n4562), .S3(n4654), .Z(n2827) );
  HS65_LH_FA1X4 U2867 ( .A0(n1326), .B0(n677), .CI(n692), .CO(n674), .S0(n675)
         );
  HS65_LHS_XOR2X6 U2868 ( .A(n4686), .B(n2787), .Z(n1326) );
  HS65_LH_MX41X7 U2869 ( .D0(n4575), .S0(n1016), .D1(n4569), .S1(n4659), .D2(
        n4572), .S2(n4661), .D3(n4578), .S3(n4662), .Z(n2787) );
  HS65_LH_FA1X4 U2870 ( .A0(n1359), .B0(n693), .CI(n708), .CO(n690), .S0(n691)
         );
  HS65_LHS_XOR2X6 U2871 ( .A(n4683), .B(n2746), .Z(n1359) );
  HS65_LH_MX41X7 U2872 ( .D0(n4586), .S0(n1014), .D1(n4580), .S1(n4662), .D2(
        n4583), .S2(n4665), .D3(n4588), .S3(n4666), .Z(n2746) );
  HS65_LH_FA1X4 U2873 ( .A0(n1391), .B0(n691), .CI(n262), .CO(n261), .S0(
        product[28]) );
  HS65_LHS_XOR2X6 U2874 ( .A(n4681), .B(n2707), .Z(n1391) );
  HS65_LH_MX41X7 U2875 ( .D0(n1011), .S0(n4494), .D1(n4591), .S1(n4669), .D2(
        n4670), .S2(n4595), .D3(n4672), .S3(n4599), .Z(n2707) );
  HS65_LH_FA1X4 U2876 ( .A0(n1259), .B0(n627), .CI(n642), .CO(n624), .S0(n625)
         );
  HS65_LHS_XOR2X6 U2877 ( .A(n4692), .B(n2869), .Z(n1259) );
  HS65_LH_MX41X7 U2878 ( .D0(n4556), .S0(n1019), .D1(n4551), .S1(n4652), .D2(
        n4554), .S2(n4655), .D3(n4559), .S3(n4656), .Z(n2869) );
  HS65_LH_FA1X4 U2879 ( .A0(n1292), .B0(n643), .CI(n658), .CO(n640), .S0(n641)
         );
  HS65_LHS_XOR2X6 U2880 ( .A(n4689), .B(n2828), .Z(n1292) );
  HS65_LH_MX41X7 U2881 ( .D0(n4567), .S0(n1017), .D1(n4612), .S1(n4660), .D2(
        n4565), .S2(n4659), .D3(n4562), .S3(n4656), .Z(n2828) );
  HS65_LH_FA1X4 U2882 ( .A0(n1325), .B0(n659), .CI(n674), .CO(n656), .S0(n657)
         );
  HS65_LHS_XOR2X6 U2883 ( .A(n4685), .B(n2788), .Z(n1325) );
  HS65_LH_MX41X7 U2884 ( .D0(n4575), .S0(n1015), .D1(n4569), .S1(n4661), .D2(
        n4572), .S2(n4663), .D3(n4577), .S3(n4664), .Z(n2788) );
  HS65_LH_FA1X4 U2885 ( .A0(n1358), .B0(n675), .CI(n690), .CO(n672), .S0(n673)
         );
  HS65_LHS_XOR2X6 U2886 ( .A(n19), .B(n2747), .Z(n1358) );
  HS65_LH_MX41X7 U2887 ( .D0(n4586), .S0(n1013), .D1(n4580), .S1(n4664), .D2(
        n4584), .S2(n4667), .D3(n4589), .S3(n4668), .Z(n2747) );
  HS65_LH_FA1X4 U2888 ( .A0(n1390), .B0(n673), .CI(n261), .CO(n260), .S0(
        product[29]) );
  HS65_LHS_XOR2X6 U2889 ( .A(n7), .B(n2708), .Z(n1390) );
  HS65_LH_MX41X7 U2890 ( .D0(n1010), .S0(n4494), .D1(n4670), .S1(n4592), .D2(
        n4672), .S2(n4595), .D3(n4674), .S3(n4600), .Z(n2708) );
  HS65_LH_FA1X4 U2891 ( .A0(n1291), .B0(n625), .CI(n640), .CO(n622), .S0(n623)
         );
  HS65_LHS_XOR2X6 U2892 ( .A(n4689), .B(n2829), .Z(n1291) );
  HS65_LH_MX41X7 U2893 ( .D0(n4567), .S0(n1016), .D1(n4612), .S1(n4663), .D2(
        n4564), .S2(n4661), .D3(n4562), .S3(n4658), .Z(n2829) );
  HS65_LH_FA1X4 U2894 ( .A0(n1324), .B0(n641), .CI(n656), .CO(n638), .S0(n639)
         );
  HS65_LHS_XOR2X6 U2895 ( .A(n4685), .B(n2789), .Z(n1324) );
  HS65_LH_MX41X7 U2896 ( .D0(n4575), .S0(n1014), .D1(n4569), .S1(n4662), .D2(
        n4572), .S2(n4665), .D3(n4577), .S3(n4666), .Z(n2789) );
  HS65_LH_FA1X4 U2897 ( .A0(n1357), .B0(n657), .CI(n672), .CO(n654), .S0(n655)
         );
  HS65_LHS_XOR2X6 U2898 ( .A(n4683), .B(n2748), .Z(n1357) );
  HS65_LH_MX41X7 U2899 ( .D0(n4586), .S0(n1012), .D1(n4580), .S1(n4667), .D2(
        n4584), .S2(n4669), .D3(n4589), .S3(n4670), .Z(n2748) );
  HS65_LH_FA1X4 U2900 ( .A0(n1389), .B0(n655), .CI(n260), .CO(n259), .S0(
        product[30]) );
  HS65_LHS_XOR2X6 U2901 ( .A(n4681), .B(n2709), .Z(n1389) );
  HS65_LH_MX41X7 U2902 ( .D0(n1009), .S0(n4494), .D1(n4672), .S1(n4592), .D2(
        n4674), .S2(n4595), .D3(n4676), .S3(n4599), .Z(n2709) );
  HS65_LH_FA1X4 U2903 ( .A0(n1323), .B0(n623), .CI(n638), .CO(n620), .S0(n621)
         );
  HS65_LHS_XOR2X6 U2904 ( .A(n4685), .B(n2790), .Z(n1323) );
  HS65_LH_MX41X7 U2905 ( .D0(n4575), .S0(n1013), .D1(n4569), .S1(n4664), .D2(
        n4573), .S2(n4667), .D3(n4578), .S3(n4668), .Z(n2790) );
  HS65_LH_FA1X4 U2906 ( .A0(n1356), .B0(n639), .CI(n654), .CO(n636), .S0(n637)
         );
  HS65_LHS_XOR2X6 U2907 ( .A(n4683), .B(n2749), .Z(n1356) );
  HS65_LH_MX41X7 U2908 ( .D0(n4586), .S0(n1011), .D1(n4580), .S1(n4669), .D2(
        n4583), .S2(n4671), .D3(n4589), .S3(n4672), .Z(n2749) );
  HS65_LH_FA1X4 U2909 ( .A0(n1388), .B0(n637), .CI(n259), .CO(n258), .S0(
        product[31]) );
  HS65_LHS_XOR2X6 U2910 ( .A(n4680), .B(n2710), .Z(n1388) );
  HS65_LH_MX41X7 U2911 ( .D0(n1008), .S0(n4493), .D1(n4674), .S1(n4591), .D2(
        n4676), .S2(n4594), .D3(n4598), .S3(n4678), .Z(n2710) );
  HS65_LH_FA1X4 U2912 ( .A0(n1355), .B0(n621), .CI(n636), .CO(n618), .S0(n619)
         );
  HS65_LHS_XOR2X6 U2913 ( .A(n19), .B(n2750), .Z(n1355) );
  HS65_LH_MX41X7 U2914 ( .D0(n4586), .S0(n1010), .D1(n4580), .S1(n4671), .D2(
        n4583), .S2(n4673), .D3(n4588), .S3(n4674), .Z(n2750) );
  HS65_LH_FA1X4 U2915 ( .A0(n1204), .B0(n787), .CI(n798), .CO(n784), .S0(n785)
         );
  HS65_LHS_XOR2X6 U2916 ( .A(n4698), .B(n2940), .Z(n1204) );
  HS65_LH_MX41X7 U2917 ( .D0(n2933), .S0(n1034), .D1(n4528), .S1(n4623), .D2(
        n4533), .S2(n4625), .D3(n4538), .S3(n4626), .Z(n2940) );
  HS65_LH_FA1X4 U2918 ( .A0(n599), .B0(n616), .CI(n1129), .CO(n596), .S0(n597)
         );
  HS65_LHS_XOR2X6 U2919 ( .A(n4704), .B(n3031), .Z(n1129) );
  HS65_LH_MX41X7 U2920 ( .D0(n4512), .S0(n1029), .D1(n4506), .S1(n4632), .D2(
        n4510), .S2(n4635), .D3(n4515), .S3(n4636), .Z(n3031) );
  HS65_LH_FA1X4 U2921 ( .A0(n477), .B0(n491), .CI(n1122), .CO(n474), .S0(n475)
         );
  HS65_LHS_XOR2X6 U2922 ( .A(n4703), .B(n3038), .Z(n1122) );
  HS65_LH_MX41X7 U2923 ( .D0(n4512), .S0(n1022), .D1(n4506), .S1(n4647), .D2(
        n4509), .S2(n4649), .D3(n4514), .S3(n4650), .Z(n3038) );
  HS65_LH_FA1X4 U2924 ( .A0(n473), .B0(n487), .CI(n1186), .CO(n470), .S0(n471)
         );
  HS65_LHS_XOR2X6 U2925 ( .A(n4698), .B(n2958), .Z(n1186) );
  HS65_LH_MX41X7 U2926 ( .D0(n4534), .S0(n1016), .D1(n4528), .S1(n4659), .D2(
        n4531), .S2(n4661), .D3(n4536), .S3(n4662), .Z(n2958) );
  HS65_LH_FA1X4 U2927 ( .A0(n581), .B0(n1096), .CI(n596), .CO(n578), .S0(n579)
         );
  HS65_LHS_XOR2X6 U2928 ( .A(n4707), .B(n3072), .Z(n1096) );
  HS65_LH_MX41X7 U2929 ( .D0(n3062), .S0(n1031), .D1(n4496), .S1(n4629), .D2(
        n4499), .S2(n4631), .D3(n4504), .S3(n4632), .Z(n3072) );
  HS65_LH_FA1X4 U2930 ( .A0(n595), .B0(n612), .CI(n1193), .CO(n592), .S0(n593)
         );
  HS65_LHS_XOR2X6 U2931 ( .A(n4697), .B(n2951), .Z(n1193) );
  HS65_LH_MX41X7 U2932 ( .D0(n4534), .S0(n1023), .D1(n4528), .S1(n4644), .D2(
        n4531), .S2(n4647), .D3(n4536), .S3(n4648), .Z(n2951) );
  HS65_LH_FA1X4 U2933 ( .A0(n563), .B0(n1095), .CI(n578), .CO(n560), .S0(n561)
         );
  HS65_LHS_XOR2X6 U2934 ( .A(n4707), .B(n3073), .Z(n1095) );
  HS65_LH_MX41X7 U2935 ( .D0(n3062), .S0(n1030), .D1(n4496), .S1(n4630), .D2(
        n4499), .S2(n4633), .D3(n4504), .S3(n4634), .Z(n3073) );
  HS65_LH_FA1X4 U2936 ( .A0(n561), .B0(n1127), .CI(n1159), .CO(n558), .S0(n559) );
  HS65_LHS_XOR2X6 U2937 ( .A(n4700), .B(n2993), .Z(n1159) );
  HS65_LHS_XOR2X6 U2938 ( .A(n4704), .B(n3033), .Z(n1127) );
  HS65_LH_MX41X7 U2939 ( .D0(n4523), .S0(n1024), .D1(n4525), .S1(n4647), .D2(
        n4517), .S2(n4643), .D3(n4520), .S3(n4644), .Z(n2993) );
  HS65_LH_FA1X4 U2940 ( .A0(n591), .B0(n608), .CI(n1257), .CO(n588), .S0(n589)
         );
  HS65_LHS_XOR2X6 U2941 ( .A(n4691), .B(n2871), .Z(n1257) );
  HS65_LH_MX41X7 U2942 ( .D0(n4556), .S0(n1017), .D1(n4550), .S1(n4656), .D2(
        n4553), .S2(n4659), .D3(n4558), .S3(n4660), .Z(n2871) );
  HS65_LH_FA1X4 U2943 ( .A0(n589), .B0(n606), .CI(n1289), .CO(n586), .S0(n587)
         );
  HS65_LHS_XOR2X6 U2944 ( .A(n4688), .B(n2831), .Z(n1289) );
  HS65_LH_MX41X7 U2945 ( .D0(n4567), .S0(n1014), .D1(n4611), .S1(n4666), .D2(
        n4564), .S2(n4665), .D3(n4561), .S3(n4662), .Z(n2831) );
  HS65_LH_FA1X4 U2946 ( .A0(n587), .B0(n604), .CI(n1321), .CO(n584), .S0(n585)
         );
  HS65_LHS_XOR2X6 U2947 ( .A(n4685), .B(n2792), .Z(n1321) );
  HS65_LH_MX41X7 U2948 ( .D0(n4575), .S0(n1011), .D1(n4569), .S1(n4668), .D2(
        n4572), .S2(n4671), .D3(n4577), .S3(n4672), .Z(n2792) );
  HS65_LH_FA1X4 U2949 ( .A0(n551), .B0(n1287), .CI(n566), .CO(n548), .S0(n549)
         );
  HS65_LHS_XOR2X6 U2950 ( .A(n4688), .B(n2833), .Z(n1287) );
  HS65_LH_MX41X7 U2951 ( .D0(n4567), .S0(n1012), .D1(n4611), .S1(n4670), .D2(
        n4564), .S2(n4669), .D3(n4561), .S3(n4666), .Z(n2833) );
  HS65_LH_FA1X4 U2952 ( .A0(n521), .B0(n537), .CI(n1221), .CO(n518), .S0(n519)
         );
  HS65_LHS_XOR2X6 U2953 ( .A(n4694), .B(n2915), .Z(n1221) );
  HS65_LH_MX41X7 U2954 ( .D0(n4545), .S0(n1016), .D1(n4539), .S1(n4659), .D2(
        n4542), .S2(n4661), .D3(n4547), .S3(n4662), .Z(n2915) );
  HS65_LH_FA1X4 U2955 ( .A0(n517), .B0(n533), .CI(n1285), .CO(n514), .S0(n515)
         );
  HS65_LHS_XOR2X6 U2956 ( .A(n4688), .B(n2835), .Z(n1285) );
  HS65_LH_MX41X7 U2957 ( .D0(n4567), .S0(n1010), .D1(n4611), .S1(n4674), .D2(
        n4564), .S2(n4673), .D3(n4561), .S3(n4670), .Z(n2835) );
  HS65_LH_FA1X4 U2958 ( .A0(n469), .B0(n483), .CI(n1250), .CO(n466), .S0(n467)
         );
  HS65_LHS_XOR2X6 U2959 ( .A(n4691), .B(n2878), .Z(n1250) );
  HS65_LH_MX41X7 U2960 ( .D0(n4556), .S0(n1010), .D1(n4550), .S1(n4671), .D2(
        n4554), .S2(n4673), .D3(n4559), .S3(n4674), .Z(n2878) );
  HS65_LH_FA1X4 U2961 ( .A0(n430), .B0(n442), .CI(n1151), .CO(n427), .S0(n428)
         );
  HS65_LHS_XOR2X6 U2962 ( .A(n4700), .B(n3001), .Z(n1151) );
  HS65_LH_MX41X7 U2963 ( .D0(n4523), .S0(n1016), .D1(n4525), .S1(n4663), .D2(
        n4517), .S2(n4659), .D3(n4520), .S3(n4660), .Z(n3001) );
  HS65_LH_FA1X4 U2964 ( .A0(n426), .B0(n438), .CI(n1215), .CO(n423), .S0(n424)
         );
  HS65_LHS_XOR2X6 U2965 ( .A(n4694), .B(n2921), .Z(n1215) );
  HS65_LH_MX41X7 U2966 ( .D0(n4545), .S0(n1010), .D1(n4539), .S1(n4670), .D2(
        n4542), .S2(n4673), .D3(n4547), .S3(n4674), .Z(n2921) );
  HS65_LH_FA1X4 U2967 ( .A0(n394), .B0(n404), .CI(n1116), .CO(n391), .S0(n392)
         );
  HS65_LHS_XOR2X6 U2968 ( .A(n4703), .B(n3044), .Z(n1116) );
  HS65_LH_MX41X7 U2969 ( .D0(n4512), .S0(n1016), .D1(n4506), .S1(n4658), .D2(
        n4509), .S2(n4661), .D3(n4514), .S3(n4662), .Z(n3044) );
  HS65_LH_FA1X4 U2970 ( .A0(n390), .B0(n400), .CI(n1180), .CO(n387), .S0(n388)
         );
  HS65_LHS_XOR2X6 U2971 ( .A(n4698), .B(n2964), .Z(n1180) );
  HS65_LH_MX41X7 U2972 ( .D0(n2933), .S0(n1010), .D1(n4529), .S1(n4671), .D2(
        n4532), .S2(n4673), .D3(n4537), .S3(n4674), .Z(n2964) );
  HS65_LH_FA1X4 U2973 ( .A0(n359), .B0(n367), .CI(n1145), .CO(n356), .S0(n357)
         );
  HS65_LHS_XOR2X6 U2974 ( .A(n4700), .B(n3007), .Z(n1145) );
  HS65_LH_MX41X7 U2975 ( .D0(n4523), .S0(n1010), .D1(n4525), .S1(n4675), .D2(
        n4517), .S2(n4671), .D3(n4520), .S3(n4672), .Z(n3007) );
  HS65_LH_FA1X4 U2976 ( .A0(n335), .B0(n341), .CI(n1110), .CO(n332), .S0(n333)
         );
  HS65_LHS_XOR2X6 U2977 ( .A(n4704), .B(n3050), .Z(n1110) );
  HS65_LH_MX41X7 U2978 ( .D0(n4512), .S0(n1010), .D1(n4506), .S1(n4671), .D2(
        n4509), .S2(n4673), .D3(n4514), .S3(n4674), .Z(n3050) );
  HS65_LH_FA1X4 U2979 ( .A0(n571), .B0(n1256), .CI(n586), .CO(n568), .S0(n569)
         );
  HS65_LHS_XOR2X6 U2980 ( .A(n4691), .B(n2872), .Z(n1256) );
  HS65_LH_MX41X7 U2981 ( .D0(n4556), .S0(n1016), .D1(n4550), .S1(n4659), .D2(
        n4553), .S2(n4661), .D3(n4558), .S3(n4662), .Z(n2872) );
  HS65_LH_FA1X4 U2982 ( .A0(n525), .B0(n541), .CI(n1157), .CO(n522), .S0(n523)
         );
  HS65_LHS_XOR2X6 U2983 ( .A(n4700), .B(n2995), .Z(n1157) );
  HS65_LH_MX41X7 U2984 ( .D0(n4523), .S0(n1022), .D1(n4525), .S1(n4650), .D2(
        n4517), .S2(n4647), .D3(n4520), .S3(n4648), .Z(n2995) );
  HS65_LH_FA1X4 U2985 ( .A0(n601), .B0(n1386), .CI(n257), .CO(n256), .S0(
        product[33]) );
  HS65_LHS_XOR2X6 U2986 ( .A(n4682), .B(n2716), .Z(n1386) );
  HS65_LH_AOI22X6 U2987 ( .A(n4493), .B(n1006), .C(n4591), .D(n4678), .Z(n2716) );
  HS65_LH_FA1X4 U2988 ( .A0(n569), .B0(n1288), .CI(n584), .CO(n566), .S0(n567)
         );
  HS65_LHS_XOR2X6 U2989 ( .A(n4688), .B(n2832), .Z(n1288) );
  HS65_LH_MX41X7 U2990 ( .D0(n4567), .S0(n1013), .D1(n4612), .S1(n4668), .D2(
        n4565), .S2(n4667), .D3(n4561), .S3(n4664), .Z(n2832) );
  HS65_LH_FA1X4 U2991 ( .A0(n4709), .B0(n1061), .CI(n1093), .CO(n526), .S0(
        n527) );
  HS65_LH_MX41X7 U2992 ( .D0(n1031), .S0(n4490), .D1(n4632), .S1(n4607), .D2(
        n4630), .S2(n4602), .D3(n4628), .S3(n4609), .Z(n1061) );
  HS65_LHS_XOR2X6 U2993 ( .A(n4706), .B(n3075), .Z(n1093) );
  HS65_LH_MX41X7 U2994 ( .D0(n4501), .S0(n1028), .D1(n4495), .S1(n4635), .D2(
        n4498), .S2(n4637), .D3(n4503), .S3(n4638), .Z(n3075) );
  HS65_LH_FA1X4 U2995 ( .A0(n4713), .B0(n446), .CI(n1087), .CO(n431), .S0(n432) );
  HS65_LHS_XOR2X6 U2996 ( .A(n4706), .B(n3081), .Z(n1087) );
  HS65_LH_MX41X7 U2997 ( .D0(n4501), .S0(n1022), .D1(n4495), .S1(n4647), .D2(
        n4498), .S2(n4649), .D3(n4503), .S3(n4650), .Z(n3081) );
  HS65_LH_FA1X4 U2998 ( .A0(n4714), .B0(n371), .CI(n1081), .CO(n360), .S0(n361) );
  HS65_LHS_XOR2X6 U2999 ( .A(n4706), .B(n3087), .Z(n1081) );
  HS65_LH_MX41X7 U3000 ( .D0(n4501), .S0(n1016), .D1(n4495), .S1(n4659), .D2(
        n4498), .S2(n4661), .D3(n4503), .S3(n4662), .Z(n3087) );
  HS65_LH_FA1X4 U3001 ( .A0(n4715), .B0(n320), .CI(n1075), .CO(n313), .S0(n314) );
  HS65_LHS_XOR2X6 U3002 ( .A(n4707), .B(n3093), .Z(n1075) );
  HS65_LH_MX41X7 U3003 ( .D0(n4501), .S0(n1010), .D1(n4495), .S1(n4671), .D2(
        n4498), .S2(n4673), .D3(n4504), .S3(n4674), .Z(n3093) );
  HS65_LH_FA1X4 U3004 ( .A0(n1065), .B0(n4680), .CI(n1097), .CO(n598), .S0(
        n599) );
  HS65_LH_MX41X7 U3005 ( .D0(n1035), .S0(n4492), .D1(n4624), .S1(n4608), .D2(
        n4622), .S2(n4604), .D3(n4620), .S3(n4609), .Z(n1065) );
  HS65_LHS_XOR2X6 U3006 ( .A(n4707), .B(n3071), .Z(n1097) );
  HS65_LH_MX41X7 U3007 ( .D0(n3062), .S0(n1032), .D1(n4496), .S1(n4627), .D2(
        n4499), .S2(n4629), .D3(n4504), .S3(n4630), .Z(n3071) );
  HS65_LH_FA1X4 U3008 ( .A0(n1064), .B0(n4680), .CI(n598), .CO(n580), .S0(n581) );
  HS65_LH_MX41X7 U3009 ( .D0(n1034), .S0(n4490), .D1(n4626), .S1(n4608), .D2(
        n4624), .S2(n4602), .D3(n4622), .S3(n4609), .Z(n1064) );
  HS65_LH_FA1X4 U3010 ( .A0(n1060), .B0(n4709), .CI(n526), .CO(n508), .S0(n509) );
  HS65_LH_MX41X7 U3011 ( .D0(n1030), .S0(n4491), .D1(n4634), .S1(n4607), .D2(
        n4632), .S2(n4603), .D3(n4630), .S3(n4609), .Z(n1060) );
  HS65_LH_FA1X4 U3012 ( .A0(n1055), .B0(n4713), .CI(n431), .CO(n417), .S0(n418) );
  HS65_LH_MX41X7 U3013 ( .D0(n1024), .S0(n4491), .D1(n4644), .S1(n4602), .D2(
        n4642), .S2(n4610), .D3(n4646), .S3(n4606), .Z(n1055) );
  HS65_LH_FA1X4 U3014 ( .A0(n1050), .B0(n4714), .CI(n360), .CO(n350), .S0(n351) );
  HS65_LH_MX41X7 U3015 ( .D0(n1018), .S0(n4490), .D1(n4654), .S1(n4609), .D2(
        n4656), .S2(n4602), .D3(n4658), .S3(n4606), .Z(n1050) );
  HS65_LH_FA1X4 U3016 ( .A0(n1045), .B0(n4715), .CI(n313), .CO(n307), .S0(n308) );
  HS65_LH_MX41X7 U3017 ( .D0(n1012), .S0(n4491), .D1(n4666), .S1(n4610), .D2(
        n4668), .S2(n4603), .D3(n4670), .S3(n4607), .Z(n1045) );
  HS65_LH_MX41X7 U3018 ( .D0(n4567), .S0(n1009), .D1(n4612), .S1(n4677), .D2(
        n4564), .S2(n4675), .D3(n4561), .S3(n4672), .Z(n2836) );
  HS65_LH_MX41X7 U3019 ( .D0(n4512), .S0(n1028), .D1(n4507), .S1(n4634), .D2(
        n4510), .S2(n4637), .D3(n4515), .S3(n4638), .Z(n3032) );
  HS65_LH_MX41X7 U3020 ( .D0(n4512), .S0(n1027), .D1(n4507), .S1(n4636), .D2(
        n4510), .S2(n4639), .D3(n4515), .S3(n4640), .Z(n3033) );
  HS65_LH_MX41X7 U3021 ( .D0(n4534), .S0(n1022), .D1(n4528), .S1(n4647), .D2(
        n4531), .S2(n4649), .D3(n4536), .S3(n4650), .Z(n2952) );
  HS65_LH_MX41X7 U3022 ( .D0(n4534), .S0(n1021), .D1(n4528), .S1(n4649), .D2(
        n4532), .S2(n4651), .D3(n4536), .S3(n4652), .Z(n2953) );
  HS65_LH_MX41X7 U3023 ( .D0(n3062), .S0(n1027), .D1(n4496), .S1(n4637), .D2(
        n4499), .S2(n4639), .D3(n4504), .S3(n4640), .Z(n3076) );
  HS65_LH_MX41X7 U3024 ( .D0(n2762), .S0(n1010), .D1(n4570), .S1(n4670), .D2(
        n4573), .S2(n4673), .D3(n4578), .S3(n4674), .Z(n2793) );
  HS65_LH_MX41X7 U3025 ( .D0(n4545), .S0(n1015), .D1(n4539), .S1(n4661), .D2(
        n4542), .S2(n4663), .D3(n4547), .S3(n4664), .Z(n2916) );
  HS65_LH_MX41X7 U3026 ( .D0(n4512), .S0(n1021), .D1(n4506), .S1(n4648), .D2(
        n4509), .S2(n4651), .D3(n4515), .S3(n4652), .Z(n3039) );
  HS65_LH_MX41X7 U3027 ( .D0(n4534), .S0(n1015), .D1(n4528), .S1(n4660), .D2(
        n4531), .S2(n4663), .D3(n4536), .S3(n4664), .Z(n2959) );
  HS65_LH_MX41X7 U3028 ( .D0(n4501), .S0(n1021), .D1(n4495), .S1(n4648), .D2(
        n4499), .S2(n4651), .D3(n4504), .S3(n4652), .Z(n3082) );
  HS65_LH_MX41X7 U3029 ( .D0(n4545), .S0(n1009), .D1(n4539), .S1(n4672), .D2(
        n4542), .S2(n4675), .D3(n4547), .S3(n4676), .Z(n2922) );
  HS65_LH_MX41X7 U3030 ( .D0(n4512), .S0(n1015), .D1(n4506), .S1(n4661), .D2(
        n4509), .S2(n4663), .D3(n4514), .S3(n4664), .Z(n3045) );
  HS65_LH_MX41X7 U3031 ( .D0(n2933), .S0(n1009), .D1(n4529), .S1(n4672), .D2(
        n4532), .S2(n4675), .D3(n4537), .S3(n4677), .Z(n2965) );
  HS65_LH_MX41X7 U3032 ( .D0(n4501), .S0(n1015), .D1(n4495), .S1(n4660), .D2(
        n4498), .S2(n4663), .D3(n4503), .S3(n4664), .Z(n3088) );
  HS65_LH_MX41X7 U3033 ( .D0(n4512), .S0(n1009), .D1(n4506), .S1(n4673), .D2(
        n4509), .S2(n4675), .D3(n4514), .S3(n4676), .Z(n3051) );
  HS65_LH_MX41X7 U3034 ( .D0(n4501), .S0(n1009), .D1(n4496), .S1(n4673), .D2(
        n4499), .S2(n4675), .D3(n4504), .S3(n4676), .Z(n3094) );
  HS65_LH_MX41X7 U3035 ( .D0(n2762), .S0(n1009), .D1(n4570), .S1(n4673), .D2(
        n4573), .S2(n4675), .D3(n4579), .S3(n4677), .Z(n2794) );
  HS65_LH_MX41X7 U3036 ( .D0(n2847), .S0(n1009), .D1(n4551), .S1(n4673), .D2(
        n4554), .S2(n4675), .D3(n4560), .S3(n4677), .Z(n2879) );
  HS65_LH_MX41X7 U3037 ( .D0(n2976), .S0(n1021), .D1(n4526), .S1(n4652), .D2(
        n4518), .S2(n4649), .D3(n4521), .S3(n4650), .Z(n2996) );
  HS65_LH_MX41X7 U3038 ( .D0(n4523), .S0(n1015), .D1(n4525), .S1(n4664), .D2(
        n4517), .S2(n4661), .D3(n4520), .S3(n4662), .Z(n3002) );
  HS65_LH_MX41X7 U3039 ( .D0(n2976), .S0(n1009), .D1(n4526), .S1(n4677), .D2(
        n4518), .S2(n4673), .D3(n4521), .S3(n4674), .Z(n3008) );
  HS65_LH_FA1X4 U3040 ( .A0(n4622), .B0(n4624), .CI(n1003), .CO(n1002), .S0(
        n1035) );
  HS65_LH_FA1X4 U3041 ( .A0(n4624), .B0(n4626), .CI(n1002), .CO(n1001), .S0(
        n1034) );
  HS65_LH_FA1X4 U3042 ( .A0(n4626), .B0(n4628), .CI(n1001), .CO(n1000), .S0(
        n1033) );
  HS65_LH_FA1X4 U3043 ( .A0(n4628), .B0(n4630), .CI(n1000), .CO(n999), .S0(
        n1032) );
  HS65_LH_FA1X4 U3044 ( .A0(n4630), .B0(n4632), .CI(n999), .CO(n998), .S0(
        n1031) );
  HS65_LH_FA1X4 U3045 ( .A0(n4632), .B0(n4634), .CI(n998), .CO(n997), .S0(
        n1030) );
  HS65_LH_FA1X4 U3046 ( .A0(n4634), .B0(n4636), .CI(n997), .CO(n996), .S0(
        n1029) );
  HS65_LH_FA1X4 U3047 ( .A0(n4636), .B0(n4638), .CI(n996), .CO(n995), .S0(
        n1028) );
  HS65_LH_FA1X4 U3048 ( .A0(n4638), .B0(n4640), .CI(n995), .CO(n994), .S0(
        n1027) );
  HS65_LH_FA1X4 U3049 ( .A0(n4640), .B0(n4642), .CI(n994), .CO(n993), .S0(
        n1026) );
  HS65_LH_FA1X4 U3050 ( .A0(n4642), .B0(n4644), .CI(n993), .CO(n992), .S0(
        n1025) );
  HS65_LH_FA1X4 U3051 ( .A0(n4644), .B0(n4646), .CI(n992), .CO(n991), .S0(
        n1024) );
  HS65_LH_FA1X4 U3052 ( .A0(n4646), .B0(n4648), .CI(n991), .CO(n990), .S0(
        n1023) );
  HS65_LH_FA1X4 U3053 ( .A0(n4648), .B0(n4650), .CI(n990), .CO(n989), .S0(
        n1022) );
  HS65_LH_FA1X4 U3054 ( .A0(n4650), .B0(n4652), .CI(n989), .CO(n988), .S0(
        n1021) );
  HS65_LH_FA1X4 U3055 ( .A0(n4652), .B0(n4654), .CI(n988), .CO(n987), .S0(
        n1020) );
  HS65_LH_FA1X4 U3056 ( .A0(n4654), .B0(n4656), .CI(n987), .CO(n986), .S0(
        n1019) );
  HS65_LH_FA1X4 U3057 ( .A0(n4656), .B0(n4658), .CI(n986), .CO(n985), .S0(
        n1018) );
  HS65_LH_FA1X4 U3058 ( .A0(n4658), .B0(n4660), .CI(n985), .CO(n984), .S0(
        n1017) );
  HS65_LH_FA1X4 U3059 ( .A0(n4662), .B0(n4664), .CI(n983), .CO(n982), .S0(
        n1015) );
  HS65_LH_FA1X4 U3060 ( .A0(n4664), .B0(n4666), .CI(n982), .CO(n981), .S0(
        n1014) );
  HS65_LH_FA1X4 U3061 ( .A0(n4666), .B0(n4668), .CI(n981), .CO(n980), .S0(
        n1013) );
  HS65_LH_FA1X4 U3062 ( .A0(n4668), .B0(n4670), .CI(n980), .CO(n979), .S0(
        n1012) );
  HS65_LH_FA1X4 U3063 ( .A0(n4670), .B0(n4672), .CI(n979), .CO(n978), .S0(
        n1011) );
  HS65_LH_FA1X4 U3064 ( .A0(n4672), .B0(n4674), .CI(n978), .CO(n977), .S0(
        n1010) );
  HS65_LH_FA1X4 U3065 ( .A0(n297), .B0(n4708), .CI(n1041), .CO(n293), .S0(n294) );
  HS65_LH_MX41X7 U3066 ( .D0(n1008), .S0(n4492), .D1(n4674), .S1(n4609), .D2(
        n4676), .S2(n4604), .D3(n4606), .S3(n4679), .Z(n1041) );
  HS65_LH_FA1X4 U3067 ( .A0(n557), .B0(n1191), .CI(n1223), .CO(n554), .S0(n555) );
  HS65_LHS_XOR2X6 U3068 ( .A(n4694), .B(n2913), .Z(n1223) );
  HS65_LHS_XOR2X6 U3069 ( .A(n4697), .B(n2953), .Z(n1191) );
  HS65_LH_MX41X7 U3070 ( .D0(n4545), .S0(n1018), .D1(n4539), .S1(n4655), .D2(
        n4542), .S2(n4657), .D3(n4547), .S3(n4658), .Z(n2913) );
  HS65_LH_FA1X4 U3071 ( .A0(n509), .B0(n1092), .CI(n1124), .CO(n506), .S0(n507) );
  HS65_LHS_XOR2X6 U3072 ( .A(n4704), .B(n3036), .Z(n1124) );
  HS65_LHS_XOR2X6 U3073 ( .A(n4707), .B(n3076), .Z(n1092) );
  HS65_LH_MX41X7 U3074 ( .D0(n4512), .S0(n1024), .D1(n4506), .S1(n4642), .D2(
        n4509), .S2(n4645), .D3(n4515), .S3(n4646), .Z(n3036) );
  HS65_LH_FA1X4 U3075 ( .A0(n553), .B0(n1255), .CI(n568), .CO(n550), .S0(n551)
         );
  HS65_LHS_XOR2X6 U3076 ( .A(n4691), .B(n2873), .Z(n1255) );
  HS65_LH_MX41X7 U3077 ( .D0(n4556), .S0(n1015), .D1(n4550), .S1(n4661), .D2(
        n4553), .S2(n4663), .D3(n4558), .S3(n4664), .Z(n2873) );
  HS65_LH_FA1X4 U3078 ( .A0(n505), .B0(n1156), .CI(n1188), .CO(n502), .S0(n503) );
  HS65_LHS_XOR2X6 U3079 ( .A(n4698), .B(n2956), .Z(n1188) );
  HS65_LHS_XOR2X6 U3080 ( .A(n4701), .B(n2996), .Z(n1156) );
  HS65_LH_MX41X7 U3081 ( .D0(n4534), .S0(n1018), .D1(n4528), .S1(n4655), .D2(
        n4531), .S2(n4657), .D3(n4536), .S3(n4658), .Z(n2956) );
  HS65_LH_FA1X4 U3082 ( .A0(n501), .B0(n1220), .CI(n1252), .CO(n498), .S0(n499) );
  HS65_LHS_XOR2X6 U3083 ( .A(n4691), .B(n2876), .Z(n1252) );
  HS65_LHS_XOR2X6 U3084 ( .A(n4695), .B(n2916), .Z(n1220) );
  HS65_LH_MX41X7 U3085 ( .D0(n4556), .S0(n1012), .D1(n4550), .S1(n4667), .D2(
        n4553), .S2(n4669), .D3(n4558), .S3(n4670), .Z(n2876) );
  HS65_LH_FA1X4 U3086 ( .A0(n459), .B0(n1121), .CI(n1153), .CO(n456), .S0(n457) );
  HS65_LHS_XOR2X6 U3087 ( .A(n4700), .B(n2999), .Z(n1153) );
  HS65_LHS_XOR2X6 U3088 ( .A(n4704), .B(n3039), .Z(n1121) );
  HS65_LH_MX41X7 U3089 ( .D0(n4523), .S0(n1018), .D1(n4525), .S1(n4658), .D2(
        n4517), .S2(n4655), .D3(n4520), .S3(n4656), .Z(n2999) );
  HS65_LH_FA1X4 U3090 ( .A0(n455), .B0(n1185), .CI(n1217), .CO(n452), .S0(n453) );
  HS65_LHS_XOR2X6 U3091 ( .A(n4694), .B(n2919), .Z(n1217) );
  HS65_LHS_XOR2X6 U3092 ( .A(n4697), .B(n2959), .Z(n1185) );
  HS65_LH_MX41X7 U3093 ( .D0(n4545), .S0(n1012), .D1(n4539), .S1(n4666), .D2(
        n4543), .S2(n4669), .D3(n4548), .S3(n4670), .Z(n2919) );
  HS65_LH_FA1X4 U3094 ( .A0(n418), .B0(n1086), .CI(n1118), .CO(n415), .S0(n416) );
  HS65_LHS_XOR2X6 U3095 ( .A(n4703), .B(n3042), .Z(n1118) );
  HS65_LHS_XOR2X6 U3096 ( .A(n4707), .B(n3082), .Z(n1086) );
  HS65_LH_MX41X7 U3097 ( .D0(n4512), .S0(n1018), .D1(n4506), .S1(n4654), .D2(
        n4509), .S2(n4657), .D3(n4514), .S3(n4658), .Z(n3042) );
  HS65_LH_FA1X4 U3098 ( .A0(n414), .B0(n1150), .CI(n1182), .CO(n411), .S0(n412) );
  HS65_LHS_XOR2X6 U3099 ( .A(n4697), .B(n2962), .Z(n1182) );
  HS65_LHS_XOR2X6 U3100 ( .A(n4700), .B(n3002), .Z(n1150) );
  HS65_LH_MX41X7 U3101 ( .D0(n4534), .S0(n1012), .D1(n4528), .S1(n4666), .D2(
        n4531), .S2(n4669), .D3(n4536), .S3(n4670), .Z(n2962) );
  HS65_LH_FA1X4 U3102 ( .A0(n380), .B0(n1115), .CI(n1147), .CO(n377), .S0(n378) );
  HS65_LHS_XOR2X6 U3103 ( .A(n4700), .B(n3005), .Z(n1147) );
  HS65_LHS_XOR2X6 U3104 ( .A(n4703), .B(n3045), .Z(n1115) );
  HS65_LH_MX41X7 U3105 ( .D0(n4523), .S0(n1012), .D1(n4525), .S1(n4671), .D2(
        n4518), .S2(n4667), .D3(n4521), .S3(n4668), .Z(n3005) );
  HS65_LH_FA1X4 U3106 ( .A0(n351), .B0(n1080), .CI(n1112), .CO(n348), .S0(n349) );
  HS65_LHS_XOR2X6 U3107 ( .A(n4703), .B(n3048), .Z(n1112) );
  HS65_LHS_XOR2X6 U3108 ( .A(n4707), .B(n3088), .Z(n1080) );
  HS65_LH_MX41X7 U3109 ( .D0(n4512), .S0(n1012), .D1(n4506), .S1(n4666), .D2(
        n4510), .S2(n4669), .D3(n4514), .S3(n4670), .Z(n3048) );
  HS65_LH_FA1X4 U3110 ( .A0(n1063), .B0(n4680), .CI(n580), .CO(n562), .S0(n563) );
  HS65_LH_MX41X7 U3111 ( .D0(n1033), .S0(n4492), .D1(n4628), .S1(n4608), .D2(
        n4626), .S2(n4603), .D3(n4624), .S3(n4609), .Z(n1063) );
  HS65_LH_FA1X4 U3112 ( .A0(n1057), .B0(n4710), .CI(n1089), .CO(n460), .S0(
        n461) );
  HS65_LH_MX41X7 U3113 ( .D0(n1027), .S0(n4491), .D1(n4606), .S1(n4640), .D2(
        n4638), .S2(n4603), .D3(n4636), .S3(n4609), .Z(n1057) );
  HS65_LHS_XOR2X6 U3114 ( .A(n4706), .B(n3079), .Z(n1089) );
  HS65_LH_MX41X7 U3115 ( .D0(n4501), .S0(n1024), .D1(n4495), .S1(n4642), .D2(
        n4498), .S2(n4645), .D3(n4503), .S3(n4646), .Z(n3079) );
  HS65_LH_FA1X4 U3116 ( .A0(n1052), .B0(n4711), .CI(n1083), .CO(n381), .S0(
        n382) );
  HS65_LH_MX41X7 U3117 ( .D0(n1021), .S0(n4490), .D1(n4648), .S1(n4610), .D2(
        n4650), .S2(n4602), .D3(n4652), .S3(n4606), .Z(n1052) );
  HS65_LHS_XOR2X6 U3118 ( .A(n4706), .B(n3085), .Z(n1083) );
  HS65_LH_MX41X7 U3119 ( .D0(n4501), .S0(n1018), .D1(n4495), .S1(n4654), .D2(
        n4498), .S2(n4657), .D3(n4503), .S3(n4658), .Z(n3085) );
  HS65_LH_FA1X4 U3120 ( .A0(n1047), .B0(n4712), .CI(n1077), .CO(n326), .S0(
        n327) );
  HS65_LH_MX41X7 U3121 ( .D0(n1015), .S0(n4490), .D1(n4660), .S1(n4610), .D2(
        n4662), .S2(n4602), .D3(n4664), .S3(n4606), .Z(n1047) );
  HS65_LHS_XOR2X6 U3122 ( .A(n4706), .B(n3091), .Z(n1077) );
  HS65_LH_MX41X7 U3123 ( .D0(n4501), .S0(n1012), .D1(n4495), .S1(n4666), .D2(
        n4498), .S2(n4669), .D3(n4503), .S3(n4670), .Z(n3091) );
  HS65_LH_FA1X4 U3124 ( .A0(n1042), .B0(n4716), .CI(n1071), .CO(n295), .S0(
        n296) );
  HS65_LH_MX41X7 U3125 ( .D0(n1009), .S0(n4490), .D1(n4672), .S1(n4609), .D2(
        n4674), .S2(n4602), .D3(n4676), .S3(n4606), .Z(n1042) );
  HS65_LHS_XOR2X6 U3126 ( .A(n4708), .B(n3102), .Z(n1071) );
  HS65_LH_AOI22X6 U3127 ( .A(n4501), .B(n1006), .C(n4495), .D(n4678), .Z(n3102) );
  HS65_LH_IVX9 U3128 ( .A(n31), .Z(n4687) );
  HS65_LH_IVX9 U3129 ( .A(n55), .Z(n4693) );
  HS65_LH_IVX9 U3130 ( .A(n67), .Z(n4696) );
  HS65_LH_IVX9 U3131 ( .A(n115), .Z(n4708) );
  HS65_LH_IVX9 U3132 ( .A(n79), .Z(n4699) );
  HS65_LH_IVX9 U3133 ( .A(n43), .Z(n4690) );
  HS65_LH_IVX9 U3134 ( .A(n103), .Z(n4705) );
  HS65_LH_IVX9 U3135 ( .A(n91), .Z(n4702) );
  HS65_LH_IVX9 U3136 ( .A(n4587), .Z(n4586) );
  HS65_LH_IVX9 U3137 ( .A(n4576), .Z(n4575) );
  HS65_LH_IVX9 U3138 ( .A(n4568), .Z(n4567) );
  HS65_LH_IVX9 U3139 ( .A(n4557), .Z(n4556) );
  HS65_LH_IVX9 U3140 ( .A(n4546), .Z(n4545) );
  HS65_LH_IVX9 U3141 ( .A(n4535), .Z(n4534) );
  HS65_LH_IVX9 U3142 ( .A(n4524), .Z(n4523) );
  HS65_LH_IVX9 U3143 ( .A(n4513), .Z(n4512) );
  HS65_LH_IVX9 U3144 ( .A(n4502), .Z(n4501) );
  HS65_LH_BFX9 U3145 ( .A(b[30]), .Z(n4676) );
  HS65_LH_AND2X4 U3146 ( .A(n4594), .B(n4679), .Z(n2715) );
  HS65_LH_BFX9 U3147 ( .A(n2723), .Z(n4580) );
  HS65_LH_BFX9 U3148 ( .A(n2766), .Z(n4569) );
  HS65_LH_BFX9 U3149 ( .A(n2851), .Z(n4550) );
  HS65_LH_BFX9 U3150 ( .A(n2894), .Z(n4539) );
  HS65_LH_BFX9 U3151 ( .A(n2937), .Z(n4528) );
  HS65_LH_BFX9 U3152 ( .A(n3023), .Z(n4506) );
  HS65_LH_BFX9 U3153 ( .A(n3066), .Z(n4495) );
  HS65_LH_BFX9 U3154 ( .A(n2808), .Z(n4561) );
  HS65_LH_BFX9 U3155 ( .A(n2980), .Z(n4517) );
  HS65_LH_BFX9 U3156 ( .A(b[31]), .Z(n4678) );
  HS65_LH_BFX9 U3157 ( .A(n2980), .Z(n4518) );
  HS65_LH_BFX9 U3158 ( .A(n2723), .Z(n4581) );
  HS65_LH_BFX9 U3159 ( .A(n3066), .Z(n4496) );
  HS65_LH_BFX9 U3160 ( .A(n2894), .Z(n4540) );
  HS65_LH_BFX9 U3161 ( .A(n2766), .Z(n4570) );
  HS65_LH_BFX9 U3162 ( .A(n3023), .Z(n4507) );
  HS65_LH_BFX9 U3163 ( .A(n2851), .Z(n4551) );
  HS65_LH_BFX9 U3164 ( .A(n2937), .Z(n4529) );
  HS65_LH_BFX9 U3165 ( .A(n2808), .Z(n4562) );
  HS65_LH_BFX9 U3166 ( .A(b[3]), .Z(n4622) );
  HS65_LH_BFX9 U3167 ( .A(b[23]), .Z(n4662) );
  HS65_LH_BFX9 U3168 ( .A(b[2]), .Z(n4620) );
  HS65_LH_BFX9 U3169 ( .A(b[22]), .Z(n4660) );
  HS65_LH_BFX9 U3170 ( .A(b[29]), .Z(n4674) );
  HS65_LH_BFX9 U3171 ( .A(b[0]), .Z(n4614) );
  HS65_LH_BFX9 U3172 ( .A(b[1]), .Z(n4618) );
  HS65_LH_BFX9 U3173 ( .A(n4718), .Z(n4493) );
  HS65_LH_BFX9 U3174 ( .A(n2417), .Z(n4611) );
  HS65_LH_BFX9 U3175 ( .A(n2417), .Z(n4612) );
  HS65_LH_BFX9 U3176 ( .A(n2975), .Z(n4526) );
  HS65_LH_BFX9 U3177 ( .A(n2975), .Z(n4525) );
  HS65_LH_BFX9 U3178 ( .A(n2932), .Z(n4537) );
  HS65_LH_BFX9 U3179 ( .A(n2718), .Z(n4589) );
  HS65_LH_BFX9 U3180 ( .A(n2846), .Z(n4559) );
  HS65_LH_BFX9 U3181 ( .A(n3061), .Z(n4504) );
  HS65_LH_BFX9 U3182 ( .A(n2761), .Z(n4577) );
  HS65_LH_BFX9 U3183 ( .A(n2761), .Z(n4578) );
  HS65_LH_BFX9 U3184 ( .A(n2718), .Z(n4588) );
  HS65_LH_BFX9 U3185 ( .A(n3018), .Z(n4515) );
  HS65_LH_BFX9 U3186 ( .A(n2889), .Z(n4547) );
  HS65_LH_BFX9 U3187 ( .A(n2846), .Z(n4558) );
  HS65_LH_BFX9 U3188 ( .A(n2889), .Z(n4548) );
  HS65_LH_BFX9 U3189 ( .A(n2932), .Z(n4536) );
  HS65_LH_BFX9 U3190 ( .A(n3018), .Z(n4514) );
  HS65_LH_BFX9 U3191 ( .A(n3061), .Z(n4503) );
  HS65_LH_BFX9 U3192 ( .A(n4717), .Z(n4491) );
  HS65_LH_BFX9 U3193 ( .A(b[31]), .Z(n4679) );
  HS65_LH_BFX9 U3194 ( .A(n4717), .Z(n4490) );
  HS65_LH_BFX9 U3195 ( .A(b[3]), .Z(n4623) );
  HS65_LH_BFX9 U3196 ( .A(b[2]), .Z(n4621) );
  HS65_LH_BFX9 U3197 ( .A(b[23]), .Z(n4663) );
  HS65_LH_BFX9 U3198 ( .A(b[30]), .Z(n4677) );
  HS65_LH_BFX9 U3199 ( .A(b[22]), .Z(n4661) );
  HS65_LH_BFX9 U3200 ( .A(b[29]), .Z(n4675) );
  HS65_LH_BFX9 U3201 ( .A(b[1]), .Z(n4619) );
  HS65_LH_BFX9 U3202 ( .A(n4718), .Z(n4494) );
  HS65_LH_BFX9 U3203 ( .A(n4582), .Z(n4584) );
  HS65_LH_BFX9 U3204 ( .A(n4571), .Z(n4573) );
  HS65_LH_BFX9 U3205 ( .A(n4563), .Z(n4565) );
  HS65_LH_BFX9 U3206 ( .A(n4552), .Z(n4554) );
  HS65_LH_BFX9 U3207 ( .A(n4497), .Z(n4499) );
  HS65_LH_BFX9 U3208 ( .A(n4571), .Z(n4572) );
  HS65_LH_BFX9 U3209 ( .A(n4563), .Z(n4564) );
  HS65_LH_BFX9 U3210 ( .A(n4582), .Z(n4583) );
  HS65_LH_BFX9 U3211 ( .A(n4541), .Z(n4542) );
  HS65_LH_BFX9 U3212 ( .A(n4552), .Z(n4553) );
  HS65_LH_BFX9 U3213 ( .A(n4541), .Z(n4543) );
  HS65_LH_BFX9 U3214 ( .A(n4508), .Z(n4509) );
  HS65_LH_BFX9 U3215 ( .A(n4530), .Z(n4532) );
  HS65_LH_BFX9 U3216 ( .A(n4530), .Z(n4531) );
  HS65_LH_BFX9 U3217 ( .A(n4508), .Z(n4510) );
  HS65_LH_BFX9 U3218 ( .A(n4497), .Z(n4498) );
  HS65_LH_BFX9 U3219 ( .A(n4601), .Z(n4602) );
  HS65_LH_BFX9 U3220 ( .A(n4519), .Z(n4520) );
  HS65_LH_BFX9 U3221 ( .A(n4519), .Z(n4521) );
  HS65_LH_BFX9 U3222 ( .A(n4601), .Z(n4603) );
  HS65_LH_BFX9 U3223 ( .A(n2975), .Z(n4527) );
  HS65_LH_BFX9 U3224 ( .A(n2718), .Z(n4590) );
  HS65_LH_BFX9 U3225 ( .A(n2761), .Z(n4579) );
  HS65_LH_BFX9 U3226 ( .A(n2846), .Z(n4560) );
  HS65_LH_BFX9 U3227 ( .A(n2889), .Z(n4549) );
  HS65_LH_BFX9 U3228 ( .A(n2932), .Z(n4538) );
  HS65_LH_BFX9 U3229 ( .A(n3018), .Z(n4516) );
  HS65_LH_BFX9 U3230 ( .A(n3061), .Z(n4505) );
  HS65_LH_BFX9 U3231 ( .A(n2417), .Z(n4613) );
  HS65_LH_BFX9 U3232 ( .A(n4717), .Z(n4492) );
  HS65_LH_BFX9 U3233 ( .A(n4582), .Z(n4585) );
  HS65_LH_BFX9 U3234 ( .A(n4571), .Z(n4574) );
  HS65_LH_BFX9 U3235 ( .A(n4552), .Z(n4555) );
  HS65_LH_BFX9 U3236 ( .A(n4541), .Z(n4544) );
  HS65_LH_BFX9 U3237 ( .A(n4530), .Z(n4533) );
  HS65_LH_BFX9 U3238 ( .A(n4508), .Z(n4511) );
  HS65_LH_BFX9 U3239 ( .A(n4497), .Z(n4500) );
  HS65_LH_BFX9 U3240 ( .A(n4563), .Z(n4566) );
  HS65_LH_BFX9 U3241 ( .A(n4519), .Z(n4522) );
  HS65_LH_BFX9 U3242 ( .A(n4601), .Z(n4604) );
  HS65_LH_IVX9 U3243 ( .A(n2673), .Z(n4717) );
  HS65_LH_IVX9 U3244 ( .A(n2713), .Z(n4718) );
  HS65_LH_IVX9 U3245 ( .A(n2719), .Z(n4587) );
  HS65_LH_NOR2AX3 U3246 ( .A(n2753), .B(n2754), .Z(n2719) );
  HS65_LH_IVX9 U3247 ( .A(n2762), .Z(n4576) );
  HS65_LH_NOR2AX3 U3248 ( .A(n2796), .B(n2797), .Z(n2762) );
  HS65_LH_IVX9 U3249 ( .A(n2804), .Z(n4568) );
  HS65_LH_NOR2AX3 U3250 ( .A(n2838), .B(n2839), .Z(n2804) );
  HS65_LH_IVX9 U3251 ( .A(n2847), .Z(n4557) );
  HS65_LH_NOR2AX3 U3252 ( .A(n2881), .B(n2882), .Z(n2847) );
  HS65_LH_IVX9 U3253 ( .A(n2890), .Z(n4546) );
  HS65_LH_NOR2AX3 U3254 ( .A(n2924), .B(n2925), .Z(n2890) );
  HS65_LH_IVX9 U3255 ( .A(n2933), .Z(n4535) );
  HS65_LH_NOR2AX3 U3256 ( .A(n2967), .B(n2968), .Z(n2933) );
  HS65_LH_IVX9 U3257 ( .A(n2976), .Z(n4524) );
  HS65_LH_NOR2AX3 U3258 ( .A(n3010), .B(n3011), .Z(n2976) );
  HS65_LH_IVX9 U3259 ( .A(n3019), .Z(n4513) );
  HS65_LH_NOR2AX3 U3260 ( .A(n3053), .B(n3054), .Z(n3019) );
  HS65_LH_IVX9 U3261 ( .A(n3062), .Z(n4502) );
  HS65_LH_NOR2AX3 U3262 ( .A(n3096), .B(n3097), .Z(n3062) );
  HS65_LH_IVX9 U3263 ( .A(n4682), .Z(n4680) );
  HS65_LH_IVX9 U3264 ( .A(n7), .Z(n4682) );
  HS65_LH_IVX9 U3265 ( .A(n4682), .Z(n4681) );
  HS65_LH_FA1X4 U3266 ( .A0(n1387), .B0(n619), .CI(n258), .CO(n257), .S0(
        product[32]) );
  HS65_LHS_XOR2X6 U3267 ( .A(n4681), .B(n2712), .Z(n1387) );
  HS65_LH_OAI21X3 U3268 ( .A(n4719), .B(n2713), .C(n2714), .Z(n2712) );
  HS65_LH_OAI22X6 U3269 ( .A(n4676), .B(n2715), .C(n4591), .D(n2715), .Z(n2714) );
  HS65_LH_OA12X9 U3270 ( .A(n2673), .B(n4719), .C(n2674), .Z(n292) );
  HS65_LH_OAI22X6 U3271 ( .A(n4676), .B(n2675), .C(n4609), .D(n2675), .Z(n2674) );
  HS65_LH_AND2X4 U3272 ( .A(n4678), .B(n4602), .Z(n2675) );
  HS65_LH_BFX9 U3273 ( .A(n2670), .Z(n4609) );
  HS65_LH_BFX9 U3274 ( .A(n2681), .Z(n4591) );
  HS65_LH_BFX9 U3275 ( .A(n2672), .Z(n4601) );
  HS65_LH_NOR2AX3 U3276 ( .A(n3104), .B(n3103), .Z(n2672) );
  HS65_LH_BFX9 U3277 ( .A(n2721), .Z(n4582) );
  HS65_LH_NOR2X6 U3278 ( .A(n2753), .B(n2758), .Z(n2721) );
  HS65_LH_BFX9 U3279 ( .A(n2764), .Z(n4571) );
  HS65_LH_NOR2X6 U3280 ( .A(n2796), .B(n2801), .Z(n2764) );
  HS65_LH_BFX9 U3281 ( .A(n2806), .Z(n4563) );
  HS65_LH_NOR2X6 U3282 ( .A(n2838), .B(n2843), .Z(n2806) );
  HS65_LH_BFX9 U3283 ( .A(n2849), .Z(n4552) );
  HS65_LH_NOR2X6 U3284 ( .A(n2881), .B(n2886), .Z(n2849) );
  HS65_LH_BFX9 U3285 ( .A(n2892), .Z(n4541) );
  HS65_LH_NOR2X6 U3286 ( .A(n2924), .B(n2929), .Z(n2892) );
  HS65_LH_BFX9 U3287 ( .A(n2935), .Z(n4530) );
  HS65_LH_NOR2X6 U3288 ( .A(n2967), .B(n2972), .Z(n2935) );
  HS65_LH_BFX9 U3289 ( .A(n2978), .Z(n4519) );
  HS65_LH_NOR2X6 U3290 ( .A(n3010), .B(n3015), .Z(n2978) );
  HS65_LH_BFX9 U3291 ( .A(n3021), .Z(n4508) );
  HS65_LH_NOR2X6 U3292 ( .A(n3053), .B(n3058), .Z(n3021) );
  HS65_LH_BFX9 U3293 ( .A(n3064), .Z(n4497) );
  HS65_LH_NOR2X6 U3294 ( .A(n3096), .B(n3101), .Z(n3064) );
  HS65_LH_BFX9 U3295 ( .A(n2681), .Z(n4592) );
  HS65_LH_BFX9 U3296 ( .A(b[27]), .Z(n4670) );
  HS65_LH_BFX9 U3297 ( .A(b[19]), .Z(n4654) );
  HS65_LH_BFX9 U3298 ( .A(b[15]), .Z(n4646) );
  HS65_LH_BFX9 U3299 ( .A(b[4]), .Z(n4624) );
  HS65_LH_BFX9 U3300 ( .A(b[5]), .Z(n4626) );
  HS65_LH_BFX9 U3301 ( .A(b[17]), .Z(n4650) );
  HS65_LH_BFX9 U3302 ( .A(b[7]), .Z(n4630) );
  HS65_LH_BFX9 U3303 ( .A(b[11]), .Z(n4638) );
  HS65_LH_BFX9 U3304 ( .A(b[21]), .Z(n4658) );
  HS65_LH_BFX9 U3305 ( .A(b[9]), .Z(n4634) );
  HS65_LH_BFX9 U3306 ( .A(b[28]), .Z(n4672) );
  HS65_LH_BFX9 U3307 ( .A(b[25]), .Z(n4666) );
  HS65_LH_BFX9 U3308 ( .A(b[18]), .Z(n4652) );
  HS65_LH_BFX9 U3309 ( .A(b[26]), .Z(n4668) );
  HS65_LH_BFX9 U3310 ( .A(b[13]), .Z(n4642) );
  HS65_LH_BFX9 U3311 ( .A(b[24]), .Z(n4664) );
  HS65_LH_BFX9 U3312 ( .A(b[20]), .Z(n4656) );
  HS65_LH_BFX9 U3313 ( .A(b[6]), .Z(n4628) );
  HS65_LH_BFX9 U3314 ( .A(b[10]), .Z(n4636) );
  HS65_LH_BFX9 U3315 ( .A(b[8]), .Z(n4632) );
  HS65_LH_BFX9 U3316 ( .A(b[16]), .Z(n4648) );
  HS65_LH_BFX9 U3317 ( .A(b[12]), .Z(n4640) );
  HS65_LH_BFX9 U3318 ( .A(b[14]), .Z(n4644) );
  HS65_LH_BFX9 U3319 ( .A(n2670), .Z(n4610) );
  HS65_LH_BFX9 U3320 ( .A(b[27]), .Z(n4671) );
  HS65_LH_BFX9 U3321 ( .A(b[19]), .Z(n4655) );
  HS65_LH_BFX9 U3322 ( .A(b[25]), .Z(n4667) );
  HS65_LH_BFX9 U3323 ( .A(b[15]), .Z(n4647) );
  HS65_LH_BFX9 U3324 ( .A(b[4]), .Z(n4625) );
  HS65_LH_BFX9 U3325 ( .A(b[5]), .Z(n4627) );
  HS65_LH_BFX9 U3326 ( .A(b[17]), .Z(n4651) );
  HS65_LH_BFX9 U3327 ( .A(b[7]), .Z(n4631) );
  HS65_LH_BFX9 U3328 ( .A(b[11]), .Z(n4639) );
  HS65_LH_BFX9 U3329 ( .A(b[21]), .Z(n4659) );
  HS65_LH_BFX9 U3330 ( .A(b[12]), .Z(n4641) );
  HS65_LH_BFX9 U3331 ( .A(b[9]), .Z(n4635) );
  HS65_LH_BFX9 U3332 ( .A(b[28]), .Z(n4673) );
  HS65_LH_BFX9 U3333 ( .A(b[13]), .Z(n4643) );
  HS65_LH_BFX9 U3334 ( .A(b[18]), .Z(n4653) );
  HS65_LH_BFX9 U3335 ( .A(b[26]), .Z(n4669) );
  HS65_LH_BFX9 U3336 ( .A(b[24]), .Z(n4665) );
  HS65_LH_BFX9 U3337 ( .A(b[20]), .Z(n4657) );
  HS65_LH_BFX9 U3338 ( .A(b[14]), .Z(n4645) );
  HS65_LH_BFX9 U3339 ( .A(b[6]), .Z(n4629) );
  HS65_LH_BFX9 U3340 ( .A(b[10]), .Z(n4637) );
  HS65_LH_BFX9 U3341 ( .A(b[8]), .Z(n4633) );
  HS65_LH_BFX9 U3342 ( .A(b[16]), .Z(n4649) );
  HS65_LH_BFX9 U3343 ( .A(n4593), .Z(n4594) );
  HS65_LH_BFX9 U3344 ( .A(n4597), .Z(n4598) );
  HS65_LH_BFX9 U3345 ( .A(n4593), .Z(n4595) );
  HS65_LH_BFX9 U3346 ( .A(n4605), .Z(n4606) );
  HS65_LH_BFX9 U3347 ( .A(n4597), .Z(n4599) );
  HS65_LH_BFX9 U3348 ( .A(n4605), .Z(n4607) );
  HS65_LH_BFX9 U3349 ( .A(n4597), .Z(n4600) );
  HS65_LH_BFX9 U3350 ( .A(n4605), .Z(n4608) );
  HS65_LH_BFX9 U3351 ( .A(n4593), .Z(n4596) );
  HS65_LHS_XOR3X2 U3352 ( .A(n292), .B(n227), .C(n2669), .Z(product[63]) );
  HS65_LH_AO22X9 U3353 ( .A(n4678), .B(n4610), .C(n4490), .D(n1006), .Z(n2669)
         );
  HS65_LHS_XOR2X6 U3354 ( .A(n4706), .B(a[30]), .Z(n3103) );
  HS65_LHS_XOR2X6 U3355 ( .A(n4685), .B(a[9]), .Z(n2838) );
  HS65_LHS_XOR2X6 U3356 ( .A(n4691), .B(a[15]), .Z(n2924) );
  HS65_LHS_XOR2X6 U3357 ( .A(n4680), .B(a[3]), .Z(n2753) );
  HS65_LHS_XOR2X6 U3358 ( .A(n4695), .B(a[18]), .Z(n2967) );
  HS65_LHS_XOR2X6 U3359 ( .A(n4688), .B(a[12]), .Z(n2881) );
  HS65_LHS_XOR2X6 U3360 ( .A(n4697), .B(a[21]), .Z(n3010) );
  HS65_LHS_XOR2X6 U3361 ( .A(n4703), .B(a[27]), .Z(n3096) );
  HS65_LHS_XOR2X6 U3362 ( .A(n4700), .B(a[24]), .Z(n3053) );
  HS65_LHS_XOR2X6 U3363 ( .A(n19), .B(a[6]), .Z(n2796) );
  HS65_LHS_XOR2X6 U3364 ( .A(n4681), .B(a[1]), .Z(n2711) );
  HS65_LHS_XNOR2X6 U3365 ( .A(n31), .B(a[7]), .Z(n2797) );
  HS65_LHS_XNOR2X6 U3366 ( .A(n55), .B(a[13]), .Z(n2882) );
  HS65_LHS_XNOR2X6 U3367 ( .A(n43), .B(a[10]), .Z(n2839) );
  HS65_LHS_XNOR2X6 U3368 ( .A(n67), .B(a[16]), .Z(n2925) );
  HS65_LHS_XNOR2X6 U3369 ( .A(n79), .B(a[19]), .Z(n2968) );
  HS65_LHS_XNOR2X6 U3370 ( .A(n103), .B(a[25]), .Z(n3054) );
  HS65_LHS_XNOR2X6 U3371 ( .A(n115), .B(a[28]), .Z(n3097) );
  HS65_LHS_XNOR2X6 U3372 ( .A(n91), .B(a[22]), .Z(n3011) );
  HS65_LHS_XNOR2X6 U3373 ( .A(n19), .B(a[4]), .Z(n2754) );
  HS65_LHS_XOR2X6 U3374 ( .A(a[31]), .B(a[30]), .Z(n3104) );
  HS65_LHS_XNOR2X6 U3375 ( .A(a[4]), .B(a[3]), .Z(n2758) );
  HS65_LHS_XNOR2X6 U3376 ( .A(a[7]), .B(a[6]), .Z(n2801) );
  HS65_LHS_XNOR2X6 U3377 ( .A(a[9]), .B(a[10]), .Z(n2843) );
  HS65_LHS_XNOR2X6 U3378 ( .A(a[13]), .B(a[12]), .Z(n2886) );
  HS65_LHS_XNOR2X6 U3379 ( .A(a[16]), .B(a[15]), .Z(n2929) );
  HS65_LHS_XNOR2X6 U3380 ( .A(a[19]), .B(a[18]), .Z(n2972) );
  HS65_LHS_XNOR2X6 U3381 ( .A(a[22]), .B(a[21]), .Z(n3015) );
  HS65_LHS_XNOR2X6 U3382 ( .A(a[25]), .B(a[24]), .Z(n3058) );
  HS65_LHS_XNOR2X6 U3383 ( .A(a[28]), .B(a[27]), .Z(n3101) );
  HS65_LH_NAND2X7 U3384 ( .A(a[0]), .B(n2711), .Z(n2713) );
  HS65_LH_NAND2X7 U3385 ( .A(a[31]), .B(n3103), .Z(n2673) );
  HS65_LH_BFX9 U3386 ( .A(n2677), .Z(n4597) );
  HS65_LH_NOR2AX3 U3387 ( .A(a[0]), .B(n2711), .Z(n2677) );
  HS65_LH_BFX9 U3388 ( .A(n2671), .Z(n4605) );
  HS65_LH_NOR2AX3 U3389 ( .A(n3103), .B(a[31]), .Z(n2671) );
  HS65_LH_BFX9 U3390 ( .A(n2679), .Z(n4593) );
  HS65_LH_NOR2AX3 U3391 ( .A(a[1]), .B(a[0]), .Z(n2679) );
endmodule


module alu ( clk, rst_n, .alu_i({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , 
        \alu_i[SRC_B][31] , \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , 
        \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , 
        \alu_i[SRC_B][25] , \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , 
        \alu_i[SRC_B][22] , \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , 
        \alu_i[SRC_B][19] , \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , 
        \alu_i[SRC_B][16] , \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , 
        \alu_i[SRC_B][13] , \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , 
        \alu_i[SRC_B][10] , \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , 
        \alu_i[SRC_B][7] , \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , 
        \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , 
        \alu_i[SRC_B][1] , \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , 
        \alu_i[OP][2] , \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , 
        \alu_i[SHAMT][3] , \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , 
        \alu_i[SHAMT][0] }), .alu_o({\alu_o[BRANCH] , \alu_o[RESULT][31] , 
        \alu_o[RESULT][30] , \alu_o[RESULT][29] , \alu_o[RESULT][28] , 
        \alu_o[RESULT][27] , \alu_o[RESULT][26] , \alu_o[RESULT][25] , 
        \alu_o[RESULT][24] , \alu_o[RESULT][23] , \alu_o[RESULT][22] , 
        \alu_o[RESULT][21] , \alu_o[RESULT][20] , \alu_o[RESULT][19] , 
        \alu_o[RESULT][18] , \alu_o[RESULT][17] , \alu_o[RESULT][16] , 
        \alu_o[RESULT][15] , \alu_o[RESULT][14] , \alu_o[RESULT][13] , 
        \alu_o[RESULT][12] , \alu_o[RESULT][11] , \alu_o[RESULT][10] , 
        \alu_o[RESULT][9] , \alu_o[RESULT][8] , \alu_o[RESULT][7] , 
        \alu_o[RESULT][6] , \alu_o[RESULT][5] , \alu_o[RESULT][4] , 
        \alu_o[RESULT][3] , \alu_o[RESULT][2] , \alu_o[RESULT][1] , 
        \alu_o[RESULT][0] }) );
  input clk, rst_n, \alu_i[SRC_A][31] , \alu_i[SRC_A][30] , \alu_i[SRC_A][29] ,
         \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , \alu_i[SRC_A][26] ,
         \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , \alu_i[SRC_A][23] ,
         \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , \alu_i[SRC_A][20] ,
         \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , \alu_i[SRC_A][17] ,
         \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , \alu_i[SRC_A][14] ,
         \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , \alu_i[SRC_A][11] ,
         \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , \alu_i[SRC_A][8] ,
         \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , \alu_i[SRC_A][5] ,
         \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , \alu_i[SRC_A][2] ,
         \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , \alu_i[SRC_B][31] ,
         \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , \alu_i[SRC_B][28] ,
         \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , \alu_i[SRC_B][25] ,
         \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , \alu_i[SRC_B][22] ,
         \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , \alu_i[SRC_B][19] ,
         \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , \alu_i[SRC_B][16] ,
         \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , \alu_i[SRC_B][13] ,
         \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , \alu_i[SRC_B][10] ,
         \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , \alu_i[SRC_B][7] ,
         \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , \alu_i[SRC_B][4] ,
         \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , \alu_i[SRC_B][1] ,
         \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , \alu_i[OP][2] ,
         \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , \alu_i[SHAMT][3] ,
         \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , \alu_i[SHAMT][0] ;
  output \alu_o[BRANCH] , \alu_o[RESULT][31] , \alu_o[RESULT][30] ,
         \alu_o[RESULT][29] , \alu_o[RESULT][28] , \alu_o[RESULT][27] ,
         \alu_o[RESULT][26] , \alu_o[RESULT][25] , \alu_o[RESULT][24] ,
         \alu_o[RESULT][23] , \alu_o[RESULT][22] , \alu_o[RESULT][21] ,
         \alu_o[RESULT][20] , \alu_o[RESULT][19] , \alu_o[RESULT][18] ,
         \alu_o[RESULT][17] , \alu_o[RESULT][16] , \alu_o[RESULT][15] ,
         \alu_o[RESULT][14] , \alu_o[RESULT][13] , \alu_o[RESULT][12] ,
         \alu_o[RESULT][11] , \alu_o[RESULT][10] , \alu_o[RESULT][9] ,
         \alu_o[RESULT][8] , \alu_o[RESULT][7] , \alu_o[RESULT][6] ,
         \alu_o[RESULT][5] , \alu_o[RESULT][4] , \alu_o[RESULT][3] ,
         \alu_o[RESULT][2] , \alu_o[RESULT][1] , \alu_o[RESULT][0] ;
  wire   \HI_LO_c[HI][31] , \HI_LO_c[HI][30] , \HI_LO_c[HI][29] ,
         \HI_LO_c[HI][28] , \HI_LO_c[HI][27] , \HI_LO_c[HI][26] ,
         \HI_LO_c[HI][25] , \HI_LO_c[HI][24] , \HI_LO_c[HI][23] ,
         \HI_LO_c[HI][22] , \HI_LO_c[HI][21] , \HI_LO_c[HI][20] ,
         \HI_LO_c[HI][19] , \HI_LO_c[HI][18] , \HI_LO_c[HI][17] ,
         \HI_LO_c[HI][16] , \HI_LO_c[HI][15] , \HI_LO_c[HI][14] ,
         \HI_LO_c[HI][13] , \HI_LO_c[HI][12] , \HI_LO_c[HI][11] ,
         \HI_LO_c[HI][10] , \HI_LO_c[HI][9] , \HI_LO_c[HI][8] ,
         \HI_LO_c[HI][7] , \HI_LO_c[HI][6] , \HI_LO_c[HI][5] ,
         \HI_LO_c[HI][4] , \HI_LO_c[HI][3] , \HI_LO_c[HI][2] ,
         \HI_LO_c[HI][1] , \HI_LO_c[HI][0] , \HI_LO_c[LO][31] ,
         \HI_LO_c[LO][30] , \HI_LO_c[LO][29] , \HI_LO_c[LO][28] ,
         \HI_LO_c[LO][27] , \HI_LO_c[LO][26] , \HI_LO_c[LO][25] ,
         \HI_LO_c[LO][24] , \HI_LO_c[LO][23] , \HI_LO_c[LO][22] ,
         \HI_LO_c[LO][21] , \HI_LO_c[LO][20] , \HI_LO_c[LO][19] ,
         \HI_LO_c[LO][18] , \HI_LO_c[LO][17] , \HI_LO_c[LO][16] ,
         \HI_LO_c[LO][15] , \HI_LO_c[LO][14] , \HI_LO_c[LO][13] ,
         \HI_LO_c[LO][12] , \HI_LO_c[LO][11] , \HI_LO_c[LO][10] ,
         \HI_LO_c[LO][9] , \HI_LO_c[LO][8] , \HI_LO_c[LO][7] ,
         \HI_LO_c[LO][6] , \HI_LO_c[LO][5] , \HI_LO_c[LO][4] ,
         \HI_LO_c[LO][3] , \HI_LO_c[LO][2] , \HI_LO_c[LO][1] ,
         \HI_LO_c[LO][0] , N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N647, N648,
         N713, N714, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801;

  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][31]  ( .D(n525), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][30]  ( .D(n524), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][29]  ( .D(n523), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][28]  ( .D(n522), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][27]  ( .D(n521), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][26]  ( .D(n520), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][25]  ( .D(n519), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][24]  ( .D(n518), .CP(clk), .RN(n1748), .Q(
        \HI_LO_c[HI][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][23]  ( .D(n517), .CP(clk), .RN(n1748), .Q(
        \HI_LO_c[HI][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][22]  ( .D(n516), .CP(clk), .RN(n1748), .Q(
        \HI_LO_c[HI][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][21]  ( .D(n515), .CP(clk), .RN(n1748), .Q(
        \HI_LO_c[HI][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][20]  ( .D(n514), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][19]  ( .D(n513), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][18]  ( .D(n512), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][17]  ( .D(n511), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][16]  ( .D(n510), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][15]  ( .D(n509), .CP(clk), .RN(n1747), .Q(
        \HI_LO_c[HI][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][14]  ( .D(n508), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][13]  ( .D(n507), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][12]  ( .D(n506), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][11]  ( .D(n505), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][10]  ( .D(n504), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][9]  ( .D(n503), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][8]  ( .D(n502), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][7]  ( .D(n501), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][6]  ( .D(n500), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][5]  ( .D(n499), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[HI][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][4]  ( .D(n498), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][3]  ( .D(n497), .CP(clk), .RN(n1746), .Q(
        \HI_LO_c[HI][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][2]  ( .D(n496), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[HI][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][1]  ( .D(n495), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[HI][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][0]  ( .D(n494), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[HI][0] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][31]  ( .D(n493), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][30]  ( .D(n492), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][29]  ( .D(n491), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][28]  ( .D(n490), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][27]  ( .D(n489), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][26]  ( .D(n488), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][25]  ( .D(n487), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][24]  ( .D(n486), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][23]  ( .D(n485), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][22]  ( .D(n484), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][21]  ( .D(n483), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][20]  ( .D(n482), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][19]  ( .D(n481), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][18]  ( .D(n480), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][17]  ( .D(n479), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][16]  ( .D(n478), .CP(clk), .RN(n1744), .Q(
        \HI_LO_c[LO][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][15]  ( .D(n477), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][14]  ( .D(n476), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][13]  ( .D(n475), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][12]  ( .D(n474), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][11]  ( .D(n473), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][10]  ( .D(n472), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][9]  ( .D(n471), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][8]  ( .D(n470), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][7]  ( .D(n469), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][6]  ( .D(n468), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][5]  ( .D(n467), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][4]  ( .D(n466), .CP(clk), .RN(n1743), .Q(
        \HI_LO_c[LO][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][3]  ( .D(n465), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][2]  ( .D(n464), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][1]  ( .D(n463), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][0]  ( .D(n462), .CP(clk), .RN(n1745), .Q(
        \HI_LO_c[LO][0] ) );
  alu_DW_cmp_0 lt_136 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n1731, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({\alu_i[SRC_B][31] , 
        \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , n1727, n1726, n1725, n1724, 
        n1723, \alu_i[SRC_B][23] , \alu_i[SRC_B][22] , n1720, n1719, n1718, 
        n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, 
        n1707, n1706, n1705, n1704, n1703, \alu_i[SRC_B][3] , 
        \alu_i[SRC_B][2] , \alu_i[SRC_B][1] , \alu_i[SRC_B][0] }), .TC(1'b1), 
        .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N647) );
  alu_DW01_sub_0 sub_68 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n1731, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({\alu_i[SRC_B][31] , 
        \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , n1727, n1726, n1725, n1724, 
        n1723, \alu_i[SRC_B][23] , \alu_i[SRC_B][22] , n1720, n1719, n1718, 
        n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, 
        n1707, n1706, n1705, n1704, n1703, \alu_i[SRC_B][3] , 
        \alu_i[SRC_B][2] , \alu_i[SRC_B][1] , \alu_i[SRC_B][0] }), .CI(1'b0), 
        .DIFF({N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, 
        N139, N138, N137, N136, N135, N134, N133, N132, N131, N130}) );
  alu_DW01_cmp6_0 r325 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n1731, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({\alu_i[SRC_B][31] , 
        \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , n1727, n1726, n1725, n1724, 
        n1723, \alu_i[SRC_B][23] , \alu_i[SRC_B][22] , n1720, n1719, n1718, 
        n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, 
        n1707, n1706, n1705, n1704, n1703, \alu_i[SRC_B][3] , 
        \alu_i[SRC_B][2] , \alu_i[SRC_B][1] , \alu_i[SRC_B][0] }), .TC(1'b0), 
        .LT(N648), .EQ(N713), .NE(N714) );
  alu_DW01_add_0 r321 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n1731, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({\alu_i[SRC_B][31] , 
        \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , n1727, n1726, n1725, n1724, 
        n1723, \alu_i[SRC_B][23] , \alu_i[SRC_B][22] , n1720, n1719, n1718, 
        n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, 
        n1707, n1706, n1705, n1704, n1703, \alu_i[SRC_B][3] , 
        \alu_i[SRC_B][2] , \alu_i[SRC_B][1] , \alu_i[SRC_B][0] }), .CI(1'b0), 
        .SUM({N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98}) );
  alu_DW_mult_uns_0 mult_71 ( .a({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n1731, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .b({\alu_i[SRC_B][31] , 
        \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , n1727, n1726, n1725, n1724, 
        n1723, \alu_i[SRC_B][23] , \alu_i[SRC_B][22] , n1720, n1719, n1718, 
        n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, 
        n1707, n1706, n1705, n1704, n1703, \alu_i[SRC_B][3] , 
        \alu_i[SRC_B][2] , \alu_i[SRC_B][1] , \alu_i[SRC_B][0] }), .product({
        N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, 
        N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, 
        N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, 
        N165, N164, N163, N162}) );
  HS65_LH_IVX9 U7 ( .A(n421), .Z(n1641) );
  HS65_LH_IVX9 U8 ( .A(n317), .Z(n1642) );
  HS65_LH_NAND4ABX3 U9 ( .A(n87), .B(n88), .C(n89), .D(n90), .Z(n86) );
  HS65_LH_BFX9 U10 ( .A(\alu_i[SRC_B][19] ), .Z(n1718) );
  HS65_LH_BFX9 U11 ( .A(\alu_i[SRC_B][27] ), .Z(n1726) );
  HS65_LH_BFX9 U12 ( .A(\alu_i[SRC_B][26] ), .Z(n1725) );
  HS65_LH_BFX9 U13 ( .A(\alu_i[SRC_B][10] ), .Z(n1709) );
  HS65_LH_BFX9 U14 ( .A(\alu_i[SRC_B][12] ), .Z(n1711) );
  HS65_LH_BFX9 U15 ( .A(\alu_i[SRC_B][13] ), .Z(n1712) );
  HS65_LH_BFX9 U16 ( .A(\alu_i[SRC_B][14] ), .Z(n1713) );
  HS65_LH_BFX9 U17 ( .A(\alu_i[SRC_B][16] ), .Z(n1715) );
  HS65_LH_BFX9 U18 ( .A(\alu_i[SRC_B][17] ), .Z(n1716) );
  HS65_LH_BFX9 U19 ( .A(\alu_i[SRC_B][18] ), .Z(n1717) );
  HS65_LH_BFX9 U20 ( .A(\alu_i[SRC_B][20] ), .Z(n1719) );
  HS65_LH_BFX9 U21 ( .A(\alu_i[SRC_B][21] ), .Z(n1720) );
  HS65_LH_BFX9 U22 ( .A(\alu_i[SRC_B][24] ), .Z(n1723) );
  HS65_LH_BFX9 U23 ( .A(\alu_i[SRC_B][25] ), .Z(n1724) );
  HS65_LH_BFX9 U24 ( .A(\alu_i[SRC_B][11] ), .Z(n1710) );
  HS65_LH_BFX9 U25 ( .A(\alu_i[SRC_B][28] ), .Z(n1727) );
  HS65_LH_BFX9 U26 ( .A(\alu_i[SRC_B][15] ), .Z(n1714) );
  HS65_LH_BFX9 U27 ( .A(\alu_i[SRC_B][4] ), .Z(n1703) );
  HS65_LH_BFX9 U28 ( .A(\alu_i[SRC_B][6] ), .Z(n1705) );
  HS65_LH_BFX9 U29 ( .A(\alu_i[SRC_B][7] ), .Z(n1706) );
  HS65_LH_BFX9 U30 ( .A(\alu_i[SRC_B][5] ), .Z(n1704) );
  HS65_LH_BFX9 U31 ( .A(\alu_i[SRC_B][8] ), .Z(n1707) );
  HS65_LH_BFX9 U32 ( .A(\alu_i[SRC_B][9] ), .Z(n1708) );
  HS65_LH_IVX9 U33 ( .A(n1686), .Z(n1685) );
  HS65_LH_IVX9 U34 ( .A(n1686), .Z(n1684) );
  HS65_LH_IVX9 U35 ( .A(n1694), .Z(n1689) );
  HS65_LH_IVX9 U36 ( .A(n1694), .Z(n1690) );
  HS65_LH_IVX9 U37 ( .A(n1694), .Z(n1691) );
  HS65_LH_IVX9 U38 ( .A(n1693), .Z(n1692) );
  HS65_LH_AOI12X2 U39 ( .A(n1651), .B(n1642), .C(n1682), .Z(n235) );
  HS65_LH_AOI12X2 U40 ( .A(n1651), .B(n1641), .C(n1682), .Z(n206) );
  HS65_LH_IVX9 U41 ( .A(n421), .Z(n1751) );
  HS65_LH_IVX9 U42 ( .A(n317), .Z(n1749) );
  HS65_LH_IVX9 U43 ( .A(n1682), .Z(n1680) );
  HS65_LH_IVX9 U44 ( .A(n1682), .Z(n1681) );
  HS65_LH_BFX9 U45 ( .A(n1687), .Z(n1694) );
  HS65_LH_BFX9 U46 ( .A(n1687), .Z(n1693) );
  HS65_LH_BFX9 U47 ( .A(n1793), .Z(n1663) );
  HS65_LH_BFX9 U48 ( .A(n1793), .Z(n1662) );
  HS65_LH_BFX9 U49 ( .A(n1795), .Z(n1665) );
  HS65_LH_BFX9 U50 ( .A(n1792), .Z(n1660) );
  HS65_LH_BFX9 U51 ( .A(n1792), .Z(n1661) );
  HS65_LH_IVX9 U52 ( .A(n1683), .Z(n1686) );
  HS65_LH_BFX9 U53 ( .A(n1687), .Z(n1695) );
  HS65_LH_BFX9 U54 ( .A(n1688), .Z(n1696) );
  HS65_LH_BFX9 U55 ( .A(n1688), .Z(n1697) );
  HS65_LH_BFX9 U56 ( .A(n1795), .Z(n1666) );
  HS65_LH_BFX9 U57 ( .A(n1793), .Z(n1664) );
  HS65_LH_BFX9 U58 ( .A(n1688), .Z(n1698) );
  HS65_LH_IVX9 U59 ( .A(n94), .Z(n1793) );
  HS65_LH_IVX9 U60 ( .A(n96), .Z(n1792) );
  HS65_LH_IVX9 U61 ( .A(n91), .Z(n1795) );
  HS65_LH_AND2X4 U62 ( .A(n379), .B(n1799), .Z(n211) );
  HS65_LH_NAND2X7 U63 ( .A(n1752), .B(n1756), .Z(n421) );
  HS65_LH_NOR2AX3 U64 ( .A(n1670), .B(n421), .Z(n204) );
  HS65_LH_NAND2X7 U65 ( .A(n1750), .B(n1756), .Z(n317) );
  HS65_LH_NOR4ABX2 U66 ( .A(n91), .B(n92), .C(n1672), .D(n93), .Z(n90) );
  HS65_LH_NAND3X5 U67 ( .A(n94), .B(n1679), .C(n96), .Z(n93) );
  HS65_LH_BFX9 U68 ( .A(n92), .Z(n1683) );
  HS65_LH_NAND2X7 U69 ( .A(n97), .B(n1799), .Z(n92) );
  HS65_LH_IVX9 U70 ( .A(n1672), .Z(n1671) );
  HS65_LH_IVX9 U71 ( .A(n119), .Z(n1672) );
  HS65_LH_BFX9 U72 ( .A(n98), .Z(n1677) );
  HS65_LH_BFX9 U73 ( .A(n1768), .Z(n1651) );
  HS65_LH_IVX9 U74 ( .A(n1679), .Z(n1682) );
  HS65_LH_BFX9 U75 ( .A(n1768), .Z(n1652) );
  HS65_LH_IVX9 U76 ( .A(n101), .Z(n1798) );
  HS65_LH_BFX9 U77 ( .A(n98), .Z(n1678) );
  HS65_LH_BFX9 U78 ( .A(n86), .Z(n1687) );
  HS65_LH_BFX9 U79 ( .A(n86), .Z(n1688) );
  HS65_LH_BFX9 U80 ( .A(n1768), .Z(n1653) );
  HS65_LH_BFX9 U81 ( .A(n1654), .Z(n1656) );
  HS65_LH_BFX9 U82 ( .A(n1655), .Z(n1658) );
  HS65_LH_BFX9 U83 ( .A(n1654), .Z(n1657) );
  HS65_LH_BFX9 U84 ( .A(n1655), .Z(n1659) );
  HS65_LH_CB4I6X9 U85 ( .A(n1799), .B(n99), .C(n1794), .D(n1676), .Z(n88) );
  HS65_LH_AOI13X5 U86 ( .A(n101), .B(n102), .C(n103), .D(n1796), .Z(n87) );
  HS65_LH_AOI12X2 U87 ( .A(n97), .B(n1798), .C(n1677), .Z(n89) );
  HS65_LH_NAND3X5 U88 ( .A(n432), .B(n1801), .C(n433), .Z(n119) );
  HS65_LH_IVX9 U89 ( .A(n396), .Z(n1768) );
  HS65_LH_NOR2X6 U90 ( .A(n1801), .B(n1797), .Z(n97) );
  HS65_LH_AO32X4 U91 ( .A(n104), .B(n1801), .C(n432), .D(n1798), .E(n379), .Z(
        n98) );
  HS65_LH_AOI222X2 U92 ( .A(n1751), .B(n194), .C(n111), .D(n130), .E(n1643), 
        .F(n131), .Z(n185) );
  HS65_LH_AOI222X2 U93 ( .A(n109), .B(n110), .C(n111), .D(n112), .E(n1644), 
        .F(n114), .Z(n108) );
  HS65_LH_AOI222X2 U94 ( .A(n275), .B(n182), .C(n214), .D(n181), .E(n211), .F(
        \alu_i[SRC_B][1] ), .Z(n368) );
  HS65_LH_AOI222X2 U95 ( .A(n275), .B(n160), .C(n214), .D(n161), .E(n211), .F(
        \alu_i[SRC_B][2] ), .Z(n361) );
  HS65_LH_AOI222X2 U96 ( .A(n275), .B(n144), .C(n214), .D(n142), .E(n211), .F(
        \alu_i[SRC_B][3] ), .Z(n354) );
  HS65_LH_AOI222X2 U97 ( .A(n1754), .B(n241), .C(n1643), .D(n166), .E(
        \alu_i[SRC_B][3] ), .F(n200), .Z(n240) );
  HS65_LH_AOI222X2 U98 ( .A(n111), .B(n114), .C(n1751), .D(n177), .E(n122), 
        .F(n112), .Z(n176) );
  HS65_LH_AOI212X4 U99 ( .A(n120), .B(n168), .C(n1751), .D(n171), .E(n420), 
        .Z(n415) );
  HS65_LH_AO22X9 U100 ( .A(n160), .B(n212), .C(n172), .D(n111), .Z(n420) );
  HS65_LH_AOI212X4 U101 ( .A(n273), .B(n142), .C(n212), .D(n215), .E(n274), 
        .Z(n268) );
  HS65_LH_AO22X9 U102 ( .A(n213), .B(n145), .C(n216), .D(n1749), .Z(n274) );
  HS65_LH_AOI212X4 U103 ( .A(n145), .B(n160), .C(n1749), .D(n161), .E(n162), 
        .Z(n159) );
  HS65_LH_AO22X9 U104 ( .A(n163), .B(n120), .C(n164), .D(n109), .Z(n162) );
  HS65_LH_AOI212X4 U105 ( .A(n120), .B(n141), .C(n1749), .D(n142), .E(n143), 
        .Z(n140) );
  HS65_LH_AO22X9 U106 ( .A(n144), .B(n1645), .C(n146), .D(n113), .Z(n143) );
  HS65_LH_IVX9 U107 ( .A(n434), .Z(n1752) );
  HS65_LH_IVX9 U108 ( .A(n190), .Z(n1750) );
  HS65_LH_AND2X4 U109 ( .A(n364), .B(n1750), .Z(n214) );
  HS65_LH_MX41X7 U110 ( .D0(\alu_i[SRC_B][3] ), .S0(n1652), .D1(
        \alu_i[SRC_B][2] ), .S1(n1649), .D2(n1656), .S2(\alu_i[SRC_B][1] ), 
        .D3(n1668), .S3(\alu_i[SRC_B][0] ), .Z(n144) );
  HS65_LH_NAND3X5 U111 ( .A(n1794), .B(n1801), .C(n104), .Z(n96) );
  HS65_LH_AND2X4 U112 ( .A(n364), .B(n1752), .Z(n122) );
  HS65_LH_NOR2X6 U113 ( .A(n1801), .B(n427), .Z(n379) );
  HS65_LH_NAND3X5 U114 ( .A(n433), .B(n1801), .C(n1794), .Z(n94) );
  HS65_LH_NOR2X6 U115 ( .A(n433), .B(n99), .Z(n101) );
  HS65_LH_IVX9 U116 ( .A(n307), .Z(n1756) );
  HS65_LH_IVX9 U117 ( .A(n102), .Z(n1799) );
  HS65_LH_MX41X7 U118 ( .D0(n1757), .S0(n164), .D1(n364), .S1(n168), .D2(n1756), .S2(n172), .D3(n1759), .S3(n163), .Z(n241) );
  HS65_LH_MX41X7 U119 ( .D0(n1757), .S0(n136), .D1(n1759), .S1(n132), .D2(n364), .S2(n129), .D3(n1756), .S3(n128), .Z(n375) );
  HS65_LH_MX41X7 U120 ( .D0(n1756), .S0(n297), .D1(n1757), .S1(n296), .D2(
        n1759), .S2(n181), .D3(n364), .S3(n182), .Z(n254) );
  HS65_LH_NAND2X7 U121 ( .A(n104), .B(n379), .Z(n91) );
  HS65_LH_MX41X7 U122 ( .D0(n364), .S0(n144), .D1(n1757), .S1(n276), .D2(n1759), .S2(n142), .D3(n1756), .S3(n277), .Z(n224) );
  HS65_LH_MX41X7 U123 ( .D0(n364), .S0(n121), .D1(n1757), .S1(n123), .D2(n1759), .S2(n110), .D3(n1756), .S3(n112), .Z(n350) );
  HS65_LH_MX41X7 U124 ( .D0(n1757), .S0(n288), .D1(n364), .S1(n160), .D2(n1759), .S2(n161), .D3(n1756), .S3(n283), .Z(n236) );
  HS65_LH_OAI21X3 U125 ( .A(\alu_i[SRC_B][29] ), .B(n1685), .C(n1680), .Z(n253) );
  HS65_LH_OAI21X3 U126 ( .A(\alu_i[SRC_B][30] ), .B(n1685), .C(n1680), .Z(n234) );
  HS65_LH_OAI21X3 U127 ( .A(\alu_i[SRC_B][31] ), .B(n1685), .C(n1680), .Z(n219) );
  HS65_LH_AO222X4 U128 ( .A(n123), .B(n1756), .C(n110), .D(n1757), .E(n121), 
        .F(n1759), .Z(n178) );
  HS65_LH_AO222X4 U129 ( .A(n181), .B(n1757), .C(n182), .D(n1759), .E(n296), 
        .F(n1756), .Z(n116) );
  HS65_LH_IVX9 U130 ( .A(n427), .Z(n1794) );
  HS65_LH_BFX9 U131 ( .A(n95), .Z(n1679) );
  HS65_LH_NAND2X7 U132 ( .A(n97), .B(n104), .Z(n95) );
  HS65_LH_IVX9 U133 ( .A(n432), .Z(n1797) );
  HS65_LH_BFX9 U134 ( .A(n1673), .Z(n1674) );
  HS65_LH_IVX9 U135 ( .A(n343), .Z(n1762) );
  HS65_LH_BFX9 U136 ( .A(n1673), .Z(n1675) );
  HS65_LH_BFX9 U137 ( .A(n1770), .Z(n1655) );
  HS65_LH_BFX9 U138 ( .A(n1770), .Z(n1654) );
  HS65_LH_BFX9 U139 ( .A(n1667), .Z(n1669) );
  HS65_LH_BFX9 U140 ( .A(n1667), .Z(n1668) );
  HS65_LH_BFX9 U141 ( .A(n1667), .Z(n1670) );
  HS65_LH_BFX9 U142 ( .A(n1767), .Z(n1647) );
  HS65_LH_AO22X9 U143 ( .A(n163), .B(n109), .C(n161), .D(n1646), .Z(n419) );
  HS65_LH_BFX9 U144 ( .A(n1767), .Z(n1649) );
  HS65_LH_BFX9 U145 ( .A(n1767), .Z(n1650) );
  HS65_LH_BFX9 U146 ( .A(n1767), .Z(n1648) );
  HS65_LH_AO22X9 U147 ( .A(n248), .B(n1749), .C(n178), .D(n1752), .Z(n334) );
  HS65_LH_AO22X9 U148 ( .A(n261), .B(n1749), .C(n133), .D(n1755), .Z(n304) );
  HS65_LH_AO22X9 U149 ( .A(n250), .B(n1749), .C(n116), .D(n1755), .Z(n295) );
  HS65_LH_AO12X9 U150 ( .A(n1651), .B(n275), .C(n211), .Z(n377) );
  HS65_LH_BFX9 U151 ( .A(n1673), .Z(n1676) );
  HS65_LH_OAI222X2 U152 ( .A(n221), .B(n1700), .C(n1699), .D(n220), .E(n396), 
        .F(n1701), .Z(n160) );
  HS65_LH_IVX9 U153 ( .A(n221), .Z(n1767) );
  HS65_LH_OAI222X2 U154 ( .A(n221), .B(n1729), .C(n220), .D(n1730), .E(n396), 
        .F(n1728), .Z(n121) );
  HS65_LH_NAND3X5 U155 ( .A(n97), .B(n1753), .C(n99), .Z(n190) );
  HS65_LH_NOR2X6 U156 ( .A(n434), .B(n193), .Z(n111) );
  HS65_LH_OAI22X6 U157 ( .A(n396), .B(n1729), .C(n221), .D(n1730), .Z(n168) );
  HS65_LH_OAI22X6 U158 ( .A(n396), .B(n1700), .C(n221), .D(n1699), .Z(n182) );
  HS65_LH_NAND3X5 U159 ( .A(n433), .B(n1753), .C(n97), .Z(n434) );
  HS65_LH_NOR2X6 U160 ( .A(n190), .B(n193), .Z(n212) );
  HS65_LH_NOR2AX3 U161 ( .A(\alu_i[OP][0] ), .B(n1800), .Z(n433) );
  HS65_LH_NOR2X6 U162 ( .A(n434), .B(n306), .Z(n1643) );
  HS65_LH_NOR2X6 U163 ( .A(n434), .B(n306), .Z(n113) );
  HS65_LH_NOR2X6 U164 ( .A(n434), .B(n306), .Z(n1644) );
  HS65_LH_OAI222X2 U165 ( .A(n1762), .B(n306), .C(n1758), .D(n189), .E(n1764), 
        .F(n307), .Z(n265) );
  HS65_LH_IVX9 U166 ( .A(n310), .Z(n1764) );
  HS65_LH_OAI21X3 U167 ( .A(n221), .B(n421), .C(n96), .Z(n200) );
  HS65_LH_NOR2X6 U168 ( .A(n1761), .B(n1758), .Z(n364) );
  HS65_LH_NOR2X6 U169 ( .A(n192), .B(n306), .Z(n120) );
  HS65_LH_OAI32X5 U170 ( .A(n427), .B(\alu_i[OP][2] ), .C(n428), .D(n429), .E(
        n1791), .Z(n426) );
  HS65_LH_AOI12X2 U171 ( .A(n1686), .B(n1699), .C(n1682), .Z(n429) );
  HS65_LH_AOI22X6 U172 ( .A(N648), .B(n99), .C(N647), .D(n1799), .Z(n428) );
  HS65_LH_NOR2X6 U173 ( .A(n305), .B(n307), .Z(n275) );
  HS65_LH_NOR2X6 U174 ( .A(n190), .B(n306), .Z(n145) );
  HS65_LH_NOR2X6 U175 ( .A(\alu_i[OP][0] ), .B(\alu_i[OP][1] ), .Z(n104) );
  HS65_LH_NOR2X6 U176 ( .A(n190), .B(n306), .Z(n1646) );
  HS65_LH_OAI212X5 U177 ( .A(n1763), .B(n306), .C(n1762), .D(n307), .E(n308), 
        .Z(n133) );
  HS65_LH_IVX9 U178 ( .A(n309), .Z(n1763) );
  HS65_LH_NAND3X5 U179 ( .A(n1651), .B(\alu_i[SRC_B][0] ), .C(n1759), .Z(n308)
         );
  HS65_LH_NOR2X6 U180 ( .A(n190), .B(n306), .Z(n1645) );
  HS65_LH_NOR2X6 U181 ( .A(n305), .B(n306), .Z(n273) );
  HS65_LH_AOI222X2 U182 ( .A(n211), .B(n1711), .C(n212), .D(n259), .E(n214), 
        .F(n260), .Z(n258) );
  HS65_LH_AOI222X2 U183 ( .A(n211), .B(n1712), .C(n212), .D(n248), .E(n214), 
        .F(n249), .Z(n247) );
  HS65_LH_AOI222X2 U184 ( .A(n211), .B(n1713), .C(n212), .D(n229), .E(n214), 
        .F(n230), .Z(n228) );
  HS65_LH_AOI222X2 U185 ( .A(n1754), .B(n199), .C(n1644), .D(n148), .E(n1703), 
        .F(n200), .Z(n198) );
  HS65_LH_NOR2X6 U186 ( .A(n192), .B(n307), .Z(n109) );
  HS65_LH_NAND2X7 U187 ( .A(n1771), .B(n1769), .Z(n396) );
  HS65_LH_NOR2X6 U188 ( .A(n1800), .B(\alu_i[OP][0] ), .Z(n99) );
  HS65_LH_AOI212X4 U189 ( .A(n273), .B(n144), .C(n1646), .D(n215), .E(n315), 
        .Z(n314) );
  HS65_LH_OAI212X5 U190 ( .A(n316), .B(n1722), .C(n1766), .D(n317), .E(n318), 
        .Z(n315) );
  HS65_LH_IVX9 U191 ( .A(n213), .Z(n1766) );
  HS65_LH_CBI4I1X5 U192 ( .A(n1686), .B(n1722), .C(n1682), .D(
        \alu_i[SRC_A][23] ), .Z(n318) );
  HS65_LH_AOI212X4 U193 ( .A(n211), .B(n1703), .C(n212), .D(n310), .E(n342), 
        .Z(n337) );
  HS65_LH_AO22X9 U194 ( .A(n343), .B(n214), .C(n260), .D(n145), .Z(n342) );
  HS65_LH_AOI212X4 U195 ( .A(n273), .B(n161), .C(n212), .D(n230), .E(n282), 
        .Z(n281) );
  HS65_LH_AO22X9 U196 ( .A(n1709), .B(n211), .C(n283), .D(n214), .Z(n282) );
  HS65_LH_NOR2X6 U197 ( .A(n1730), .B(n396), .Z(n150) );
  HS65_LH_AOI212X4 U198 ( .A(\alu_i[SRC_A][23] ), .B(n1672), .C(n1686), .D(
        n1738), .E(n1682), .Z(n316) );
  HS65_LH_IVX9 U199 ( .A(\alu_i[OP][2] ), .Z(n1801) );
  HS65_LH_NAND2X7 U200 ( .A(n1758), .B(n1761), .Z(n307) );
  HS65_LH_OAI212X5 U201 ( .A(\alu_i[SRC_A][20] ), .B(n92), .C(n119), .D(n1737), 
        .E(n1681), .Z(n339) );
  HS65_LH_OAI212X5 U202 ( .A(\alu_i[SRC_A][11] ), .B(n1684), .C(n119), .D(
        n1734), .E(n95), .Z(n410) );
  HS65_LH_MX41X7 U203 ( .D0(n1706), .S0(n1652), .D1(n1705), .S1(n1649), .D2(
        n1704), .S2(n1658), .D3(n1703), .S3(n1669), .Z(n142) );
  HS65_LH_MX41X7 U204 ( .D0(n1705), .S0(n1653), .D1(n1704), .S1(n1650), .D2(
        n1703), .S2(n1658), .D3(\alu_i[SRC_B][3] ), .S3(n1670), .Z(n161) );
  HS65_LH_MX41X7 U205 ( .D0(n1727), .S0(n1653), .D1(\alu_i[SRC_B][29] ), .S1(
        n1650), .D2(\alu_i[SRC_B][30] ), .S2(n1659), .D3(\alu_i[SRC_B][31] ), 
        .S3(n1670), .Z(n129) );
  HS65_LH_OAI212X5 U206 ( .A(n220), .B(n1728), .C(n221), .D(n1729), .E(n222), 
        .Z(n218) );
  HS65_LH_AOI12X2 U207 ( .A(n1727), .B(n1668), .C(n150), .Z(n222) );
  HS65_LH_OAI212X5 U208 ( .A(\alu_i[SRC_A][29] ), .B(n1683), .C(n1671), .D(
        n1740), .E(n235), .Z(n251) );
  HS65_LH_OAI212X5 U209 ( .A(\alu_i[SRC_B][1] ), .B(n92), .C(n119), .D(n1700), 
        .E(n1681), .Z(n348) );
  HS65_LH_OAI212X5 U210 ( .A(\alu_i[SRC_B][2] ), .B(n1683), .C(n1671), .D(
        n1701), .E(n1680), .Z(n242) );
  HS65_LH_OAI212X5 U211 ( .A(\alu_i[SRC_B][3] ), .B(n92), .C(n119), .D(n1702), 
        .E(n1680), .Z(n202) );
  HS65_LH_OAI212X5 U212 ( .A(\alu_i[SRC_A][5] ), .B(n1684), .C(n1671), .D(
        n1732), .E(n1680), .Z(n179) );
  HS65_LH_OAI212X5 U213 ( .A(\alu_i[SRC_A][8] ), .B(n1684), .C(n1671), .D(
        n1733), .E(n1680), .Z(n134) );
  HS65_LH_OAI212X5 U214 ( .A(\alu_i[SRC_A][14] ), .B(n1684), .C(n119), .D(
        n1735), .E(n1679), .Z(n390) );
  HS65_LH_OAI212X5 U215 ( .A(\alu_i[SRC_A][17] ), .B(n1684), .C(n119), .D(
        n1736), .E(n1681), .Z(n369) );
  HS65_LH_MX41X7 U216 ( .D0(n1723), .S0(n1653), .D1(n1724), .S1(n1767), .D2(
        n1725), .S2(n1659), .D3(n1726), .S3(n1670), .Z(n132) );
  HS65_LH_IVX9 U217 ( .A(n192), .Z(n1754) );
  HS65_LH_IVX9 U218 ( .A(n305), .Z(n1755) );
  HS65_LH_NOR3X4 U219 ( .A(n104), .B(\alu_i[OP][3] ), .C(\alu_i[OP][2] ), .Z(
        n103) );
  HS65_LH_MX41X7 U220 ( .D0(n1725), .S0(n1653), .D1(n1726), .S1(n1650), .D2(
        n1727), .S2(n1658), .D3(\alu_i[SRC_B][29] ), .S3(n1670), .Z(n163) );
  HS65_LH_NOR2X6 U221 ( .A(n421), .B(n220), .Z(n203) );
  HS65_LH_MX41X7 U222 ( .D0(n1711), .S0(n1653), .D1(n1712), .S1(n1650), .D2(
        n1713), .S2(n1659), .D3(n1714), .S3(n1670), .Z(n130) );
  HS65_LH_MX41X7 U223 ( .D0(n1724), .S0(n1652), .D1(n1725), .S1(n1649), .D2(
        n1726), .S2(n1657), .D3(n1727), .S3(n1669), .Z(n110) );
  HS65_LH_MX41X7 U224 ( .D0(\alu_i[SRC_B][22] ), .S0(n1653), .D1(
        \alu_i[SRC_B][23] ), .S1(n1650), .D2(n1723), .S2(n1659), .D3(n1724), 
        .S3(n1670), .Z(n164) );
  HS65_LH_MX41X7 U225 ( .D0(n1719), .S0(n1651), .D1(n1720), .S1(n1647), .D2(
        \alu_i[SRC_B][22] ), .S2(n1656), .D3(\alu_i[SRC_B][23] ), .S3(n1668), 
        .Z(n136) );
  HS65_LH_MX41X7 U226 ( .D0(n1715), .S0(n1653), .D1(n1716), .S1(n1650), .D2(
        n1717), .S2(n1659), .D3(n1718), .S3(n1670), .Z(n128) );
  HS65_LH_MX41X7 U227 ( .D0(n1716), .S0(n1652), .D1(n1717), .S1(n1649), .D2(
        n1718), .S2(n1657), .D3(n1719), .S3(n1669), .Z(n112) );
  HS65_LH_MX41X7 U228 ( .D0(n1704), .S0(n1652), .D1(n1703), .S1(n1648), .D2(
        \alu_i[SRC_B][3] ), .S2(n1657), .D3(\alu_i[SRC_B][2] ), .S3(n1669), 
        .Z(n181) );
  HS65_LH_MX41X7 U229 ( .D0(n1712), .S0(n1652), .D1(n1713), .S1(n1649), .D2(
        n1714), .S2(n1658), .D3(n1715), .S3(n1669), .Z(n114) );
  HS65_LH_MX41X7 U230 ( .D0(n1717), .S0(n1652), .D1(n1716), .S1(n1648), .D2(
        n1715), .S2(n1657), .D3(n1714), .S3(n1669), .Z(n230) );
  HS65_LH_MX41X7 U231 ( .D0(n1718), .S0(n1651), .D1(n1717), .S1(n1648), .D2(
        n1716), .S2(n1656), .D3(n1715), .S3(n1669), .Z(n215) );
  HS65_LH_NOR2X6 U232 ( .A(n192), .B(n193), .Z(n151) );
  HS65_LH_NOR2X6 U233 ( .A(\alu_i[OP][3] ), .B(\alu_i[OP][4] ), .Z(n432) );
  HS65_LH_MX41X7 U234 ( .D0(n1726), .S0(n1652), .D1(n1727), .S1(n1649), .D2(
        \alu_i[SRC_B][29] ), .S2(n1658), .D3(\alu_i[SRC_B][30] ), .S3(n1669), 
        .Z(n141) );
  HS65_LH_MX41X7 U235 ( .D0(n1709), .S0(n1653), .D1(n1647), .S1(n1708), .D2(
        n1707), .S2(n1658), .D3(n1706), .S3(n1670), .Z(n288) );
  HS65_LH_MX41X7 U236 ( .D0(n1710), .S0(n1652), .D1(n1709), .S1(n1649), .D2(
        n1656), .S2(n1708), .D3(n1707), .S3(n1669), .Z(n276) );
  HS65_LH_MX41X7 U237 ( .D0(n1718), .S0(n1653), .D1(n1719), .S1(n1650), .D2(
        n1720), .S2(n1658), .D3(\alu_i[SRC_B][22] ), .S3(n1670), .Z(n153) );
  HS65_LH_IVX9 U238 ( .A(n306), .Z(n1757) );
  HS65_LH_MX41X7 U239 ( .D0(n1715), .S0(n1652), .D1(n1714), .S1(n1648), .D2(
        n1713), .S2(n1657), .D3(n1712), .S3(n1669), .Z(n260) );
  HS65_LH_MX41X7 U240 ( .D0(\alu_i[SRC_B][23] ), .S0(n1652), .D1(n1723), .S1(
        n1650), .D2(n1724), .S2(n1658), .D3(n1725), .S3(n1670), .Z(n155) );
  HS65_LH_MX41X7 U241 ( .D0(n1707), .S0(n1653), .D1(n1647), .S1(n1708), .D2(
        n1709), .S2(n1659), .D3(n1710), .S3(n1670), .Z(n131) );
  HS65_LH_MX41X7 U242 ( .D0(n1711), .S0(n1652), .D1(n1710), .S1(n1649), .D2(
        n1709), .S2(n1658), .D3(n1668), .S3(n1708), .Z(n310) );
  HS65_LH_MX41X7 U243 ( .D0(n1716), .S0(n1651), .D1(n1715), .S1(n1648), .D2(
        n1714), .S2(n1657), .D3(n1713), .S3(n1669), .Z(n249) );
  HS65_LH_MX41X7 U244 ( .D0(n1713), .S0(n1652), .D1(n1712), .S1(n1648), .D2(
        n1711), .S2(n1657), .D3(n1710), .S3(n1669), .Z(n283) );
  HS65_LH_MX41X7 U245 ( .D0(n1714), .S0(n1652), .D1(n1713), .S1(n1648), .D2(
        n1712), .S2(n1657), .D3(n1711), .S3(n1669), .Z(n277) );
  HS65_LH_MX41X7 U246 ( .D0(\alu_i[SRC_B][23] ), .S0(n1651), .D1(
        \alu_i[SRC_B][22] ), .S1(n1647), .D2(n1720), .S2(n1656), .D3(n1719), 
        .S3(n1668), .Z(n213) );
  HS65_LH_IVX9 U247 ( .A(n193), .Z(n1759) );
  HS65_LH_MX41X7 U248 ( .D0(n1719), .S0(n1651), .D1(n1718), .S1(n1648), .D2(
        n1717), .S2(n1657), .D3(n1716), .S3(n1669), .Z(n259) );
  HS65_LH_MX41X7 U249 ( .D0(\alu_i[SRC_B][22] ), .S0(n1651), .D1(n1720), .S1(
        n1647), .D2(n1719), .S2(n1657), .D3(n1718), .S3(n1668), .Z(n229) );
  HS65_LH_IVX9 U250 ( .A(n220), .Z(n1770) );
  HS65_LH_NAND2X7 U251 ( .A(\alu_i[OP][3] ), .B(n1796), .Z(n427) );
  HS65_LH_MX41X7 U252 ( .D0(n1720), .S0(n1651), .D1(n1719), .S1(n1648), .D2(
        n1718), .S2(n1656), .D3(n1717), .S3(n1668), .Z(n248) );
  HS65_LH_MX41X7 U253 ( .D0(n1651), .S0(n1708), .D1(n1707), .S1(n1648), .D2(
        n1706), .S2(n1657), .D3(n1705), .S3(n1669), .Z(n296) );
  HS65_LH_MX41X7 U254 ( .D0(n1704), .S0(n1651), .D1(n1705), .S1(n1648), .D2(
        n1706), .S2(n1657), .D3(n1707), .S3(n1668), .Z(n177) );
  HS65_LH_MX41X7 U255 ( .D0(n1714), .S0(n1653), .D1(n1715), .S1(n1650), .D2(
        n1716), .S2(n1658), .D3(n1717), .S3(n1670), .Z(n154) );
  HS65_LH_MX41X7 U256 ( .D0(n1713), .S0(n1653), .D1(n1714), .S1(n1650), .D2(
        n1715), .S2(n1659), .D3(n1716), .S3(n1670), .Z(n170) );
  HS65_LH_MX41X7 U257 ( .D0(n1717), .S0(n1653), .D1(n1718), .S1(n1650), .D2(
        n1719), .S2(n1658), .D3(n1720), .S3(n1670), .Z(n172) );
  HS65_LH_MX41X7 U258 ( .D0(n1720), .S0(n1652), .D1(\alu_i[SRC_B][22] ), .S1(
        n1648), .D2(\alu_i[SRC_B][23] ), .S2(n1657), .D3(n1723), .S3(n1669), 
        .Z(n123) );
  HS65_LH_MX41X7 U259 ( .D0(n1703), .S0(n1652), .D1(\alu_i[SRC_B][3] ), .S1(
        n1649), .D2(n1656), .S2(\alu_i[SRC_B][2] ), .D3(n1668), .S3(
        \alu_i[SRC_B][1] ), .Z(n309) );
  HS65_LH_MX41X7 U260 ( .D0(n1651), .S0(n1708), .D1(n1709), .S1(n1648), .D2(
        n1710), .S2(n1656), .D3(n1711), .S3(n1668), .Z(n115) );
  HS65_LH_MX41X7 U261 ( .D0(n1712), .S0(n1652), .D1(n1711), .S1(n1649), .D2(
        n1710), .S2(n1657), .D3(n1709), .S3(n1669), .Z(n297) );
  HS65_LH_NAND2X7 U262 ( .A(\alu_i[OP][0] ), .B(n1800), .Z(n102) );
  HS65_LH_MX41X7 U263 ( .D0(n1707), .S0(n1652), .D1(n1706), .S1(n1649), .D2(
        n1705), .S2(n1658), .D3(n1704), .S3(n1669), .Z(n343) );
  HS65_LH_MX41X7 U264 ( .D0(n1709), .S0(n1653), .D1(n1710), .S1(n1650), .D2(
        n1711), .S2(n1658), .D3(n1712), .S3(n1670), .Z(n171) );
  HS65_LH_IVX9 U265 ( .A(\alu_i[OP][1] ), .Z(n1800) );
  HS65_LH_MX41X7 U266 ( .D0(n1710), .S0(n1652), .D1(n1711), .S1(n1649), .D2(
        n1712), .S2(n1658), .D3(n1713), .S3(n1670), .Z(n146) );
  HS65_LH_MX41X7 U267 ( .D0(n1703), .S0(n1653), .D1(n1704), .S1(n1650), .D2(
        n1705), .S2(n1659), .D3(n1706), .S3(n1670), .Z(n194) );
  HS65_LH_MX41X7 U268 ( .D0(n1706), .S0(n1652), .D1(n1707), .S1(n1649), .D2(
        n1656), .S2(n1708), .D3(n1709), .S3(n1669), .Z(n148) );
  HS65_LH_MX41X7 U269 ( .D0(n1705), .S0(n1651), .D1(n1706), .S1(n1647), .D2(
        n1707), .S2(n1656), .D3(n1668), .S3(n1708), .Z(n166) );
  HS65_LH_OAI21X3 U270 ( .A(n1720), .B(n1685), .C(n1680), .Z(n332) );
  HS65_LH_OAI21X3 U271 ( .A(n1723), .B(n1685), .C(n1680), .Z(n302) );
  HS65_LH_OAI21X3 U272 ( .A(n1724), .B(n1685), .C(n1680), .Z(n293) );
  HS65_LH_OAI21X3 U273 ( .A(n1726), .B(n1685), .C(n1680), .Z(n270) );
  HS65_LH_OAI21X3 U274 ( .A(n1709), .B(n1683), .C(n95), .Z(n417) );
  HS65_LH_IVX9 U275 ( .A(\alu_i[OP][4] ), .Z(n1796) );
  HS65_LH_MX41X7 U276 ( .D0(n1726), .S0(n1651), .D1(n1725), .S1(n1647), .D2(
        n1724), .S2(n1656), .D3(n1723), .S3(n1668), .Z(n216) );
  HS65_LH_MX41X7 U277 ( .D0(n1724), .S0(n1651), .D1(n1723), .S1(n1647), .D2(
        \alu_i[SRC_B][23] ), .S2(n1656), .D3(\alu_i[SRC_B][22] ), .S3(n1668), 
        .Z(n250) );
  HS65_LH_MX41X7 U278 ( .D0(n1723), .S0(n1651), .D1(\alu_i[SRC_B][23] ), .S1(
        n1647), .D2(\alu_i[SRC_B][22] ), .S2(n1656), .D3(n1720), .S3(n1668), 
        .Z(n261) );
  HS65_LH_OAI21X3 U279 ( .A(n1731), .B(n1685), .C(n206), .Z(n243) );
  HS65_LH_OAI21X3 U280 ( .A(n1705), .B(n1685), .C(n1679), .Z(n169) );
  HS65_LH_OAI21X3 U281 ( .A(n1707), .B(n1685), .C(n95), .Z(n135) );
  HS65_LH_OAI21X3 U282 ( .A(n1713), .B(n1685), .C(n1679), .Z(n391) );
  HS65_LH_OAI21X3 U283 ( .A(n1714), .B(n1685), .C(n95), .Z(n385) );
  HS65_LH_OAI21X3 U284 ( .A(n1715), .B(n1685), .C(n1679), .Z(n378) );
  HS65_LH_OAI21X3 U285 ( .A(n1716), .B(n1685), .C(n95), .Z(n370) );
  HS65_LH_OAI21X3 U286 ( .A(n1717), .B(n1685), .C(n1679), .Z(n363) );
  HS65_LH_OAI21X3 U287 ( .A(n1718), .B(n1685), .C(n95), .Z(n356) );
  HS65_LH_OAI21X3 U288 ( .A(n1727), .B(n1685), .C(n1680), .Z(n264) );
  HS65_LH_MX41X7 U289 ( .D0(n1725), .S0(n1651), .D1(n1724), .S1(n1647), .D2(
        n1723), .S2(n1656), .D3(\alu_i[SRC_B][23] ), .S3(n1668), .Z(n231) );
  HS65_LH_OAI21X3 U290 ( .A(n1704), .B(n1683), .C(n1679), .Z(n180) );
  HS65_LH_OAI21X3 U291 ( .A(n1706), .B(n92), .C(n95), .Z(n152) );
  HS65_LH_OAI21X3 U292 ( .A(n1708), .B(n1683), .C(n1679), .Z(n118) );
  HS65_LH_NOR3X4 U293 ( .A(n1796), .B(\alu_i[OP][3] ), .C(n435), .Z(
        \alu_o[BRANCH] ) );
  HS65_LH_AOI33X5 U294 ( .A(n104), .B(\alu_i[OP][2] ), .C(N714), .D(n433), .E(
        n1801), .F(N713), .Z(n435) );
  HS65_LH_OAI21X3 U295 ( .A(n1711), .B(n92), .C(n95), .Z(n404) );
  HS65_LH_OAI21X3 U296 ( .A(n1712), .B(n1683), .C(n1679), .Z(n398) );
  HS65_LH_AO33X9 U297 ( .A(n1760), .B(n1758), .C(n1752), .D(n1755), .E(n144), 
        .F(n1759), .Z(n272) );
  HS65_LH_AO222X4 U298 ( .A(n1659), .B(n1725), .C(n1668), .D(n1724), .E(n1647), 
        .F(n1726), .Z(n263) );
  HS65_LH_AO222X4 U299 ( .A(n1659), .B(n1726), .C(n1668), .D(n1725), .E(n1647), 
        .F(n1727), .Z(n252) );
  HS65_LH_AO222X4 U300 ( .A(n1659), .B(n1727), .C(n1668), .D(n1726), .E(n1647), 
        .F(\alu_i[SRC_B][29] ), .Z(n233) );
  HS65_LH_AO312X9 U301 ( .A(n1759), .B(n160), .C(n1755), .D(n1725), .E(n286), 
        .F(n287), .Z(n285) );
  HS65_LH_CBI4I6X5 U302 ( .A(n1725), .B(n1684), .C(n1679), .D(n1739), .Z(n287)
         );
  HS65_LH_OAI212X5 U303 ( .A(\alu_i[SRC_A][26] ), .B(n1683), .C(n1671), .D(
        n1739), .E(n1681), .Z(n286) );
  HS65_LH_BFX9 U304 ( .A(n100), .Z(n1673) );
  HS65_LH_NOR3X4 U305 ( .A(n1797), .B(\alu_i[OP][2] ), .C(n102), .Z(n100) );
  HS65_LH_BFX9 U306 ( .A(n201), .Z(n1667) );
  HS65_LH_NOR2X6 U307 ( .A(n1769), .B(n1771), .Z(n201) );
  HS65_LH_IVX9 U308 ( .A(n357), .Z(n1760) );
  HS65_LH_AO22X9 U309 ( .A(n1705), .B(n211), .C(n288), .D(n214), .Z(n327) );
  HS65_LH_AO22X9 U310 ( .A(n1706), .B(n211), .C(n276), .D(n214), .Z(n319) );
  HS65_LH_BFX9 U311 ( .A(n1741), .Z(n1743) );
  HS65_LH_BFX9 U312 ( .A(n1741), .Z(n1744) );
  HS65_LH_BFX9 U313 ( .A(n1741), .Z(n1745) );
  HS65_LH_BFX9 U314 ( .A(n1742), .Z(n1746) );
  HS65_LH_BFX9 U315 ( .A(n1742), .Z(n1747) );
  HS65_LH_BFX9 U316 ( .A(n1742), .Z(n1748) );
  HS65_LH_AO22X9 U317 ( .A(\HI_LO_c[LO][0] ), .B(n1693), .C(N162), .D(n1689), 
        .Z(n462) );
  HS65_LH_AO22X9 U318 ( .A(\HI_LO_c[HI][1] ), .B(n1696), .C(N195), .D(n1691), 
        .Z(n495) );
  HS65_LH_AO22X9 U319 ( .A(\HI_LO_c[HI][2] ), .B(n1696), .C(N196), .D(n1691), 
        .Z(n496) );
  HS65_LH_AO22X9 U320 ( .A(\HI_LO_c[HI][3] ), .B(n1696), .C(N197), .D(n1691), 
        .Z(n497) );
  HS65_LH_AO22X9 U321 ( .A(\HI_LO_c[HI][5] ), .B(n1696), .C(N199), .D(n1692), 
        .Z(n499) );
  HS65_LH_AO22X9 U322 ( .A(\HI_LO_c[HI][9] ), .B(n1696), .C(N203), .D(n1692), 
        .Z(n503) );
  HS65_LH_AO22X9 U323 ( .A(\HI_LO_c[HI][11] ), .B(n1697), .C(N205), .D(n1692), 
        .Z(n505) );
  HS65_LH_AO22X9 U324 ( .A(\HI_LO_c[HI][13] ), .B(n1697), .C(N207), .D(n1692), 
        .Z(n507) );
  HS65_LH_AO22X9 U325 ( .A(\HI_LO_c[HI][14] ), .B(n1697), .C(N208), .D(n1692), 
        .Z(n508) );
  HS65_LH_AO22X9 U326 ( .A(\HI_LO_c[HI][15] ), .B(n1697), .C(N209), .D(n1692), 
        .Z(n509) );
  HS65_LH_AO22X9 U327 ( .A(\HI_LO_c[HI][16] ), .B(n1697), .C(N210), .D(n1689), 
        .Z(n510) );
  HS65_LH_AO22X9 U328 ( .A(\HI_LO_c[HI][17] ), .B(n1697), .C(N211), .D(n1690), 
        .Z(n511) );
  HS65_LH_AO22X9 U329 ( .A(\HI_LO_c[HI][18] ), .B(n1697), .C(N212), .D(n1691), 
        .Z(n512) );
  HS65_LH_AO22X9 U330 ( .A(\HI_LO_c[HI][19] ), .B(n1697), .C(N213), .D(n1692), 
        .Z(n513) );
  HS65_LH_AO22X9 U331 ( .A(\HI_LO_c[HI][21] ), .B(n1697), .C(N215), .D(n1689), 
        .Z(n515) );
  HS65_LH_AO22X9 U332 ( .A(\HI_LO_c[HI][24] ), .B(n1697), .C(N218), .D(n1690), 
        .Z(n518) );
  HS65_LH_AO22X9 U333 ( .A(\HI_LO_c[HI][25] ), .B(n1697), .C(N219), .D(n1691), 
        .Z(n519) );
  HS65_LH_AO22X9 U334 ( .A(\HI_LO_c[HI][28] ), .B(n1697), .C(N222), .D(n1689), 
        .Z(n522) );
  HS65_LH_AO22X9 U335 ( .A(\HI_LO_c[HI][29] ), .B(n1697), .C(N223), .D(n1690), 
        .Z(n523) );
  HS65_LH_AO22X9 U336 ( .A(\HI_LO_c[HI][30] ), .B(n1698), .C(N224), .D(n1691), 
        .Z(n524) );
  HS65_LH_AO22X9 U337 ( .A(\HI_LO_c[HI][31] ), .B(n1698), .C(N225), .D(n1692), 
        .Z(n525) );
  HS65_LH_AO22X9 U338 ( .A(\HI_LO_c[LO][12] ), .B(n1695), .C(N174), .D(n1690), 
        .Z(n474) );
  HS65_LH_AO22X9 U339 ( .A(\HI_LO_c[LO][16] ), .B(n1695), .C(N178), .D(n1690), 
        .Z(n478) );
  HS65_LH_AO22X9 U340 ( .A(\HI_LO_c[HI][8] ), .B(n1696), .C(N202), .D(n1692), 
        .Z(n502) );
  HS65_LH_AO22X9 U341 ( .A(\HI_LO_c[LO][8] ), .B(n1695), .C(N170), .D(n1689), 
        .Z(n470) );
  HS65_LH_AO22X9 U342 ( .A(\HI_LO_c[LO][13] ), .B(n1695), .C(N175), .D(n1690), 
        .Z(n475) );
  HS65_LH_AO22X9 U343 ( .A(\HI_LO_c[LO][14] ), .B(n1695), .C(N176), .D(n1690), 
        .Z(n476) );
  HS65_LH_AO22X9 U344 ( .A(\HI_LO_c[LO][15] ), .B(n1695), .C(N177), .D(n1690), 
        .Z(n477) );
  HS65_LH_AO22X9 U345 ( .A(\HI_LO_c[HI][6] ), .B(n1696), .C(N200), .D(n1692), 
        .Z(n500) );
  HS65_LH_AO22X9 U346 ( .A(\HI_LO_c[HI][7] ), .B(n1696), .C(N201), .D(n1692), 
        .Z(n501) );
  HS65_LH_AO22X9 U347 ( .A(\HI_LO_c[HI][26] ), .B(n1697), .C(N220), .D(n1692), 
        .Z(n520) );
  HS65_LH_AO22X9 U348 ( .A(\HI_LO_c[LO][20] ), .B(n1695), .C(N182), .D(n1690), 
        .Z(n482) );
  HS65_LH_AO22X9 U349 ( .A(\HI_LO_c[LO][24] ), .B(n1696), .C(N186), .D(n1691), 
        .Z(n486) );
  HS65_LH_AO22X9 U350 ( .A(\HI_LO_c[LO][31] ), .B(n1696), .C(N193), .D(n1691), 
        .Z(n493) );
  HS65_LH_AO22X9 U351 ( .A(\HI_LO_c[LO][4] ), .B(n1695), .C(N166), .D(n1689), 
        .Z(n466) );
  HS65_LH_AO22X9 U352 ( .A(\HI_LO_c[LO][5] ), .B(n1695), .C(N167), .D(n1689), 
        .Z(n467) );
  HS65_LH_AO22X9 U353 ( .A(\HI_LO_c[LO][9] ), .B(n1695), .C(N171), .D(n1689), 
        .Z(n471) );
  HS65_LH_AO22X9 U354 ( .A(\HI_LO_c[LO][11] ), .B(n1695), .C(N173), .D(n1689), 
        .Z(n473) );
  HS65_LH_AO22X9 U355 ( .A(\HI_LO_c[LO][17] ), .B(n1695), .C(N179), .D(n1690), 
        .Z(n479) );
  HS65_LH_AO22X9 U356 ( .A(\HI_LO_c[LO][18] ), .B(n1695), .C(N180), .D(n1690), 
        .Z(n480) );
  HS65_LH_AO22X9 U357 ( .A(\HI_LO_c[LO][19] ), .B(n1695), .C(N181), .D(n1690), 
        .Z(n481) );
  HS65_LH_AO22X9 U358 ( .A(\HI_LO_c[LO][21] ), .B(n1695), .C(N183), .D(n1690), 
        .Z(n483) );
  HS65_LH_AO22X9 U359 ( .A(\HI_LO_c[LO][25] ), .B(n1696), .C(N187), .D(n1691), 
        .Z(n487) );
  HS65_LH_AO22X9 U360 ( .A(\HI_LO_c[LO][29] ), .B(n1696), .C(N191), .D(n1691), 
        .Z(n491) );
  HS65_LH_AO22X9 U361 ( .A(\HI_LO_c[LO][30] ), .B(n1696), .C(N192), .D(n1691), 
        .Z(n492) );
  HS65_LH_AO22X9 U362 ( .A(\HI_LO_c[LO][1] ), .B(n1694), .C(N163), .D(n1689), 
        .Z(n463) );
  HS65_LH_AO22X9 U363 ( .A(\HI_LO_c[LO][2] ), .B(n1695), .C(N164), .D(n1689), 
        .Z(n464) );
  HS65_LH_AO22X9 U364 ( .A(\HI_LO_c[LO][3] ), .B(n1695), .C(N165), .D(n1689), 
        .Z(n465) );
  HS65_LH_AO22X9 U365 ( .A(\HI_LO_c[LO][6] ), .B(n1695), .C(N168), .D(n1689), 
        .Z(n468) );
  HS65_LH_AO22X9 U366 ( .A(\HI_LO_c[LO][7] ), .B(n1695), .C(N169), .D(n1689), 
        .Z(n469) );
  HS65_LH_AO22X9 U367 ( .A(\HI_LO_c[LO][10] ), .B(n1695), .C(N172), .D(n1689), 
        .Z(n472) );
  HS65_LH_AO22X9 U368 ( .A(\HI_LO_c[LO][22] ), .B(n1696), .C(N184), .D(n1690), 
        .Z(n484) );
  HS65_LH_AO22X9 U369 ( .A(\HI_LO_c[LO][23] ), .B(n1696), .C(N185), .D(n1690), 
        .Z(n485) );
  HS65_LH_AO22X9 U370 ( .A(\HI_LO_c[LO][26] ), .B(n1696), .C(N188), .D(n1691), 
        .Z(n488) );
  HS65_LH_AO22X9 U371 ( .A(\HI_LO_c[LO][27] ), .B(n1696), .C(N189), .D(n1691), 
        .Z(n489) );
  HS65_LH_AO22X9 U372 ( .A(\HI_LO_c[HI][0] ), .B(n1696), .C(N194), .D(n1691), 
        .Z(n494) );
  HS65_LH_AO22X9 U373 ( .A(\HI_LO_c[HI][4] ), .B(n1696), .C(N198), .D(n1692), 
        .Z(n498) );
  HS65_LH_AO22X9 U374 ( .A(\HI_LO_c[HI][10] ), .B(n1697), .C(N204), .D(n1692), 
        .Z(n504) );
  HS65_LH_AO22X9 U375 ( .A(\HI_LO_c[HI][20] ), .B(n1697), .C(N214), .D(n1689), 
        .Z(n514) );
  HS65_LH_AO22X9 U376 ( .A(\HI_LO_c[HI][22] ), .B(n1697), .C(N216), .D(n1690), 
        .Z(n516) );
  HS65_LH_AO22X9 U377 ( .A(\HI_LO_c[HI][23] ), .B(n1697), .C(N217), .D(n1691), 
        .Z(n517) );
  HS65_LH_AO22X9 U378 ( .A(\HI_LO_c[HI][27] ), .B(n1697), .C(N221), .D(n1692), 
        .Z(n521) );
  HS65_LH_AO22X9 U379 ( .A(\HI_LO_c[LO][28] ), .B(n1696), .C(N190), .D(n1691), 
        .Z(n490) );
  HS65_LH_AO22X9 U380 ( .A(\HI_LO_c[HI][12] ), .B(n1697), .C(N206), .D(n1692), 
        .Z(n506) );
  HS65_LH_NAND2X7 U381 ( .A(\alu_i[SHAMT][2] ), .B(n1758), .Z(n306) );
  HS65_LH_NAND3X5 U382 ( .A(n97), .B(n433), .C(\alu_i[SHAMT][4] ), .Z(n192) );
  HS65_LH_OAI32X5 U383 ( .A(n189), .B(\alu_i[SHAMT][3] ), .C(n190), .D(n191), 
        .E(n1790), .Z(n188) );
  HS65_LH_OA12X9 U384 ( .A(n92), .B(n1703), .C(n95), .Z(n191) );
  HS65_LH_OAI32X5 U385 ( .A(n357), .B(\alu_i[SHAMT][3] ), .C(n192), .D(n412), 
        .E(n1734), .Z(n411) );
  HS65_LH_OA12X9 U386 ( .A(n1683), .B(n1710), .C(n1679), .Z(n412) );
  HS65_LH_OAI32X5 U387 ( .A(n305), .B(\alu_i[SHAMT][3] ), .C(n189), .D(n341), 
        .E(n1737), .Z(n340) );
  HS65_LH_OA12X9 U388 ( .A(n92), .B(n1719), .C(n95), .Z(n341) );
  HS65_LH_NAND3X5 U389 ( .A(n99), .B(n97), .C(\alu_i[SHAMT][4] ), .Z(n305) );
  HS65_LH_AOI222X2 U390 ( .A(n122), .B(n132), .C(n1665), .D(\HI_LO_c[LO][12] ), 
        .E(n113), .F(n128), .Z(n402) );
  HS65_LH_AOI222X2 U391 ( .A(n1662), .B(\HI_LO_c[HI][31] ), .C(N129), .D(n1677), .E(N161), .F(n1675), .Z(n209) );
  HS65_LH_AOI222X2 U392 ( .A(n1643), .B(n130), .C(n1663), .D(\HI_LO_c[HI][8] ), 
        .E(n1751), .F(n131), .Z(n126) );
  HS65_LH_AOI222X2 U393 ( .A(N114), .B(n1677), .C(n1665), .D(\HI_LO_c[LO][16] ), .E(n1752), .F(n375), .Z(n374) );
  HS65_LH_AOI222X2 U394 ( .A(N113), .B(n1677), .C(n113), .D(n153), .E(n1665), 
        .F(\HI_LO_c[LO][15] ), .Z(n383) );
  HS65_LH_AOI222X2 U395 ( .A(N111), .B(n1677), .C(n109), .D(n121), .E(n1665), 
        .F(\HI_LO_c[LO][13] ), .Z(n395) );
  HS65_LH_AOI222X2 U396 ( .A(n1665), .B(\HI_LO_c[LO][0] ), .C(
        \alu_i[SRC_B][0] ), .D(n430), .E(\alu_i[SRC_B][1] ), .F(n200), .Z(n424) );
  HS65_LH_OAI212X5 U397 ( .A(n396), .B(n421), .C(\alu_i[SRC_A][0] ), .D(n1683), 
        .E(n431), .Z(n430) );
  HS65_LH_OA12X9 U398 ( .A(n1791), .B(n119), .C(n235), .Z(n431) );
  HS65_LH_AOI222X2 U399 ( .A(n1662), .B(\HI_LO_c[HI][1] ), .C(N99), .D(n1677), 
        .E(N131), .F(n1675), .Z(n346) );
  HS65_LH_AOI222X2 U400 ( .A(N112), .B(n1677), .C(n111), .D(n164), .E(n1665), 
        .F(\HI_LO_c[LO][14] ), .Z(n389) );
  HS65_LH_AOI222X2 U401 ( .A(n1663), .B(\HI_LO_c[HI][11] ), .C(N141), .D(n1675), .E(n1660), .F(n1711), .Z(n408) );
  HS65_LH_AOI222X2 U402 ( .A(n1662), .B(\HI_LO_c[HI][21] ), .C(N151), .D(n1674), .E(n1660), .F(\alu_i[SRC_B][22] ), .Z(n330) );
  HS65_LH_AOI222X2 U403 ( .A(n1662), .B(\HI_LO_c[HI][24] ), .C(N154), .D(n1674), .E(n1661), .F(n1724), .Z(n300) );
  HS65_LH_AOI222X2 U404 ( .A(n1662), .B(\HI_LO_c[HI][25] ), .C(N155), .D(n1674), .E(n1661), .F(n1725), .Z(n291) );
  HS65_LH_AOI212X4 U405 ( .A(n273), .B(n160), .C(n1645), .D(n230), .E(n324), 
        .Z(n323) );
  HS65_LH_OAI212X5 U406 ( .A(n325), .B(n1721), .C(n1765), .D(n317), .E(n326), 
        .Z(n324) );
  HS65_LH_IVX9 U407 ( .A(n229), .Z(n1765) );
  HS65_LH_CBI4I1X5 U408 ( .A(n1686), .B(n1721), .C(n1682), .D(
        \alu_i[SRC_A][22] ), .Z(n326) );
  HS65_LH_NAND2X7 U409 ( .A(\alu_i[SHAMT][3] ), .B(n1761), .Z(n193) );
  HS65_LH_OAI22X6 U410 ( .A(\alu_i[SHAMT][2] ), .B(n141), .C(n150), .D(n1761), 
        .Z(n357) );
  HS65_LH_AOI212X4 U411 ( .A(\alu_i[SRC_A][22] ), .B(n1672), .C(n1686), .D(
        n1778), .E(n1682), .Z(n325) );
  HS65_LH_IVX9 U412 ( .A(\alu_i[SRC_A][22] ), .Z(n1778) );
  HS65_LH_NAND2X7 U413 ( .A(\alu_i[SHAMT][0] ), .B(n1769), .Z(n221) );
  HS65_LH_OAI21X3 U414 ( .A(\alu_i[SHAMT][2] ), .B(n309), .C(n405), .Z(n189)
         );
  HS65_LH_OAI21X3 U415 ( .A(n1699), .B(n396), .C(\alu_i[SHAMT][2] ), .Z(n405)
         );
  HS65_LH_OAI212X5 U416 ( .A(\alu_i[SRC_A][21] ), .B(n92), .C(n119), .D(n1779), 
        .E(n1681), .Z(n333) );
  HS65_LH_IVX9 U417 ( .A(\alu_i[SRC_A][21] ), .Z(n1779) );
  HS65_LH_OAI212X5 U418 ( .A(\alu_i[SRC_A][24] ), .B(n1683), .C(n119), .D(
        n1777), .E(n1681), .Z(n303) );
  HS65_LH_IVX9 U419 ( .A(\alu_i[SRC_A][24] ), .Z(n1777) );
  HS65_LH_OAI212X5 U420 ( .A(\alu_i[SRC_A][25] ), .B(n92), .C(n1671), .D(n1776), .E(n1681), .Z(n294) );
  HS65_LH_IVX9 U421 ( .A(\alu_i[SRC_A][25] ), .Z(n1776) );
  HS65_LH_OAI212X5 U422 ( .A(\alu_i[SRC_A][27] ), .B(n1683), .C(n1671), .D(
        n1775), .E(n1681), .Z(n271) );
  HS65_LH_IVX9 U423 ( .A(\alu_i[SRC_A][27] ), .Z(n1775) );
  HS65_LH_OAI212X5 U424 ( .A(\alu_i[SRC_A][4] ), .B(n1684), .C(n1671), .D(
        n1790), .E(n1681), .Z(n187) );
  HS65_LH_OAI212X5 U425 ( .A(\alu_i[SRC_A][10] ), .B(n1684), .C(n119), .D(
        n1786), .E(n1680), .Z(n418) );
  HS65_LH_IVX9 U426 ( .A(\alu_i[SRC_A][10] ), .Z(n1786) );
  HS65_LH_OAI212X5 U427 ( .A(\alu_i[SRC_A][28] ), .B(n92), .C(n1671), .D(n1774), .E(n235), .Z(n262) );
  HS65_LH_IVX9 U428 ( .A(\alu_i[SRC_A][28] ), .Z(n1774) );
  HS65_LH_OAI212X5 U429 ( .A(\alu_i[SRC_A][30] ), .B(n92), .C(n1671), .D(n1773), .E(n235), .Z(n232) );
  HS65_LH_IVX9 U430 ( .A(\alu_i[SRC_A][30] ), .Z(n1773) );
  HS65_LH_OAI212X5 U431 ( .A(\alu_i[SRC_A][31] ), .B(n1683), .C(n1671), .D(
        n1772), .E(n223), .Z(n217) );
  HS65_LH_IVX9 U432 ( .A(\alu_i[SRC_A][31] ), .Z(n1772) );
  HS65_LH_NOR2X6 U433 ( .A(n1682), .B(n1661), .Z(n223) );
  HS65_LH_OAI212X5 U434 ( .A(\alu_i[SRC_A][6] ), .B(n1684), .C(n1671), .D(
        n1789), .E(n1680), .Z(n167) );
  HS65_LH_IVX9 U435 ( .A(\alu_i[SRC_A][6] ), .Z(n1789) );
  HS65_LH_OAI212X5 U436 ( .A(\alu_i[SRC_A][7] ), .B(n1684), .C(n1671), .D(
        n1788), .E(n1680), .Z(n149) );
  HS65_LH_IVX9 U437 ( .A(\alu_i[SRC_A][7] ), .Z(n1788) );
  HS65_LH_OAI212X5 U438 ( .A(\alu_i[SRC_A][16] ), .B(n1684), .C(n119), .D(
        n1782), .E(n1681), .Z(n376) );
  HS65_LH_IVX9 U439 ( .A(\alu_i[SRC_A][16] ), .Z(n1782) );
  HS65_LH_OAI212X5 U440 ( .A(\alu_i[SRC_A][9] ), .B(n1684), .C(n1787), .D(n119), .E(n1681), .Z(n117) );
  HS65_LH_IVX9 U441 ( .A(\alu_i[SRC_A][9] ), .Z(n1787) );
  HS65_LH_OAI212X5 U442 ( .A(\alu_i[SRC_A][12] ), .B(n1684), .C(n119), .D(
        n1785), .E(n95), .Z(n403) );
  HS65_LH_IVX9 U443 ( .A(\alu_i[SRC_A][12] ), .Z(n1785) );
  HS65_LH_OAI212X5 U444 ( .A(\alu_i[SRC_A][13] ), .B(n1684), .C(n1671), .D(
        n1784), .E(n1681), .Z(n397) );
  HS65_LH_IVX9 U445 ( .A(\alu_i[SRC_A][13] ), .Z(n1784) );
  HS65_LH_OAI212X5 U446 ( .A(\alu_i[SRC_A][15] ), .B(n1684), .C(n119), .D(
        n1783), .E(n1681), .Z(n384) );
  HS65_LH_IVX9 U447 ( .A(\alu_i[SRC_A][15] ), .Z(n1783) );
  HS65_LH_OAI212X5 U448 ( .A(\alu_i[SRC_A][18] ), .B(n1684), .C(n1671), .D(
        n1781), .E(n1681), .Z(n362) );
  HS65_LH_IVX9 U449 ( .A(\alu_i[SRC_A][18] ), .Z(n1781) );
  HS65_LH_OAI212X5 U450 ( .A(\alu_i[SRC_A][19] ), .B(n1684), .C(n119), .D(
        n1780), .E(n1681), .Z(n355) );
  HS65_LH_IVX9 U451 ( .A(\alu_i[SRC_A][19] ), .Z(n1780) );
  HS65_LH_NAND2X7 U452 ( .A(\alu_i[SHAMT][1] ), .B(n1771), .Z(n220) );
  HS65_LH_IVX9 U453 ( .A(\alu_i[SHAMT][3] ), .Z(n1758) );
  HS65_LH_IVX9 U454 ( .A(\alu_i[SRC_B][0] ), .Z(n1699) );
  HS65_LH_IVX9 U455 ( .A(\alu_i[SRC_B][31] ), .Z(n1730) );
  HS65_LH_IVX9 U456 ( .A(\alu_i[SRC_B][1] ), .Z(n1700) );
  HS65_LH_IVX9 U457 ( .A(\alu_i[SRC_B][30] ), .Z(n1729) );
  HS65_LH_IVX9 U458 ( .A(\alu_i[SRC_B][22] ), .Z(n1721) );
  HS65_LH_IVX9 U459 ( .A(\alu_i[SRC_B][23] ), .Z(n1722) );
  HS65_LH_IVX9 U460 ( .A(\alu_i[SRC_B][29] ), .Z(n1728) );
  HS65_LH_IVX9 U461 ( .A(\alu_i[SRC_B][2] ), .Z(n1701) );
  HS65_LH_IVX9 U462 ( .A(\alu_i[SRC_B][3] ), .Z(n1702) );
  HS65_LH_AO222X4 U463 ( .A(n155), .B(n1757), .C(\alu_i[SHAMT][3] ), .D(n1760), 
        .E(n153), .F(n1756), .Z(n199) );
  HS65_LH_IVX9 U464 ( .A(\alu_i[SHAMT][2] ), .Z(n1761) );
  HS65_LH_OAI21X3 U465 ( .A(\alu_i[SRC_A][1] ), .B(n1685), .C(n206), .Z(n349)
         );
  HS65_LH_OAI21X3 U466 ( .A(\alu_i[SRC_A][3] ), .B(n92), .C(n206), .Z(n205) );
  HS65_LH_NAND4ABX3 U467 ( .A(n399), .B(n400), .C(n401), .D(n402), .Z(
        \alu_o[RESULT][12] ) );
  HS65_LH_MX41X7 U468 ( .D0(n109), .S0(n129), .D1(n1750), .S1(n265), .D2(n1711), .S2(n403), .D3(\alu_i[SRC_A][12] ), .S3(n404), .Z(n400) );
  HS65_LH_AO222X4 U469 ( .A(\HI_LO_c[HI][12] ), .B(n1664), .C(n1712), .D(n1661), .E(n130), .F(n1751), .Z(n399) );
  HS65_LH_AOI222X2 U470 ( .A(N142), .B(n1674), .C(n111), .D(n136), .E(N110), 
        .F(n1677), .Z(n401) );
  HS65_LH_NAND4ABX3 U471 ( .A(n105), .B(n106), .C(n107), .D(n108), .Z(
        \alu_o[RESULT][9] ) );
  HS65_LH_MX41X7 U472 ( .D0(n1751), .S0(n115), .D1(n1750), .S1(n116), .D2(
        n1708), .S2(n117), .D3(\alu_i[SRC_A][9] ), .S3(n118), .Z(n106) );
  HS65_LH_MX41X7 U473 ( .D0(N107), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][9] ), .D2(n120), .S2(n121), .D3(n122), .S3(n123), .Z(n105) );
  HS65_LH_AOI222X2 U474 ( .A(n1662), .B(\HI_LO_c[HI][9] ), .C(N139), .D(n1674), 
        .E(n1660), .F(n1709), .Z(n107) );
  HS65_LH_NAND4ABX3 U475 ( .A(n365), .B(n366), .C(n367), .D(n368), .Z(
        \alu_o[RESULT][17] ) );
  HS65_LH_MX41X7 U476 ( .D0(n1749), .S0(n249), .D1(n1752), .S1(n350), .D2(
        n1716), .S2(n369), .D3(\alu_i[SRC_A][17] ), .S3(n370), .Z(n366) );
  HS65_LH_MX41X7 U477 ( .D0(N115), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][17] ), .D2(n1645), .S2(n297), .D3(n212), .S3(n296), .Z(
        n365) );
  HS65_LH_AOI222X2 U478 ( .A(n1663), .B(\HI_LO_c[HI][17] ), .C(N147), .D(n1674), .E(n1660), .F(n1717), .Z(n367) );
  HS65_LH_NAND4ABX3 U479 ( .A(n358), .B(n359), .C(n360), .D(n361), .Z(
        \alu_o[RESULT][18] ) );
  HS65_LH_MX41X7 U480 ( .D0(n1749), .S0(n230), .D1(n1752), .S1(n241), .D2(
        n1717), .S2(n362), .D3(\alu_i[SRC_A][18] ), .S3(n363), .Z(n359) );
  HS65_LH_MX41X7 U481 ( .D0(N116), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][18] ), .D2(n212), .S2(n288), .D3(n1646), .S3(n283), .Z(
        n358) );
  HS65_LH_AOI222X2 U482 ( .A(n1663), .B(\HI_LO_c[HI][18] ), .C(N148), .D(n1674), .E(n1660), .F(n1718), .Z(n360) );
  HS65_LH_NAND4ABX3 U483 ( .A(n351), .B(n352), .C(n353), .D(n354), .Z(
        \alu_o[RESULT][19] ) );
  HS65_LH_MX41X7 U484 ( .D0(n1749), .S0(n215), .D1(n1752), .S1(n199), .D2(
        n1718), .S2(n355), .D3(\alu_i[SRC_A][19] ), .S3(n356), .Z(n352) );
  HS65_LH_MX41X7 U485 ( .D0(N117), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][19] ), .D2(n212), .S2(n276), .D3(n145), .S3(n277), .Z(
        n351) );
  HS65_LH_AOI222X2 U486 ( .A(n1663), .B(\HI_LO_c[HI][19] ), .C(N149), .D(n1674), .E(n1660), .F(n1719), .Z(n353) );
  HS65_LH_NAND4ABX3 U487 ( .A(n371), .B(n372), .C(n373), .D(n374), .Z(
        \alu_o[RESULT][16] ) );
  HS65_LH_MX41X7 U488 ( .D0(n1749), .S0(n260), .D1(n1715), .S1(n376), .D2(
        \alu_i[SRC_B][0] ), .S2(n377), .D3(\alu_i[SRC_A][16] ), .S3(n378), .Z(
        n371) );
  HS65_LH_AO222X4 U489 ( .A(n343), .B(n212), .C(n309), .D(n214), .E(n310), .F(
        n1646), .Z(n372) );
  HS65_LH_AOI222X2 U490 ( .A(n1663), .B(\HI_LO_c[HI][16] ), .C(N146), .D(n1675), .E(n1660), .F(n1716), .Z(n373) );
  HS65_LH_NAND4ABX3 U491 ( .A(n255), .B(n256), .C(n257), .D(n258), .Z(
        \alu_o[RESULT][28] ) );
  HS65_LH_MX41X7 U492 ( .D0(n1645), .S0(n261), .D1(n1727), .S1(n262), .D2(
        n1749), .S2(n263), .D3(\alu_i[SRC_A][28] ), .S3(n264), .Z(n256) );
  HS65_LH_MX41X7 U493 ( .D0(N126), .S0(n1678), .D1(n1751), .S1(n129), .D2(
        n1665), .S2(\HI_LO_c[LO][28] ), .D3(n1755), .S3(n265), .Z(n255) );
  HS65_LH_AOI222X2 U494 ( .A(n1662), .B(\HI_LO_c[HI][28] ), .C(N158), .D(n1674), .E(n1661), .F(\alu_i[SRC_B][29] ), .Z(n257) );
  HS65_LH_NAND4ABX3 U495 ( .A(n244), .B(n245), .C(n246), .D(n247), .Z(
        \alu_o[RESULT][29] ) );
  HS65_LH_MX41X7 U496 ( .D0(n1646), .S0(n250), .D1(\alu_i[SRC_B][29] ), .S1(
        n251), .D2(n1749), .S2(n252), .D3(\alu_i[SRC_A][29] ), .S3(n253), .Z(
        n245) );
  HS65_LH_MX41X7 U497 ( .D0(N127), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][29] ), .D2(n1751), .S2(n121), .D3(n1755), .S3(n254), .Z(
        n244) );
  HS65_LH_AOI222X2 U498 ( .A(n1662), .B(\HI_LO_c[HI][29] ), .C(N159), .D(n1674), .E(n1660), .F(\alu_i[SRC_B][30] ), .Z(n246) );
  HS65_LH_NAND4ABX3 U499 ( .A(n225), .B(n226), .C(n227), .D(n228), .Z(
        \alu_o[RESULT][30] ) );
  HS65_LH_MX41X7 U500 ( .D0(n145), .S0(n231), .D1(\alu_i[SRC_B][30] ), .S1(
        n232), .D2(n1749), .S2(n233), .D3(\alu_i[SRC_A][30] ), .S3(n234), .Z(
        n226) );
  HS65_LH_MX41X7 U501 ( .D0(N128), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][30] ), .D2(n1751), .S2(n168), .D3(n1755), .S3(n236), .Z(
        n225) );
  HS65_LH_AOI222X2 U502 ( .A(n1662), .B(\HI_LO_c[HI][30] ), .C(N160), .D(n1674), .E(n1660), .F(\alu_i[SRC_B][31] ), .Z(n227) );
  HS65_LH_NAND4ABX3 U503 ( .A(n207), .B(n208), .C(n209), .D(n210), .Z(
        \alu_o[RESULT][31] ) );
  HS65_LH_MX41X7 U504 ( .D0(n1645), .S0(n216), .D1(\alu_i[SRC_B][31] ), .S1(
        n217), .D2(n1749), .S2(n218), .D3(\alu_i[SRC_A][31] ), .S3(n219), .Z(
        n208) );
  HS65_LH_AO222X4 U505 ( .A(n1641), .B(n150), .C(n224), .D(n1755), .E(
        \HI_LO_c[LO][31] ), .F(n1666), .Z(n207) );
  HS65_LH_AOI222X2 U506 ( .A(n211), .B(n1714), .C(n212), .D(n213), .E(n214), 
        .F(n215), .Z(n210) );
  HS65_LH_NAND4ABX3 U507 ( .A(n237), .B(n238), .C(n239), .D(n240), .Z(
        \alu_o[RESULT][2] ) );
  HS65_LH_MX41X7 U508 ( .D0(n1731), .S0(n242), .D1(n203), .S1(n1703), .D2(n204), .S2(n1704), .D3(\alu_i[SRC_B][2] ), .S3(n243), .Z(n238) );
  HS65_LH_MX41X7 U509 ( .D0(n1666), .S0(\HI_LO_c[LO][2] ), .D1(n122), .S1(n170), .D2(n111), .S2(n171), .D3(n1749), .S3(n160), .Z(n237) );
  HS65_LH_AOI222X2 U510 ( .A(n1662), .B(\HI_LO_c[HI][2] ), .C(N100), .D(n1677), 
        .E(N132), .F(n1675), .Z(n239) );
  HS65_LH_NAND4ABX3 U511 ( .A(n380), .B(n381), .C(n382), .D(n383), .Z(
        \alu_o[RESULT][15] ) );
  HS65_LH_MX41X7 U512 ( .D0(n150), .S0(n109), .D1(n1750), .S1(n224), .D2(n1714), .S2(n384), .D3(\alu_i[SRC_A][15] ), .S3(n385), .Z(n380) );
  HS65_LH_AO222X4 U513 ( .A(n155), .B(n111), .C(n141), .D(n122), .E(n154), .F(
        n1751), .Z(n381) );
  HS65_LH_AOI222X2 U514 ( .A(n1663), .B(\HI_LO_c[HI][15] ), .C(N145), .D(n1674), .E(n1660), .F(n1715), .Z(n382) );
  HS65_LH_NAND4ABX3 U515 ( .A(n195), .B(n196), .C(n197), .D(n198), .Z(
        \alu_o[RESULT][3] ) );
  HS65_LH_MX41X7 U516 ( .D0(\alu_i[SRC_A][3] ), .S0(n202), .D1(n203), .S1(
        n1704), .D2(n204), .S2(n1705), .D3(\alu_i[SRC_B][3] ), .S3(n205), .Z(
        n196) );
  HS65_LH_MX41X7 U517 ( .D0(n1666), .S0(\HI_LO_c[LO][3] ), .D1(n122), .S1(n154), .D2(n1749), .S2(n144), .D3(n111), .S3(n146), .Z(n195) );
  HS65_LH_AOI222X2 U518 ( .A(n1662), .B(\HI_LO_c[HI][3] ), .C(N101), .D(n1677), 
        .E(N133), .F(n1675), .Z(n197) );
  HS65_LH_NAND4ABX3 U519 ( .A(n124), .B(n125), .C(n126), .D(n127), .Z(
        \alu_o[RESULT][8] ) );
  HS65_LH_MX41X7 U520 ( .D0(n109), .S0(n132), .D1(n1750), .S1(n133), .D2(n1707), .S2(n134), .D3(\alu_i[SRC_A][8] ), .S3(n135), .Z(n125) );
  HS65_LH_MX41X7 U521 ( .D0(n1661), .S0(n1708), .D1(N138), .S1(n1675), .D2(
        N106), .S2(n1678), .D3(n122), .S3(n136), .Z(n124) );
  HS65_LH_AOI222X2 U522 ( .A(n111), .B(n128), .C(n120), .D(n129), .E(n1665), 
        .F(\HI_LO_c[LO][8] ), .Z(n127) );
  HS65_LH_NAND4ABX3 U523 ( .A(n173), .B(n174), .C(n175), .D(n176), .Z(
        \alu_o[RESULT][5] ) );
  HS65_LH_MX41X7 U524 ( .D0(n1643), .S0(n115), .D1(n1754), .S1(n178), .D2(
        n1704), .S2(n179), .D3(\alu_i[SRC_A][5] ), .S3(n180), .Z(n174) );
  HS65_LH_MX41X7 U525 ( .D0(N103), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][5] ), .D2(n1749), .S2(n181), .D3(n145), .S3(n182), .Z(
        n173) );
  HS65_LH_AOI222X2 U526 ( .A(n1662), .B(\HI_LO_c[HI][5] ), .C(N135), .D(n1674), 
        .E(n1660), .F(n1705), .Z(n175) );
  HS65_LH_NAND4ABX3 U527 ( .A(n392), .B(n393), .C(n394), .D(n395), .Z(
        \alu_o[RESULT][13] ) );
  HS65_LH_MX41X7 U528 ( .D0(n1751), .S0(n114), .D1(n1643), .S1(n112), .D2(
        n1712), .S2(n397), .D3(\alu_i[SRC_A][13] ), .S3(n398), .Z(n392) );
  HS65_LH_AO222X4 U529 ( .A(n110), .B(n122), .C(n254), .D(n1750), .E(n123), 
        .F(n111), .Z(n393) );
  HS65_LH_AOI222X2 U530 ( .A(n1663), .B(\HI_LO_c[HI][13] ), .C(N143), .D(n1675), .E(n1660), .F(n1713), .Z(n394) );
  HS65_LH_NAND4ABX3 U531 ( .A(n344), .B(n345), .C(n346), .D(n347), .Z(
        \alu_o[RESULT][1] ) );
  HS65_LH_MX41X7 U532 ( .D0(\alu_i[SRC_A][1] ), .S0(n348), .D1(n203), .S1(
        \alu_i[SRC_B][3] ), .D2(n204), .S2(n1703), .D3(\alu_i[SRC_B][1] ), 
        .S3(n349), .Z(n345) );
  HS65_LH_MX41X7 U533 ( .D0(n1666), .S0(\HI_LO_c[LO][1] ), .D1(n1749), .S1(
        n182), .D2(n122), .S2(n114), .D3(n1754), .S3(n350), .Z(n344) );
  HS65_LH_AOI222X2 U534 ( .A(n113), .B(n177), .C(n111), .D(n115), .E(
        \alu_i[SRC_B][2] ), .F(n200), .Z(n347) );
  HS65_LH_NAND4ABX3 U535 ( .A(n386), .B(n387), .C(n388), .D(n389), .Z(
        \alu_o[RESULT][14] ) );
  HS65_LH_MX41X7 U536 ( .D0(n109), .S0(n168), .D1(n1750), .S1(n236), .D2(n1713), .S2(n390), .D3(\alu_i[SRC_A][14] ), .S3(n391), .Z(n386) );
  HS65_LH_AO222X4 U537 ( .A(n172), .B(n1644), .C(n163), .D(n122), .E(n170), 
        .F(n1641), .Z(n387) );
  HS65_LH_AOI222X2 U538 ( .A(n1663), .B(\HI_LO_c[HI][14] ), .C(N144), .D(n1675), .E(n1660), .F(n1714), .Z(n388) );
  HS65_LH_NAND4ABX3 U539 ( .A(n406), .B(n407), .C(n408), .D(n409), .Z(
        \alu_o[RESULT][11] ) );
  HS65_LH_MX41X7 U540 ( .D0(n122), .S0(n155), .D1(n212), .S1(n144), .D2(n1751), 
        .S2(n146), .D3(n1749), .S3(n276), .Z(n407) );
  HS65_LH_MX41X7 U541 ( .D0(N109), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][11] ), .D2(n111), .S2(n153), .D3(n1644), .S3(n154), .Z(
        n406) );
  HS65_LH_AOI212X4 U542 ( .A(n1710), .B(n410), .C(n145), .D(n142), .E(n411), 
        .Z(n409) );
  HS65_LH_NAND4ABX3 U543 ( .A(n311), .B(n312), .C(n313), .D(n314), .Z(
        \alu_o[RESULT][23] ) );
  HS65_LH_MX41X7 U544 ( .D0(n1663), .S0(\HI_LO_c[HI][23] ), .D1(n1661), .S1(
        n1723), .D2(N153), .S2(n1675), .D3(N121), .S3(n1678), .Z(n312) );
  HS65_LH_MX41X7 U545 ( .D0(n1666), .S0(\HI_LO_c[LO][23] ), .D1(n1751), .S1(
        n155), .D2(n1644), .S2(n141), .D3(n150), .S3(n111), .Z(n311) );
  HS65_LH_AOI212X4 U546 ( .A(n275), .B(n142), .C(n212), .D(n277), .E(n319), 
        .Z(n313) );
  HS65_LH_NAND4ABX3 U547 ( .A(n320), .B(n321), .C(n322), .D(n323), .Z(
        \alu_o[RESULT][22] ) );
  HS65_LH_MX41X7 U548 ( .D0(n1663), .S0(\HI_LO_c[HI][22] ), .D1(n1661), .S1(
        \alu_i[SRC_B][23] ), .D2(N152), .S2(n1675), .D3(N120), .S3(n1678), .Z(
        n321) );
  HS65_LH_MX41X7 U549 ( .D0(n1666), .S0(\HI_LO_c[LO][22] ), .D1(n1751), .S1(
        n164), .D2(n111), .S2(n168), .D3(n113), .S3(n163), .Z(n320) );
  HS65_LH_AOI212X4 U550 ( .A(n275), .B(n161), .C(n212), .D(n283), .E(n327), 
        .Z(n322) );
  HS65_LH_NAND4ABX3 U551 ( .A(n278), .B(n279), .C(n280), .D(n281), .Z(
        \alu_o[RESULT][26] ) );
  HS65_LH_AO212X4 U552 ( .A(n231), .B(n1642), .C(n229), .D(n1645), .E(n285), 
        .Z(n279) );
  HS65_LH_MX41X7 U553 ( .D0(n1666), .S0(\HI_LO_c[LO][26] ), .D1(n113), .S1(
        n168), .D2(n1751), .S2(n163), .D3(n275), .S3(n288), .Z(n278) );
  HS65_LH_AOI212X4 U554 ( .A(N124), .B(n1677), .C(N156), .D(n1675), .E(n284), 
        .Z(n280) );
  HS65_LH_NAND4ABX3 U555 ( .A(n156), .B(n157), .C(n158), .D(n159), .Z(
        \alu_o[RESULT][6] ) );
  HS65_LH_MX41X7 U556 ( .D0(n1751), .S0(n166), .D1(n1705), .S1(n167), .D2(n151), .S2(n168), .D3(\alu_i[SRC_A][6] ), .S3(n169), .Z(n157) );
  HS65_LH_MX41X7 U557 ( .D0(n1666), .S0(\HI_LO_c[LO][6] ), .D1(n111), .S1(n170), .D2(n1644), .S2(n171), .D3(n122), .S3(n172), .Z(n156) );
  HS65_LH_AOI212X4 U558 ( .A(N104), .B(n1677), .C(N136), .D(n1675), .E(n165), 
        .Z(n158) );
  HS65_LH_NAND4ABX3 U559 ( .A(n137), .B(n138), .C(n139), .D(n140), .Z(
        \alu_o[RESULT][7] ) );
  HS65_LH_MX41X7 U560 ( .D0(n1751), .S0(n148), .D1(n1706), .S1(n149), .D2(n150), .S2(n151), .D3(\alu_i[SRC_A][7] ), .S3(n152), .Z(n138) );
  HS65_LH_MX41X7 U561 ( .D0(n1666), .S0(\HI_LO_c[LO][7] ), .D1(n122), .S1(n153), .D2(n111), .S2(n154), .D3(n109), .S3(n155), .Z(n137) );
  HS65_LH_AOI212X4 U562 ( .A(N105), .B(n1677), .C(N137), .D(n1675), .E(n147), 
        .Z(n139) );
  HS65_LH_NAND4ABX3 U563 ( .A(n335), .B(n336), .C(n337), .D(n338), .Z(
        \alu_o[RESULT][20] ) );
  HS65_LH_MX41X7 U564 ( .D0(n1663), .S0(\HI_LO_c[HI][20] ), .D1(n1661), .S1(
        n1720), .D2(N150), .S2(n1676), .D3(N118), .S3(n1678), .Z(n336) );
  HS65_LH_MX41X7 U565 ( .D0(n1751), .S0(n136), .D1(n1644), .S1(n132), .D2(n111), .S2(n129), .D3(n1666), .S3(\HI_LO_c[LO][20] ), .Z(n335) );
  HS65_LH_AOI212X4 U566 ( .A(n1719), .B(n339), .C(n1749), .D(n259), .E(n340), 
        .Z(n338) );
  HS65_LH_NAND4ABX3 U567 ( .A(n422), .B(n423), .C(n424), .D(n425), .Z(
        \alu_o[RESULT][0] ) );
  HS65_LH_MX41X7 U568 ( .D0(n1663), .S0(\HI_LO_c[HI][0] ), .D1(N130), .S1(
        n1675), .D2(N98), .S2(n1678), .D3(n1754), .S3(n375), .Z(n422) );
  HS65_LH_AO222X4 U569 ( .A(n194), .B(n1644), .C(n131), .D(n111), .E(n130), 
        .F(n122), .Z(n423) );
  HS65_LH_AOI212X4 U570 ( .A(n204), .B(\alu_i[SRC_B][3] ), .C(n203), .D(
        \alu_i[SRC_B][2] ), .E(n426), .Z(n425) );
  HS65_LH_NAND4ABX3 U571 ( .A(n266), .B(n267), .C(n268), .D(n269), .Z(
        \alu_o[RESULT][27] ) );
  HS65_LH_MX41X7 U572 ( .D0(n1663), .S0(\HI_LO_c[HI][27] ), .D1(n1661), .S1(
        n1727), .D2(N157), .S2(n1675), .D3(N125), .S3(n1678), .Z(n267) );
  HS65_LH_MX41X7 U573 ( .D0(n1666), .S0(\HI_LO_c[LO][27] ), .D1(n275), .S1(
        n276), .D2(n211), .S2(n1710), .D3(n214), .S3(n277), .Z(n266) );
  HS65_LH_AOI212X4 U574 ( .A(\alu_i[SRC_A][27] ), .B(n270), .C(n1726), .D(n271), .E(n272), .Z(n269) );
  HS65_LH_NAND4ABX3 U575 ( .A(n289), .B(n290), .C(n291), .D(n292), .Z(
        \alu_o[RESULT][25] ) );
  HS65_LH_MX41X7 U576 ( .D0(N123), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][25] ), .D2(n1643), .S2(n121), .D3(n1751), .S3(n110), .Z(
        n289) );
  HS65_LH_MX41X7 U577 ( .D0(n211), .S0(n1708), .D1(n214), .S1(n297), .D2(n212), 
        .S2(n249), .D3(n1646), .S3(n248), .Z(n290) );
  HS65_LH_AOI212X4 U578 ( .A(\alu_i[SRC_A][25] ), .B(n293), .C(n1724), .D(n294), .E(n295), .Z(n292) );
  HS65_LH_NAND4ABX3 U579 ( .A(n183), .B(n184), .C(n185), .D(n186), .Z(
        \alu_o[RESULT][4] ) );
  HS65_LH_MX41X7 U580 ( .D0(n1663), .S0(\HI_LO_c[HI][4] ), .D1(n1661), .S1(
        n1704), .D2(N134), .S2(n1676), .D3(N102), .S3(n1678), .Z(n183) );
  HS65_LH_MX41X7 U581 ( .D0(n122), .S0(n128), .D1(n1665), .S1(\HI_LO_c[LO][4] ), .D2(n120), .S2(n132), .D3(n109), .S3(n136), .Z(n184) );
  HS65_LH_AOI212X4 U582 ( .A(n151), .B(n129), .C(n1703), .D(n187), .E(n188), 
        .Z(n186) );
  HS65_LH_NAND4ABX3 U583 ( .A(n298), .B(n299), .C(n300), .D(n301), .Z(
        \alu_o[RESULT][24] ) );
  HS65_LH_MX41X7 U584 ( .D0(N122), .S0(n1678), .D1(n1751), .S1(n132), .D2(n113), .S2(n129), .D3(n1666), .S3(\HI_LO_c[LO][24] ), .Z(n298) );
  HS65_LH_MX41X7 U585 ( .D0(n211), .S0(n1707), .D1(n214), .S1(n310), .D2(n212), 
        .S2(n260), .D3(n1645), .S3(n259), .Z(n299) );
  HS65_LH_AOI212X4 U586 ( .A(\alu_i[SRC_A][24] ), .B(n302), .C(n1723), .D(n303), .E(n304), .Z(n301) );
  HS65_LH_NAND4ABX3 U587 ( .A(n328), .B(n329), .C(n330), .D(n331), .Z(
        \alu_o[RESULT][21] ) );
  HS65_LH_MX41X7 U588 ( .D0(n211), .S0(n1704), .D1(n214), .S1(n296), .D2(n1646), .S2(n249), .D3(n273), .S3(n182), .Z(n329) );
  HS65_LH_MX41X7 U589 ( .D0(N119), .S0(n1678), .D1(n1665), .S1(
        \HI_LO_c[LO][21] ), .D2(n212), .S2(n297), .D3(n275), .S3(n181), .Z(
        n328) );
  HS65_LH_AOI212X4 U590 ( .A(\alu_i[SRC_A][21] ), .B(n332), .C(n1720), .D(n333), .E(n334), .Z(n331) );
  HS65_LH_NAND4ABX3 U591 ( .A(n413), .B(n414), .C(n415), .D(n416), .Z(
        \alu_o[RESULT][10] ) );
  HS65_LH_MX41X7 U592 ( .D0(n1663), .S0(\HI_LO_c[HI][10] ), .D1(n1661), .S1(
        n1710), .D2(N140), .S2(n1676), .D3(N108), .S3(n1677), .Z(n414) );
  HS65_LH_MX41X7 U593 ( .D0(n1666), .S0(\HI_LO_c[LO][10] ), .D1(n122), .S1(
        n164), .D2(n1643), .S2(n170), .D3(n1642), .S3(n288), .Z(n413) );
  HS65_LH_AOI212X4 U594 ( .A(\alu_i[SRC_A][10] ), .B(n417), .C(n1709), .D(n418), .E(n419), .Z(n416) );
  HS65_LH_IVX9 U595 ( .A(\alu_i[SHAMT][1] ), .Z(n1769) );
  HS65_LH_IVX9 U596 ( .A(\alu_i[SHAMT][0] ), .Z(n1771) );
  HS65_LH_IVX9 U597 ( .A(\alu_i[SRC_A][26] ), .Z(n1739) );
  HS65_LH_IVX9 U598 ( .A(\alu_i[SRC_A][11] ), .Z(n1734) );
  HS65_LH_IVX9 U599 ( .A(\alu_i[SRC_A][20] ), .Z(n1737) );
  HS65_LH_IVX9 U600 ( .A(\alu_i[SRC_A][5] ), .Z(n1732) );
  HS65_LH_IVX9 U601 ( .A(\alu_i[SRC_A][8] ), .Z(n1733) );
  HS65_LH_IVX9 U602 ( .A(\alu_i[SRC_A][14] ), .Z(n1735) );
  HS65_LH_IVX9 U603 ( .A(\alu_i[SRC_A][17] ), .Z(n1736) );
  HS65_LH_IVX9 U604 ( .A(\alu_i[SRC_A][29] ), .Z(n1740) );
  HS65_LH_IVX9 U605 ( .A(\alu_i[SRC_A][23] ), .Z(n1738) );
  HS65_LH_BFX9 U606 ( .A(rst_n), .Z(n1741) );
  HS65_LH_BFX9 U607 ( .A(rst_n), .Z(n1742) );
  HS65_LH_BFX9 U608 ( .A(\alu_i[SRC_A][2] ), .Z(n1731) );
  HS65_LH_AO22X9 U609 ( .A(\HI_LO_c[HI][26] ), .B(n1664), .C(n1726), .D(n1661), 
        .Z(n284) );
  HS65_LH_AO22X9 U610 ( .A(\HI_LO_c[HI][6] ), .B(n1664), .C(n1706), .D(n1661), 
        .Z(n165) );
  HS65_LH_AO22X9 U611 ( .A(\HI_LO_c[HI][7] ), .B(n1664), .C(n1707), .D(n1661), 
        .Z(n147) );
  HS65_LH_IVX9 U612 ( .A(\alu_i[SHAMT][4] ), .Z(n1753) );
  HS65_LH_IVX9 U613 ( .A(\alu_i[SRC_A][4] ), .Z(n1790) );
  HS65_LH_IVX9 U614 ( .A(\alu_i[SRC_A][0] ), .Z(n1791) );
endmodule


module alu_ctrl ( .alu_ctrl_i({\alu_ctrl_i[OP][3] , \alu_ctrl_i[OP][2] , 
        \alu_ctrl_i[OP][1] , \alu_ctrl_i[OP][0] , \alu_ctrl_i[FUNCT][5] , 
        \alu_ctrl_i[FUNCT][4] , \alu_ctrl_i[FUNCT][3] , \alu_ctrl_i[FUNCT][2] , 
        \alu_ctrl_i[FUNCT][1] , \alu_ctrl_i[FUNCT][0] }), .alu_ctrl_o({
        \alu_ctrl_o[OP][4] , \alu_ctrl_o[OP][3] , \alu_ctrl_o[OP][2] , 
        \alu_ctrl_o[OP][1] , \alu_ctrl_o[OP][0] }) );
  input \alu_ctrl_i[OP][3] , \alu_ctrl_i[OP][2] , \alu_ctrl_i[OP][1] ,
         \alu_ctrl_i[OP][0] , \alu_ctrl_i[FUNCT][5] , \alu_ctrl_i[FUNCT][4] ,
         \alu_ctrl_i[FUNCT][3] , \alu_ctrl_i[FUNCT][2] ,
         \alu_ctrl_i[FUNCT][1] , \alu_ctrl_i[FUNCT][0] ;
  output \alu_ctrl_o[OP][4] , \alu_ctrl_o[OP][3] , \alu_ctrl_o[OP][2] ,
         \alu_ctrl_o[OP][1] , \alu_ctrl_o[OP][0] ;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125;

  HS65_LH_NOR2X6 U3 ( .A(n33), .B(n116), .Z(n22) );
  HS65_LH_NOR2X6 U4 ( .A(n124), .B(n125), .Z(n19) );
  HS65_LH_AOI12X2 U5 ( .A(n124), .B(n125), .C(n19), .Z(n13) );
  HS65_LH_NAND2X7 U6 ( .A(n26), .B(n22), .Z(n16) );
  HS65_LH_NAND2X7 U7 ( .A(n118), .B(n119), .Z(n33) );
  HS65_LH_NOR2X6 U8 ( .A(n25), .B(n123), .Z(n23) );
  HS65_LH_IVX9 U9 ( .A(n24), .Z(n116) );
  HS65_LH_OAI212X5 U10 ( .A(n16), .B(n20), .C(n12), .D(n118), .E(n21), .Z(
        \alu_ctrl_o[OP][2] ) );
  HS65_LH_OAI21X3 U11 ( .A(\alu_ctrl_i[FUNCT][1] ), .B(n121), .C(n125), .Z(n20) );
  HS65_LH_AOI13X5 U12 ( .A(n13), .B(n22), .C(n23), .D(n117), .Z(n21) );
  HS65_LH_IVX9 U13 ( .A(n18), .Z(n117) );
  HS65_LH_OAI212X5 U14 ( .A(\alu_ctrl_i[OP][3] ), .B(n27), .C(
        \alu_ctrl_i[FUNCT][0] ), .D(n17), .E(n31), .Z(\alu_ctrl_o[OP][0] ) );
  HS65_LH_AOI32X5 U15 ( .A(n22), .B(n32), .C(n120), .D(n24), .E(n33), .Z(n31)
         );
  HS65_LH_IVX9 U16 ( .A(n25), .Z(n120) );
  HS65_LH_AO22X9 U17 ( .A(n125), .B(\alu_ctrl_i[FUNCT][2] ), .C(n123), .D(n19), 
        .Z(n32) );
  HS65_LH_OAI211X5 U18 ( .A(n15), .B(n16), .C(n17), .D(n18), .Z(
        \alu_ctrl_o[OP][3] ) );
  HS65_LH_AOI22X6 U19 ( .A(n19), .B(n121), .C(\alu_ctrl_i[FUNCT][4] ), .D(n125), .Z(n15) );
  HS65_LH_OAI212X5 U20 ( .A(\alu_ctrl_i[OP][3] ), .B(n27), .C(n125), .D(n17), 
        .E(n28), .Z(\alu_ctrl_o[OP][1] ) );
  HS65_LH_AOI33X5 U21 ( .A(n29), .B(n124), .C(n22), .D(\alu_ctrl_i[OP][1] ), 
        .E(n24), .F(\alu_ctrl_i[OP][2] ), .Z(n28) );
  HS65_LH_OAI33X3 U22 ( .A(n30), .B(\alu_ctrl_i[FUNCT][5] ), .C(
        \alu_ctrl_i[FUNCT][2] ), .D(n123), .E(\alu_ctrl_i[FUNCT][0] ), .F(n25), 
        .Z(n29) );
  HS65_LH_AOI32X5 U23 ( .A(\alu_ctrl_i[FUNCT][3] ), .B(\alu_ctrl_i[FUNCT][0] ), 
        .C(\alu_ctrl_i[FUNCT][4] ), .D(n125), .E(n121), .Z(n30) );
  HS65_LH_NOR3X4 U24 ( .A(\alu_ctrl_i[FUNCT][3] ), .B(\alu_ctrl_i[FUNCT][5] ), 
        .C(\alu_ctrl_i[FUNCT][2] ), .Z(n26) );
  HS65_LH_NAND4ABX3 U25 ( .A(n122), .B(n34), .C(\alu_ctrl_i[FUNCT][5] ), .D(
        n22), .Z(n17) );
  HS65_LH_NAND3X5 U26 ( .A(n123), .B(n121), .C(\alu_ctrl_i[FUNCT][1] ), .Z(n34) );
  HS65_LH_IVX9 U27 ( .A(\alu_ctrl_i[FUNCT][0] ), .Z(n125) );
  HS65_LH_NAND3X5 U28 ( .A(n122), .B(n121), .C(\alu_ctrl_i[FUNCT][5] ), .Z(n25) );
  HS65_LH_CBI4I1X5 U29 ( .A(n118), .B(n11), .C(n116), .D(n12), .Z(
        \alu_ctrl_o[OP][4] ) );
  HS65_LH_NAND4ABX3 U30 ( .A(n13), .B(n14), .C(n125), .D(
        \alu_ctrl_i[FUNCT][3] ), .Z(n11) );
  HS65_LH_NAND4ABX3 U31 ( .A(\alu_ctrl_i[FUNCT][2] ), .B(
        \alu_ctrl_i[FUNCT][5] ), .C(n121), .D(n119), .Z(n14) );
  HS65_LH_NOR2X6 U32 ( .A(\alu_ctrl_i[OP][0] ), .B(\alu_ctrl_i[OP][3] ), .Z(
        n24) );
  HS65_LH_NAND3AX6 U33 ( .A(n33), .B(n26), .C(n35), .Z(n27) );
  HS65_LH_NOR3X4 U34 ( .A(n36), .B(\alu_ctrl_i[OP][0] ), .C(
        \alu_ctrl_i[FUNCT][0] ), .Z(n35) );
  HS65_LHS_XOR2X6 U35 ( .A(\alu_ctrl_i[FUNCT][4] ), .B(n124), .Z(n36) );
  HS65_LH_IVX9 U36 ( .A(\alu_ctrl_i[FUNCT][4] ), .Z(n121) );
  HS65_LH_NAND3AX6 U37 ( .A(\alu_ctrl_i[OP][3] ), .B(\alu_ctrl_i[OP][0] ), .C(
        \alu_ctrl_i[OP][1] ), .Z(n12) );
  HS65_LH_NAND3X5 U38 ( .A(n24), .B(n118), .C(\alu_ctrl_i[OP][1] ), .Z(n18) );
  HS65_LH_IVX9 U39 ( .A(\alu_ctrl_i[FUNCT][1] ), .Z(n124) );
  HS65_LH_IVX9 U40 ( .A(\alu_ctrl_i[OP][2] ), .Z(n118) );
  HS65_LH_IVX9 U41 ( .A(\alu_ctrl_i[FUNCT][2] ), .Z(n123) );
  HS65_LH_IVX9 U42 ( .A(\alu_ctrl_i[OP][1] ), .Z(n119) );
  HS65_LH_IVX9 U43 ( .A(\alu_ctrl_i[FUNCT][3] ), .Z(n122) );
endmodule


module exe_top_DW01_add_0 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [11:1] carry;

  HS65_LHS_XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Z(SUM[11]) );
  HS65_LH_FA1X4 U1_10 ( .A0(A[10]), .B0(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S0(SUM[10]) );
  HS65_LH_FA1X4 U1_9 ( .A0(A[9]), .B0(B[9]), .CI(carry[9]), .CO(carry[10]), 
        .S0(SUM[9]) );
  HS65_LH_FA1X4 U1_8 ( .A0(A[8]), .B0(B[8]), .CI(carry[8]), .CO(carry[9]), 
        .S0(SUM[8]) );
  HS65_LH_FA1X4 U1_7 ( .A0(A[7]), .B0(B[7]), .CI(carry[7]), .CO(carry[8]), 
        .S0(SUM[7]) );
  HS65_LH_FA1X4 U1_6 ( .A0(A[6]), .B0(B[6]), .CI(carry[6]), .CO(carry[7]), 
        .S0(SUM[6]) );
  HS65_LH_FA1X4 U1_5 ( .A0(A[5]), .B0(B[5]), .CI(carry[5]), .CO(carry[6]), 
        .S0(SUM[5]) );
  HS65_LH_FA1X4 U1_4 ( .A0(A[4]), .B0(B[4]), .CI(carry[4]), .CO(carry[5]), 
        .S0(SUM[4]) );
  HS65_LH_FA1X4 U1_3 ( .A0(A[3]), .B0(B[3]), .CI(carry[3]), .CO(carry[4]), 
        .S0(SUM[3]) );
  HS65_LH_FA1X4 U1_2 ( .A0(A[2]), .B0(B[2]), .CI(carry[2]), .CO(carry[3]), 
        .S0(SUM[2]) );
  HS65_LH_FA1X4 U1_1 ( .A0(A[1]), .B0(B[1]), .CI(n1), .CO(carry[2]), .S0(
        SUM[1]) );
  HS65_LH_AND2X4 U1 ( .A(A[0]), .B(B[0]), .Z(n1) );
  HS65_LHS_XOR2X6 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module exe_top ( clk, rst_n, .exe_top_i({\exe_top_i[SHAMT][4] , 
        \exe_top_i[SHAMT][3] , \exe_top_i[SHAMT][2] , \exe_top_i[SHAMT][1] , 
        \exe_top_i[SHAMT][0] , \exe_top_i[REGS_A][31] , 
        \exe_top_i[REGS_A][30] , \exe_top_i[REGS_A][29] , 
        \exe_top_i[REGS_A][28] , \exe_top_i[REGS_A][27] , 
        \exe_top_i[REGS_A][26] , \exe_top_i[REGS_A][25] , 
        \exe_top_i[REGS_A][24] , \exe_top_i[REGS_A][23] , 
        \exe_top_i[REGS_A][22] , \exe_top_i[REGS_A][21] , 
        \exe_top_i[REGS_A][20] , \exe_top_i[REGS_A][19] , 
        \exe_top_i[REGS_A][18] , \exe_top_i[REGS_A][17] , 
        \exe_top_i[REGS_A][16] , \exe_top_i[REGS_A][15] , 
        \exe_top_i[REGS_A][14] , \exe_top_i[REGS_A][13] , 
        \exe_top_i[REGS_A][12] , \exe_top_i[REGS_A][11] , 
        \exe_top_i[REGS_A][10] , \exe_top_i[REGS_A][9] , 
        \exe_top_i[REGS_A][8] , \exe_top_i[REGS_A][7] , \exe_top_i[REGS_A][6] , 
        \exe_top_i[REGS_A][5] , \exe_top_i[REGS_A][4] , \exe_top_i[REGS_A][3] , 
        \exe_top_i[REGS_A][2] , \exe_top_i[REGS_A][1] , \exe_top_i[REGS_A][0] , 
        \exe_top_i[REGS_B][31] , \exe_top_i[REGS_B][30] , 
        \exe_top_i[REGS_B][29] , \exe_top_i[REGS_B][28] , 
        \exe_top_i[REGS_B][27] , \exe_top_i[REGS_B][26] , 
        \exe_top_i[REGS_B][25] , \exe_top_i[REGS_B][24] , 
        \exe_top_i[REGS_B][23] , \exe_top_i[REGS_B][22] , 
        \exe_top_i[REGS_B][21] , \exe_top_i[REGS_B][20] , 
        \exe_top_i[REGS_B][19] , \exe_top_i[REGS_B][18] , 
        \exe_top_i[REGS_B][17] , \exe_top_i[REGS_B][16] , 
        \exe_top_i[REGS_B][15] , \exe_top_i[REGS_B][14] , 
        \exe_top_i[REGS_B][13] , \exe_top_i[REGS_B][12] , 
        \exe_top_i[REGS_B][11] , \exe_top_i[REGS_B][10] , 
        \exe_top_i[REGS_B][9] , \exe_top_i[REGS_B][8] , \exe_top_i[REGS_B][7] , 
        \exe_top_i[REGS_B][6] , \exe_top_i[REGS_B][5] , \exe_top_i[REGS_B][4] , 
        \exe_top_i[REGS_B][3] , \exe_top_i[REGS_B][2] , \exe_top_i[REGS_B][1] , 
        \exe_top_i[REGS_B][0] , \exe_top_i[ALU_SRC_B] , 
        \exe_top_i[IMMIDIATE][31] , \exe_top_i[IMMIDIATE][30] , 
        \exe_top_i[IMMIDIATE][29] , \exe_top_i[IMMIDIATE][28] , 
        \exe_top_i[IMMIDIATE][27] , \exe_top_i[IMMIDIATE][26] , 
        \exe_top_i[IMMIDIATE][25] , \exe_top_i[IMMIDIATE][24] , 
        \exe_top_i[IMMIDIATE][23] , \exe_top_i[IMMIDIATE][22] , 
        \exe_top_i[IMMIDIATE][21] , \exe_top_i[IMMIDIATE][20] , 
        \exe_top_i[IMMIDIATE][19] , \exe_top_i[IMMIDIATE][18] , 
        \exe_top_i[IMMIDIATE][17] , \exe_top_i[IMMIDIATE][16] , 
        \exe_top_i[IMMIDIATE][15] , \exe_top_i[IMMIDIATE][14] , 
        \exe_top_i[IMMIDIATE][13] , \exe_top_i[IMMIDIATE][12] , 
        \exe_top_i[IMMIDIATE][11] , \exe_top_i[IMMIDIATE][10] , 
        \exe_top_i[IMMIDIATE][9] , \exe_top_i[IMMIDIATE][8] , 
        \exe_top_i[IMMIDIATE][7] , \exe_top_i[IMMIDIATE][6] , 
        \exe_top_i[IMMIDIATE][5] , \exe_top_i[IMMIDIATE][4] , 
        \exe_top_i[IMMIDIATE][3] , \exe_top_i[IMMIDIATE][2] , 
        \exe_top_i[IMMIDIATE][1] , \exe_top_i[IMMIDIATE][0] , 
        \exe_top_i[OP][3] , \exe_top_i[OP][2] , \exe_top_i[OP][1] , 
        \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] , \exe_top_i[FUNCT][4] , 
        \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] , \exe_top_i[FUNCT][1] , 
        \exe_top_i[FUNCT][0] , \exe_top_i[PC_PLUS1][11] , 
        \exe_top_i[PC_PLUS1][10] , \exe_top_i[PC_PLUS1][9] , 
        \exe_top_i[PC_PLUS1][8] , \exe_top_i[PC_PLUS1][7] , 
        \exe_top_i[PC_PLUS1][6] , \exe_top_i[PC_PLUS1][5] , 
        \exe_top_i[PC_PLUS1][4] , \exe_top_i[PC_PLUS1][3] , 
        \exe_top_i[PC_PLUS1][2] , \exe_top_i[PC_PLUS1][1] , 
        \exe_top_i[PC_PLUS1][0] , \exe_top_i[REGDST] , \exe_top_i[RT][4] , 
        \exe_top_i[RT][3] , \exe_top_i[RT][2] , \exe_top_i[RT][1] , 
        \exe_top_i[RT][0] , \exe_top_i[RD][4] , \exe_top_i[RD][3] , 
        \exe_top_i[RD][2] , \exe_top_i[RD][1] , \exe_top_i[RD][0] }), 
    .exe_top_o({\exe_top_o[BRANCH] , \exe_top_o[BRANCH_PC][11] , 
        \exe_top_o[BRANCH_PC][10] , \exe_top_o[BRANCH_PC][9] , 
        \exe_top_o[BRANCH_PC][8] , \exe_top_o[BRANCH_PC][7] , 
        \exe_top_o[BRANCH_PC][6] , \exe_top_o[BRANCH_PC][5] , 
        \exe_top_o[BRANCH_PC][4] , \exe_top_o[BRANCH_PC][3] , 
        \exe_top_o[BRANCH_PC][2] , \exe_top_o[BRANCH_PC][1] , 
        \exe_top_o[BRANCH_PC][0] , \exe_top_o[RESULT][31] , 
        \exe_top_o[RESULT][30] , \exe_top_o[RESULT][29] , 
        \exe_top_o[RESULT][28] , \exe_top_o[RESULT][27] , 
        \exe_top_o[RESULT][26] , \exe_top_o[RESULT][25] , 
        \exe_top_o[RESULT][24] , \exe_top_o[RESULT][23] , 
        \exe_top_o[RESULT][22] , \exe_top_o[RESULT][21] , 
        \exe_top_o[RESULT][20] , \exe_top_o[RESULT][19] , 
        \exe_top_o[RESULT][18] , \exe_top_o[RESULT][17] , 
        \exe_top_o[RESULT][16] , \exe_top_o[RESULT][15] , 
        \exe_top_o[RESULT][14] , \exe_top_o[RESULT][13] , 
        \exe_top_o[RESULT][12] , \exe_top_o[RESULT][11] , 
        \exe_top_o[RESULT][10] , \exe_top_o[RESULT][9] , 
        \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] , \exe_top_o[RESULT][6] , 
        \exe_top_o[RESULT][5] , \exe_top_o[RESULT][4] , \exe_top_o[RESULT][3] , 
        \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] , \exe_top_o[RESULT][0] , 
        \exe_top_o[WRITE_REG][4] , \exe_top_o[WRITE_REG][3] , 
        \exe_top_o[WRITE_REG][2] , \exe_top_o[WRITE_REG][1] , 
        \exe_top_o[WRITE_REG][0] , \exe_top_o[DMEM_DATA][31] , 
        \exe_top_o[DMEM_DATA][30] , \exe_top_o[DMEM_DATA][29] , 
        \exe_top_o[DMEM_DATA][28] , \exe_top_o[DMEM_DATA][27] , 
        \exe_top_o[DMEM_DATA][26] , \exe_top_o[DMEM_DATA][25] , 
        \exe_top_o[DMEM_DATA][24] , \exe_top_o[DMEM_DATA][23] , 
        \exe_top_o[DMEM_DATA][22] , \exe_top_o[DMEM_DATA][21] , 
        \exe_top_o[DMEM_DATA][20] , \exe_top_o[DMEM_DATA][19] , 
        \exe_top_o[DMEM_DATA][18] , \exe_top_o[DMEM_DATA][17] , 
        \exe_top_o[DMEM_DATA][16] , \exe_top_o[DMEM_DATA][15] , 
        \exe_top_o[DMEM_DATA][14] , \exe_top_o[DMEM_DATA][13] , 
        \exe_top_o[DMEM_DATA][12] , \exe_top_o[DMEM_DATA][11] , 
        \exe_top_o[DMEM_DATA][10] , \exe_top_o[DMEM_DATA][9] , 
        \exe_top_o[DMEM_DATA][8] , \exe_top_o[DMEM_DATA][7] , 
        \exe_top_o[DMEM_DATA][6] , \exe_top_o[DMEM_DATA][5] , 
        \exe_top_o[DMEM_DATA][4] , \exe_top_o[DMEM_DATA][3] , 
        \exe_top_o[DMEM_DATA][2] , \exe_top_o[DMEM_DATA][1] , 
        \exe_top_o[DMEM_DATA][0] }) );
  input clk, rst_n, \exe_top_i[SHAMT][4] , \exe_top_i[SHAMT][3] ,
         \exe_top_i[SHAMT][2] , \exe_top_i[SHAMT][1] , \exe_top_i[SHAMT][0] ,
         \exe_top_i[REGS_A][31] , \exe_top_i[REGS_A][30] ,
         \exe_top_i[REGS_A][29] , \exe_top_i[REGS_A][28] ,
         \exe_top_i[REGS_A][27] , \exe_top_i[REGS_A][26] ,
         \exe_top_i[REGS_A][25] , \exe_top_i[REGS_A][24] ,
         \exe_top_i[REGS_A][23] , \exe_top_i[REGS_A][22] ,
         \exe_top_i[REGS_A][21] , \exe_top_i[REGS_A][20] ,
         \exe_top_i[REGS_A][19] , \exe_top_i[REGS_A][18] ,
         \exe_top_i[REGS_A][17] , \exe_top_i[REGS_A][16] ,
         \exe_top_i[REGS_A][15] , \exe_top_i[REGS_A][14] ,
         \exe_top_i[REGS_A][13] , \exe_top_i[REGS_A][12] ,
         \exe_top_i[REGS_A][11] , \exe_top_i[REGS_A][10] ,
         \exe_top_i[REGS_A][9] , \exe_top_i[REGS_A][8] ,
         \exe_top_i[REGS_A][7] , \exe_top_i[REGS_A][6] ,
         \exe_top_i[REGS_A][5] , \exe_top_i[REGS_A][4] ,
         \exe_top_i[REGS_A][3] , \exe_top_i[REGS_A][2] ,
         \exe_top_i[REGS_A][1] , \exe_top_i[REGS_A][0] ,
         \exe_top_i[REGS_B][31] , \exe_top_i[REGS_B][30] ,
         \exe_top_i[REGS_B][29] , \exe_top_i[REGS_B][28] ,
         \exe_top_i[REGS_B][27] , \exe_top_i[REGS_B][26] ,
         \exe_top_i[REGS_B][25] , \exe_top_i[REGS_B][24] ,
         \exe_top_i[REGS_B][23] , \exe_top_i[REGS_B][22] ,
         \exe_top_i[REGS_B][21] , \exe_top_i[REGS_B][20] ,
         \exe_top_i[REGS_B][19] , \exe_top_i[REGS_B][18] ,
         \exe_top_i[REGS_B][17] , \exe_top_i[REGS_B][16] ,
         \exe_top_i[REGS_B][15] , \exe_top_i[REGS_B][14] ,
         \exe_top_i[REGS_B][13] , \exe_top_i[REGS_B][12] ,
         \exe_top_i[REGS_B][11] , \exe_top_i[REGS_B][10] ,
         \exe_top_i[REGS_B][9] , \exe_top_i[REGS_B][8] ,
         \exe_top_i[REGS_B][7] , \exe_top_i[REGS_B][6] ,
         \exe_top_i[REGS_B][5] , \exe_top_i[REGS_B][4] ,
         \exe_top_i[REGS_B][3] , \exe_top_i[REGS_B][2] ,
         \exe_top_i[REGS_B][1] , \exe_top_i[REGS_B][0] ,
         \exe_top_i[ALU_SRC_B] , \exe_top_i[IMMIDIATE][31] ,
         \exe_top_i[IMMIDIATE][30] , \exe_top_i[IMMIDIATE][29] ,
         \exe_top_i[IMMIDIATE][28] , \exe_top_i[IMMIDIATE][27] ,
         \exe_top_i[IMMIDIATE][26] , \exe_top_i[IMMIDIATE][25] ,
         \exe_top_i[IMMIDIATE][24] , \exe_top_i[IMMIDIATE][23] ,
         \exe_top_i[IMMIDIATE][22] , \exe_top_i[IMMIDIATE][21] ,
         \exe_top_i[IMMIDIATE][20] , \exe_top_i[IMMIDIATE][19] ,
         \exe_top_i[IMMIDIATE][18] , \exe_top_i[IMMIDIATE][17] ,
         \exe_top_i[IMMIDIATE][16] , \exe_top_i[IMMIDIATE][15] ,
         \exe_top_i[IMMIDIATE][14] , \exe_top_i[IMMIDIATE][13] ,
         \exe_top_i[IMMIDIATE][12] , \exe_top_i[IMMIDIATE][11] ,
         \exe_top_i[IMMIDIATE][10] , \exe_top_i[IMMIDIATE][9] ,
         \exe_top_i[IMMIDIATE][8] , \exe_top_i[IMMIDIATE][7] ,
         \exe_top_i[IMMIDIATE][6] , \exe_top_i[IMMIDIATE][5] ,
         \exe_top_i[IMMIDIATE][4] , \exe_top_i[IMMIDIATE][3] ,
         \exe_top_i[IMMIDIATE][2] , \exe_top_i[IMMIDIATE][1] ,
         \exe_top_i[IMMIDIATE][0] , \exe_top_i[OP][3] , \exe_top_i[OP][2] ,
         \exe_top_i[OP][1] , \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] ,
         \exe_top_i[FUNCT][4] , \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] ,
         \exe_top_i[FUNCT][1] , \exe_top_i[FUNCT][0] ,
         \exe_top_i[PC_PLUS1][11] , \exe_top_i[PC_PLUS1][10] ,
         \exe_top_i[PC_PLUS1][9] , \exe_top_i[PC_PLUS1][8] ,
         \exe_top_i[PC_PLUS1][7] , \exe_top_i[PC_PLUS1][6] ,
         \exe_top_i[PC_PLUS1][5] , \exe_top_i[PC_PLUS1][4] ,
         \exe_top_i[PC_PLUS1][3] , \exe_top_i[PC_PLUS1][2] ,
         \exe_top_i[PC_PLUS1][1] , \exe_top_i[PC_PLUS1][0] ,
         \exe_top_i[REGDST] , \exe_top_i[RT][4] , \exe_top_i[RT][3] ,
         \exe_top_i[RT][2] , \exe_top_i[RT][1] , \exe_top_i[RT][0] ,
         \exe_top_i[RD][4] , \exe_top_i[RD][3] , \exe_top_i[RD][2] ,
         \exe_top_i[RD][1] , \exe_top_i[RD][0] ;
  output \exe_top_o[BRANCH] , \exe_top_o[BRANCH_PC][11] ,
         \exe_top_o[BRANCH_PC][10] , \exe_top_o[BRANCH_PC][9] ,
         \exe_top_o[BRANCH_PC][8] , \exe_top_o[BRANCH_PC][7] ,
         \exe_top_o[BRANCH_PC][6] , \exe_top_o[BRANCH_PC][5] ,
         \exe_top_o[BRANCH_PC][4] , \exe_top_o[BRANCH_PC][3] ,
         \exe_top_o[BRANCH_PC][2] , \exe_top_o[BRANCH_PC][1] ,
         \exe_top_o[BRANCH_PC][0] , \exe_top_o[RESULT][31] ,
         \exe_top_o[RESULT][30] , \exe_top_o[RESULT][29] ,
         \exe_top_o[RESULT][28] , \exe_top_o[RESULT][27] ,
         \exe_top_o[RESULT][26] , \exe_top_o[RESULT][25] ,
         \exe_top_o[RESULT][24] , \exe_top_o[RESULT][23] ,
         \exe_top_o[RESULT][22] , \exe_top_o[RESULT][21] ,
         \exe_top_o[RESULT][20] , \exe_top_o[RESULT][19] ,
         \exe_top_o[RESULT][18] , \exe_top_o[RESULT][17] ,
         \exe_top_o[RESULT][16] , \exe_top_o[RESULT][15] ,
         \exe_top_o[RESULT][14] , \exe_top_o[RESULT][13] ,
         \exe_top_o[RESULT][12] , \exe_top_o[RESULT][11] ,
         \exe_top_o[RESULT][10] , \exe_top_o[RESULT][9] ,
         \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] ,
         \exe_top_o[RESULT][6] , \exe_top_o[RESULT][5] ,
         \exe_top_o[RESULT][4] , \exe_top_o[RESULT][3] ,
         \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] ,
         \exe_top_o[RESULT][0] , \exe_top_o[WRITE_REG][4] ,
         \exe_top_o[WRITE_REG][3] , \exe_top_o[WRITE_REG][2] ,
         \exe_top_o[WRITE_REG][1] , \exe_top_o[WRITE_REG][0] ,
         \exe_top_o[DMEM_DATA][31] , \exe_top_o[DMEM_DATA][30] ,
         \exe_top_o[DMEM_DATA][29] , \exe_top_o[DMEM_DATA][28] ,
         \exe_top_o[DMEM_DATA][27] , \exe_top_o[DMEM_DATA][26] ,
         \exe_top_o[DMEM_DATA][25] , \exe_top_o[DMEM_DATA][24] ,
         \exe_top_o[DMEM_DATA][23] , \exe_top_o[DMEM_DATA][22] ,
         \exe_top_o[DMEM_DATA][21] , \exe_top_o[DMEM_DATA][20] ,
         \exe_top_o[DMEM_DATA][19] , \exe_top_o[DMEM_DATA][18] ,
         \exe_top_o[DMEM_DATA][17] , \exe_top_o[DMEM_DATA][16] ,
         \exe_top_o[DMEM_DATA][15] , \exe_top_o[DMEM_DATA][14] ,
         \exe_top_o[DMEM_DATA][13] , \exe_top_o[DMEM_DATA][12] ,
         \exe_top_o[DMEM_DATA][11] , \exe_top_o[DMEM_DATA][10] ,
         \exe_top_o[DMEM_DATA][9] , \exe_top_o[DMEM_DATA][8] ,
         \exe_top_o[DMEM_DATA][7] , \exe_top_o[DMEM_DATA][6] ,
         \exe_top_o[DMEM_DATA][5] , \exe_top_o[DMEM_DATA][4] ,
         \exe_top_o[DMEM_DATA][3] , \exe_top_o[DMEM_DATA][2] ,
         \exe_top_o[DMEM_DATA][1] , \exe_top_o[DMEM_DATA][0] ;
  wire   \exe_top_o[DMEM_DATA][31] , \exe_top_o[DMEM_DATA][30] ,
         \exe_top_o[DMEM_DATA][29] , \exe_top_o[DMEM_DATA][28] ,
         \exe_top_o[DMEM_DATA][27] , \exe_top_o[DMEM_DATA][26] ,
         \exe_top_o[DMEM_DATA][25] , \exe_top_o[DMEM_DATA][24] ,
         \exe_top_o[DMEM_DATA][23] , \exe_top_o[DMEM_DATA][22] ,
         \exe_top_o[DMEM_DATA][21] , \exe_top_o[DMEM_DATA][20] ,
         \exe_top_o[DMEM_DATA][19] , \exe_top_o[DMEM_DATA][18] ,
         \exe_top_o[DMEM_DATA][17] , \exe_top_o[DMEM_DATA][16] ,
         \exe_top_o[DMEM_DATA][15] , \exe_top_o[DMEM_DATA][14] ,
         \exe_top_o[DMEM_DATA][13] , \exe_top_o[DMEM_DATA][12] ,
         \exe_top_o[DMEM_DATA][11] , \exe_top_o[DMEM_DATA][10] ,
         \exe_top_o[DMEM_DATA][9] , \exe_top_o[DMEM_DATA][8] ,
         \exe_top_o[DMEM_DATA][7] , \exe_top_o[DMEM_DATA][6] ,
         \exe_top_o[DMEM_DATA][5] , \exe_top_o[DMEM_DATA][4] ,
         \exe_top_o[DMEM_DATA][3] , \exe_top_o[DMEM_DATA][2] ,
         \exe_top_o[DMEM_DATA][1] , \exe_top_o[DMEM_DATA][0] , n6, n7, n8;
  wire   [31:0] src_b;
  wire   [4:0] op_aluCtrl_alu;
  assign \exe_top_o[DMEM_DATA][31]  = \exe_top_i[REGS_B][31] ;
  assign \exe_top_o[DMEM_DATA][30]  = \exe_top_i[REGS_B][30] ;
  assign \exe_top_o[DMEM_DATA][29]  = \exe_top_i[REGS_B][29] ;
  assign \exe_top_o[DMEM_DATA][28]  = \exe_top_i[REGS_B][28] ;
  assign \exe_top_o[DMEM_DATA][27]  = \exe_top_i[REGS_B][27] ;
  assign \exe_top_o[DMEM_DATA][26]  = \exe_top_i[REGS_B][26] ;
  assign \exe_top_o[DMEM_DATA][25]  = \exe_top_i[REGS_B][25] ;
  assign \exe_top_o[DMEM_DATA][24]  = \exe_top_i[REGS_B][24] ;
  assign \exe_top_o[DMEM_DATA][23]  = \exe_top_i[REGS_B][23] ;
  assign \exe_top_o[DMEM_DATA][22]  = \exe_top_i[REGS_B][22] ;
  assign \exe_top_o[DMEM_DATA][21]  = \exe_top_i[REGS_B][21] ;
  assign \exe_top_o[DMEM_DATA][20]  = \exe_top_i[REGS_B][20] ;
  assign \exe_top_o[DMEM_DATA][19]  = \exe_top_i[REGS_B][19] ;
  assign \exe_top_o[DMEM_DATA][18]  = \exe_top_i[REGS_B][18] ;
  assign \exe_top_o[DMEM_DATA][17]  = \exe_top_i[REGS_B][17] ;
  assign \exe_top_o[DMEM_DATA][16]  = \exe_top_i[REGS_B][16] ;
  assign \exe_top_o[DMEM_DATA][15]  = \exe_top_i[REGS_B][15] ;
  assign \exe_top_o[DMEM_DATA][14]  = \exe_top_i[REGS_B][14] ;
  assign \exe_top_o[DMEM_DATA][13]  = \exe_top_i[REGS_B][13] ;
  assign \exe_top_o[DMEM_DATA][12]  = \exe_top_i[REGS_B][12] ;
  assign \exe_top_o[DMEM_DATA][11]  = \exe_top_i[REGS_B][11] ;
  assign \exe_top_o[DMEM_DATA][10]  = \exe_top_i[REGS_B][10] ;
  assign \exe_top_o[DMEM_DATA][9]  = \exe_top_i[REGS_B][9] ;
  assign \exe_top_o[DMEM_DATA][8]  = \exe_top_i[REGS_B][8] ;
  assign \exe_top_o[DMEM_DATA][7]  = \exe_top_i[REGS_B][7] ;
  assign \exe_top_o[DMEM_DATA][6]  = \exe_top_i[REGS_B][6] ;
  assign \exe_top_o[DMEM_DATA][5]  = \exe_top_i[REGS_B][5] ;
  assign \exe_top_o[DMEM_DATA][4]  = \exe_top_i[REGS_B][4] ;
  assign \exe_top_o[DMEM_DATA][3]  = \exe_top_i[REGS_B][3] ;
  assign \exe_top_o[DMEM_DATA][2]  = \exe_top_i[REGS_B][2] ;
  assign \exe_top_o[DMEM_DATA][1]  = \exe_top_i[REGS_B][1] ;
  assign \exe_top_o[DMEM_DATA][0]  = \exe_top_i[REGS_B][0] ;

  alu alu_inst ( .clk(clk), .rst_n(rst_n), .alu_i({\exe_top_i[REGS_A][31] , 
        \exe_top_i[REGS_A][30] , \exe_top_i[REGS_A][29] , 
        \exe_top_i[REGS_A][28] , \exe_top_i[REGS_A][27] , 
        \exe_top_i[REGS_A][26] , \exe_top_i[REGS_A][25] , 
        \exe_top_i[REGS_A][24] , \exe_top_i[REGS_A][23] , 
        \exe_top_i[REGS_A][22] , \exe_top_i[REGS_A][21] , 
        \exe_top_i[REGS_A][20] , \exe_top_i[REGS_A][19] , 
        \exe_top_i[REGS_A][18] , \exe_top_i[REGS_A][17] , 
        \exe_top_i[REGS_A][16] , \exe_top_i[REGS_A][15] , 
        \exe_top_i[REGS_A][14] , \exe_top_i[REGS_A][13] , 
        \exe_top_i[REGS_A][12] , \exe_top_i[REGS_A][11] , 
        \exe_top_i[REGS_A][10] , \exe_top_i[REGS_A][9] , 
        \exe_top_i[REGS_A][8] , \exe_top_i[REGS_A][7] , \exe_top_i[REGS_A][6] , 
        \exe_top_i[REGS_A][5] , \exe_top_i[REGS_A][4] , \exe_top_i[REGS_A][3] , 
        \exe_top_i[REGS_A][2] , \exe_top_i[REGS_A][1] , \exe_top_i[REGS_A][0] , 
        src_b, op_aluCtrl_alu, \exe_top_i[SHAMT][4] , \exe_top_i[SHAMT][3] , 
        \exe_top_i[SHAMT][2] , \exe_top_i[SHAMT][1] , \exe_top_i[SHAMT][0] }), 
        .alu_o({\exe_top_o[BRANCH] , \exe_top_o[RESULT][31] , 
        \exe_top_o[RESULT][30] , \exe_top_o[RESULT][29] , 
        \exe_top_o[RESULT][28] , \exe_top_o[RESULT][27] , 
        \exe_top_o[RESULT][26] , \exe_top_o[RESULT][25] , 
        \exe_top_o[RESULT][24] , \exe_top_o[RESULT][23] , 
        \exe_top_o[RESULT][22] , \exe_top_o[RESULT][21] , 
        \exe_top_o[RESULT][20] , \exe_top_o[RESULT][19] , 
        \exe_top_o[RESULT][18] , \exe_top_o[RESULT][17] , 
        \exe_top_o[RESULT][16] , \exe_top_o[RESULT][15] , 
        \exe_top_o[RESULT][14] , \exe_top_o[RESULT][13] , 
        \exe_top_o[RESULT][12] , \exe_top_o[RESULT][11] , 
        \exe_top_o[RESULT][10] , \exe_top_o[RESULT][9] , 
        \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] , \exe_top_o[RESULT][6] , 
        \exe_top_o[RESULT][5] , \exe_top_o[RESULT][4] , \exe_top_o[RESULT][3] , 
        \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] , \exe_top_o[RESULT][0] }) );
  alu_ctrl alu_ctrl_inst ( .alu_ctrl_i({\exe_top_i[OP][3] , \exe_top_i[OP][2] , 
        \exe_top_i[OP][1] , \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] , 
        \exe_top_i[FUNCT][4] , \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] , 
        \exe_top_i[FUNCT][1] , \exe_top_i[FUNCT][0] }), .alu_ctrl_o(
        op_aluCtrl_alu) );
  exe_top_DW01_add_0 add_43 ( .A({\exe_top_i[PC_PLUS1][11] , 
        \exe_top_i[PC_PLUS1][10] , \exe_top_i[PC_PLUS1][9] , 
        \exe_top_i[PC_PLUS1][8] , \exe_top_i[PC_PLUS1][7] , 
        \exe_top_i[PC_PLUS1][6] , \exe_top_i[PC_PLUS1][5] , 
        \exe_top_i[PC_PLUS1][4] , \exe_top_i[PC_PLUS1][3] , 
        \exe_top_i[PC_PLUS1][2] , \exe_top_i[PC_PLUS1][1] , 
        \exe_top_i[PC_PLUS1][0] }), .B({\exe_top_i[IMMIDIATE][11] , 
        \exe_top_i[IMMIDIATE][10] , \exe_top_i[IMMIDIATE][9] , 
        \exe_top_i[IMMIDIATE][8] , \exe_top_i[IMMIDIATE][7] , 
        \exe_top_i[IMMIDIATE][6] , \exe_top_i[IMMIDIATE][5] , 
        \exe_top_i[IMMIDIATE][4] , \exe_top_i[IMMIDIATE][3] , 
        \exe_top_i[IMMIDIATE][2] , \exe_top_i[IMMIDIATE][1] , 
        \exe_top_i[IMMIDIATE][0] }), .CI(1'b0), .SUM({
        \exe_top_o[BRANCH_PC][11] , \exe_top_o[BRANCH_PC][10] , 
        \exe_top_o[BRANCH_PC][9] , \exe_top_o[BRANCH_PC][8] , 
        \exe_top_o[BRANCH_PC][7] , \exe_top_o[BRANCH_PC][6] , 
        \exe_top_o[BRANCH_PC][5] , \exe_top_o[BRANCH_PC][4] , 
        \exe_top_o[BRANCH_PC][3] , \exe_top_o[BRANCH_PC][2] , 
        \exe_top_o[BRANCH_PC][1] , \exe_top_o[BRANCH_PC][0] }) );
  HS65_LH_AO22X9 U42 ( .A(\exe_top_i[IMMIDIATE][19] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][19] ), .D(n6), .Z(
        src_b[19]) );
  HS65_LH_AO22X9 U43 ( .A(\exe_top_i[IMMIDIATE][27] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][27] ), .D(n7), .Z(
        src_b[27]) );
  HS65_LH_AO22X9 U44 ( .A(\exe_top_i[IMMIDIATE][25] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][25] ), .D(n7), .Z(
        src_b[25]) );
  HS65_LH_AO22X9 U45 ( .A(\exe_top_i[IMMIDIATE][12] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][12] ), .D(n6), .Z(
        src_b[12]) );
  HS65_LH_AO22X9 U46 ( .A(\exe_top_i[IMMIDIATE][15] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][15] ), .D(n6), .Z(
        src_b[15]) );
  HS65_LH_AO22X9 U47 ( .A(\exe_top_i[IMMIDIATE][13] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][13] ), .D(n6), .Z(
        src_b[13]) );
  HS65_LH_AO22X9 U48 ( .A(\exe_top_i[IMMIDIATE][4] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][4] ), .D(n6), .Z(
        src_b[4]) );
  HS65_LH_AO22X9 U49 ( .A(\exe_top_i[IMMIDIATE][18] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][18] ), .D(n6), .Z(
        src_b[18]) );
  HS65_LH_AO22X9 U50 ( .A(\exe_top_i[IMMIDIATE][5] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][5] ), .D(n7), .Z(
        src_b[5]) );
  HS65_LH_AO22X9 U51 ( .A(\exe_top_i[IMMIDIATE][26] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][26] ), .D(n7), .Z(
        src_b[26]) );
  HS65_LH_AO22X9 U52 ( .A(\exe_top_i[IMMIDIATE][17] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][17] ), .D(n6), .Z(
        src_b[17]) );
  HS65_LH_AO22X9 U53 ( .A(\exe_top_i[IMMIDIATE][24] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][24] ), .D(n7), .Z(
        src_b[24]) );
  HS65_LH_AO22X9 U54 ( .A(\exe_top_i[IMMIDIATE][20] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][20] ), .D(n7), .Z(
        src_b[20]) );
  HS65_LH_AO22X9 U55 ( .A(\exe_top_i[IMMIDIATE][7] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][7] ), .D(n6), .Z(
        src_b[7]) );
  HS65_LH_AO22X9 U56 ( .A(\exe_top_i[IMMIDIATE][11] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][11] ), .D(n6), .Z(
        src_b[11]) );
  HS65_LH_AO22X9 U57 ( .A(\exe_top_i[IMMIDIATE][21] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][21] ), .D(n7), .Z(
        src_b[21]) );
  HS65_LH_AO22X9 U58 ( .A(\exe_top_i[IMMIDIATE][9] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][9] ), .D(n7), .Z(
        src_b[9]) );
  HS65_LH_AO22X9 U59 ( .A(\exe_top_i[IMMIDIATE][28] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][28] ), .D(n7), .Z(
        src_b[28]) );
  HS65_LH_AO22X9 U60 ( .A(\exe_top_i[IMMIDIATE][0] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][0] ), .D(n6), .Z(
        src_b[0]) );
  HS65_LH_AO22X9 U61 ( .A(\exe_top_i[IMMIDIATE][31] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][31] ), .D(n6), .Z(
        src_b[31]) );
  HS65_LH_AO22X9 U62 ( .A(\exe_top_i[IMMIDIATE][1] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][1] ), .D(n6), .Z(
        src_b[1]) );
  HS65_LH_AO22X9 U63 ( .A(\exe_top_i[IMMIDIATE][30] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][30] ), .D(n7), .Z(
        src_b[30]) );
  HS65_LH_AO22X9 U64 ( .A(\exe_top_i[IMMIDIATE][22] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][22] ), .D(n7), .Z(
        src_b[22]) );
  HS65_LH_AO22X9 U65 ( .A(\exe_top_i[IMMIDIATE][23] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][23] ), .D(n7), .Z(
        src_b[23]) );
  HS65_LH_AO22X9 U66 ( .A(\exe_top_i[IMMIDIATE][29] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][29] ), .D(n7), .Z(
        src_b[29]) );
  HS65_LH_AO22X9 U67 ( .A(\exe_top_i[IMMIDIATE][2] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][2] ), .D(n7), .Z(
        src_b[2]) );
  HS65_LH_AO22X9 U68 ( .A(\exe_top_i[IMMIDIATE][3] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][3] ), .D(n7), .Z(
        src_b[3]) );
  HS65_LH_AO22X9 U69 ( .A(\exe_top_i[IMMIDIATE][14] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][14] ), .D(n6), .Z(
        src_b[14]) );
  HS65_LH_AO22X9 U70 ( .A(\exe_top_i[IMMIDIATE][6] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][6] ), .D(n6), .Z(
        src_b[6]) );
  HS65_LH_AO22X9 U71 ( .A(\exe_top_i[IMMIDIATE][10] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][10] ), .D(n6), .Z(
        src_b[10]) );
  HS65_LH_AO22X9 U72 ( .A(\exe_top_i[IMMIDIATE][8] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][8] ), .D(n7), .Z(
        src_b[8]) );
  HS65_LH_AO22X9 U73 ( .A(\exe_top_i[IMMIDIATE][16] ), .B(
        \exe_top_i[ALU_SRC_B] ), .C(\exe_top_o[DMEM_DATA][16] ), .D(n6), .Z(
        src_b[16]) );
  HS65_LH_IVX9 U74 ( .A(\exe_top_i[REGDST] ), .Z(n8) );
  HS65_LH_AO22X9 U75 ( .A(\exe_top_i[RT][0] ), .B(n8), .C(\exe_top_i[RD][0] ), 
        .D(\exe_top_i[REGDST] ), .Z(\exe_top_o[WRITE_REG][0] ) );
  HS65_LH_AO22X9 U76 ( .A(\exe_top_i[RT][1] ), .B(n8), .C(\exe_top_i[RD][1] ), 
        .D(\exe_top_i[REGDST] ), .Z(\exe_top_o[WRITE_REG][1] ) );
  HS65_LH_AO22X9 U77 ( .A(\exe_top_i[RT][2] ), .B(n8), .C(\exe_top_i[RD][2] ), 
        .D(\exe_top_i[REGDST] ), .Z(\exe_top_o[WRITE_REG][2] ) );
  HS65_LH_AO22X9 U78 ( .A(\exe_top_i[RT][3] ), .B(n8), .C(\exe_top_i[RD][3] ), 
        .D(\exe_top_i[REGDST] ), .Z(\exe_top_o[WRITE_REG][3] ) );
  HS65_LH_AO22X9 U79 ( .A(\exe_top_i[RT][4] ), .B(n8), .C(\exe_top_i[REGDST] ), 
        .D(\exe_top_i[RD][4] ), .Z(\exe_top_o[WRITE_REG][4] ) );
  HS65_LH_IVX9 U80 ( .A(\exe_top_i[ALU_SRC_B] ), .Z(n6) );
  HS65_LH_IVX9 U81 ( .A(\exe_top_i[ALU_SRC_B] ), .Z(n7) );
endmodule

