VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
 MACRO prCellClass STRING ;
 MACRO prCellType STRING ;
 MACRO symmetry STRING ;
END PROPERTYDEFINITIONS

UNITS
 DATABASE MICRONS 1000 ;
END UNITS

MACRO ST_SPHDL_1024x32m8_L
 CLASS BLOCK ;
   SIZE 304.800 BY 99.400 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.250 0.050 148.350 0.570 ;
   LAYER M3 ;
    RECT 148.250 0.050 148.350 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.850 0.050 148.950 0.570 ;
   LAYER M3 ;
    RECT 148.850 0.050 148.950 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 149.450 0.050 149.550 0.570 ;
   LAYER M3 ;
    RECT 149.450 0.050 149.550 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 155.850 0.050 155.950 0.570 ;
   LAYER M3 ;
    RECT 155.850 0.050 155.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 156.450 0.050 156.550 0.570 ;
   LAYER M3 ;
    RECT 156.450 0.050 156.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 150.250 0.050 150.350 0.570 ;
   LAYER M3 ;
    RECT 150.250 0.050 150.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 151.850 0.050 151.950 0.570 ;
   LAYER M3 ;
    RECT 151.850 0.050 151.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN A[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 146.050 0.050 146.150 0.570 ;
   LAYER M3 ;
    RECT 146.050 0.050 146.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.916 LAYER M2 ;
  ANTENNAMAXAREACAR 13.057 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.347 LAYER M3 ;
 END A[7]
 PIN A[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 147.450 0.050 147.550 0.570 ;
   LAYER M3 ;
    RECT 147.450 0.050 147.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.924 LAYER M2 ;
  ANTENNAMAXAREACAR 13.892 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.282 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.376 LAYER M3 ;
 END A[8]
 PIN A[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 137.450 0.050 137.550 0.570 ;
   LAYER M3 ;
    RECT 137.450 0.050 137.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.251 LAYER M2 ;
  ANTENNAGATEAREA 0.251 LAYER M3 ;
  ANTENNAMAXAREACAR 3.203 LAYER M2 ;
  ANTENNAMAXAREACAR 9.213 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.586 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.511 LAYER M3 ;
 END A[9]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 160.650 0.050 160.750 0.570 ;
   LAYER M3 ;
    RECT 160.650 0.050 160.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 162.050 0.050 162.150 0.570 ;
   LAYER M3 ;
    RECT 162.050 0.050 162.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 91.250 0.050 91.350 0.570 ;
   LAYER M3 ;
    RECT 91.250 0.050 91.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[10]
 PIN D[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 95.450 0.050 95.550 0.570 ;
   LAYER M3 ;
    RECT 95.450 0.050 95.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[11]
 PIN D[12]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 108.050 0.050 108.150 0.570 ;
   LAYER M3 ;
    RECT 108.050 0.050 108.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[12]
 PIN D[13]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 112.250 0.050 112.350 0.570 ;
   LAYER M3 ;
    RECT 112.250 0.050 112.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[13]
 PIN D[14]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 124.850 0.050 124.950 0.570 ;
   LAYER M3 ;
    RECT 124.850 0.050 124.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[14]
 PIN D[15]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 129.050 0.050 129.150 0.570 ;
   LAYER M3 ;
    RECT 129.050 0.050 129.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[15]
 PIN D[16]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 174.250 0.050 174.350 0.570 ;
   LAYER M3 ;
    RECT 174.250 0.050 174.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[16]
 PIN D[17]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 178.250 0.050 178.350 0.570 ;
   LAYER M3 ;
    RECT 178.250 0.050 178.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[17]
 PIN D[18]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 191.050 0.050 191.150 0.570 ;
   LAYER M3 ;
    RECT 191.050 0.050 191.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[18]
 PIN D[19]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 195.050 0.050 195.150 0.570 ;
   LAYER M3 ;
    RECT 195.050 0.050 195.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[19]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[20]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 207.850 0.050 207.950 0.570 ;
   LAYER M3 ;
    RECT 207.850 0.050 207.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[20]
 PIN D[21]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 211.850 0.050 211.950 0.570 ;
   LAYER M3 ;
    RECT 211.850 0.050 211.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[21]
 PIN D[22]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 224.650 0.050 224.750 0.570 ;
   LAYER M3 ;
    RECT 224.650 0.050 224.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[22]
 PIN D[23]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 228.650 0.050 228.750 0.570 ;
   LAYER M3 ;
    RECT 228.650 0.050 228.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[23]
 PIN D[24]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 241.450 0.050 241.550 0.570 ;
   LAYER M3 ;
    RECT 241.450 0.050 241.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[24]
 PIN D[25]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 245.450 0.050 245.550 0.570 ;
   LAYER M3 ;
    RECT 245.450 0.050 245.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[25]
 PIN D[26]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 258.250 0.050 258.350 0.570 ;
   LAYER M3 ;
    RECT 258.250 0.050 258.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[26]
 PIN D[27]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 262.250 0.050 262.350 0.570 ;
   LAYER M3 ;
    RECT 262.250 0.050 262.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[27]
 PIN D[28]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 275.050 0.050 275.150 0.570 ;
   LAYER M3 ;
    RECT 275.050 0.050 275.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[28]
 PIN D[29]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 279.050 0.050 279.150 0.570 ;
   LAYER M3 ;
    RECT 279.050 0.050 279.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[29]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[30]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 291.850 0.050 291.950 0.570 ;
   LAYER M3 ;
    RECT 291.850 0.050 291.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[30]
 PIN D[31]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 295.850 0.050 295.950 0.570 ;
   LAYER M3 ;
    RECT 295.850 0.050 295.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[31]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 40.850 0.050 40.950 0.570 ;
   LAYER M3 ;
    RECT 40.850 0.050 40.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 45.050 0.050 45.150 0.570 ;
   LAYER M3 ;
    RECT 45.050 0.050 45.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 57.650 0.050 57.750 0.570 ;
   LAYER M3 ;
    RECT 57.650 0.050 57.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 61.850 0.050 61.950 0.570 ;
   LAYER M3 ;
    RECT 61.850 0.050 61.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN D[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 74.450 0.050 74.550 0.570 ;
   LAYER M3 ;
    RECT 74.450 0.050 74.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[8]
 PIN D[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 78.650 0.050 78.750 0.570 ;
   LAYER M3 ;
    RECT 78.650 0.050 78.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[9]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[10]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 89.850 0.050 89.950 0.570 ;
   LAYER M3 ;
    RECT 89.850 0.050 89.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[10]
 PIN Q[11]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 96.850 0.050 96.950 0.570 ;
   LAYER M3 ;
    RECT 96.850 0.050 96.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[11]
 PIN Q[12]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 106.650 0.050 106.750 0.570 ;
   LAYER M3 ;
    RECT 106.650 0.050 106.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[12]
 PIN Q[13]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 113.650 0.050 113.750 0.570 ;
   LAYER M3 ;
    RECT 113.650 0.050 113.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[13]
 PIN Q[14]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 123.450 0.050 123.550 0.570 ;
   LAYER M3 ;
    RECT 123.450 0.050 123.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[14]
 PIN Q[15]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 130.450 0.050 130.550 0.570 ;
   LAYER M3 ;
    RECT 130.450 0.050 130.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[15]
 PIN Q[16]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 172.850 0.050 172.950 0.570 ;
   LAYER M3 ;
    RECT 172.850 0.050 172.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[16]
 PIN Q[17]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 179.650 0.050 179.750 0.570 ;
   LAYER M3 ;
    RECT 179.650 0.050 179.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[17]
 PIN Q[18]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 189.650 0.050 189.750 0.570 ;
   LAYER M3 ;
    RECT 189.650 0.050 189.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[18]
 PIN Q[19]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 196.450 0.050 196.550 0.570 ;
   LAYER M3 ;
    RECT 196.450 0.050 196.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[19]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[20]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 206.450 0.050 206.550 0.570 ;
   LAYER M3 ;
    RECT 206.450 0.050 206.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[20]
 PIN Q[21]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 213.250 0.050 213.350 0.570 ;
   LAYER M3 ;
    RECT 213.250 0.050 213.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[21]
 PIN Q[22]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 223.250 0.050 223.350 0.570 ;
   LAYER M3 ;
    RECT 223.250 0.050 223.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[22]
 PIN Q[23]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 230.050 0.050 230.150 0.570 ;
   LAYER M3 ;
    RECT 230.050 0.050 230.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[23]
 PIN Q[24]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 240.050 0.050 240.150 0.570 ;
   LAYER M3 ;
    RECT 240.050 0.050 240.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[24]
 PIN Q[25]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 246.850 0.050 246.950 0.570 ;
   LAYER M3 ;
    RECT 246.850 0.050 246.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[25]
 PIN Q[26]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 256.850 0.050 256.950 0.570 ;
   LAYER M3 ;
    RECT 256.850 0.050 256.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[26]
 PIN Q[27]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 263.650 0.050 263.750 0.570 ;
   LAYER M3 ;
    RECT 263.650 0.050 263.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[27]
 PIN Q[28]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 273.650 0.050 273.750 0.570 ;
   LAYER M3 ;
    RECT 273.650 0.050 273.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[28]
 PIN Q[29]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 280.450 0.050 280.550 0.570 ;
   LAYER M3 ;
    RECT 280.450 0.050 280.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[29]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[30]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 290.450 0.050 290.550 0.570 ;
   LAYER M3 ;
    RECT 290.450 0.050 290.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[30]
 PIN Q[31]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 297.250 0.050 297.350 0.570 ;
   LAYER M3 ;
    RECT 297.250 0.050 297.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[31]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 39.450 0.050 39.550 0.570 ;
   LAYER M3 ;
    RECT 39.450 0.050 39.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 46.450 0.050 46.550 0.570 ;
   LAYER M3 ;
    RECT 46.450 0.050 46.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 56.250 0.050 56.350 0.570 ;
   LAYER M3 ;
    RECT 56.250 0.050 56.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 63.250 0.050 63.350 0.570 ;
   LAYER M3 ;
    RECT 63.250 0.050 63.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN Q[8]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 73.050 0.050 73.150 0.570 ;
   LAYER M3 ;
    RECT 73.050 0.050 73.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[8]
 PIN Q[9]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 80.050 0.050 80.150 0.570 ;
   LAYER M3 ;
    RECT 80.050 0.050 80.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[9]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 303.050 0.050 303.150 0.570 ;
   LAYER M3 ;
    RECT 303.050 0.050 303.150 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 161.250 0.050 161.350 0.570 ;
   LAYER M3 ;
    RECT 161.250 0.050 161.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 153.250 0.050 153.350 0.570 ;
   LAYER M3 ;
    RECT 153.250 0.050 153.350 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 0.495 1.725 303.920 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 303.920 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 303.920 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 303.920 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 303.920 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 303.920 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 303.920 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 303.920 23.605 ;
   LAYER M4 ;
    RECT 302.535 25.290 302.915 98.575 ;
   LAYER M4 ;
    RECT 301.495 25.290 302.195 98.575 ;
   LAYER M4 ;
    RECT 299.395 25.290 300.095 98.575 ;
   LAYER M4 ;
    RECT 297.295 25.290 297.995 98.575 ;
   LAYER M4 ;
    RECT 295.195 25.290 295.895 98.575 ;
   LAYER M4 ;
    RECT 293.095 25.290 293.795 98.575 ;
   LAYER M4 ;
    RECT 292.045 25.400 292.745 98.575 ;
   LAYER M4 ;
    RECT 290.995 25.290 291.695 98.575 ;
   LAYER M4 ;
    RECT 288.895 25.290 289.595 98.575 ;
   LAYER M4 ;
    RECT 286.795 25.290 287.495 98.575 ;
   LAYER M4 ;
    RECT 284.695 25.290 285.395 98.575 ;
   LAYER M4 ;
    RECT 282.595 25.290 283.295 98.575 ;
   LAYER M4 ;
    RECT 280.495 25.290 281.195 98.575 ;
   LAYER M4 ;
    RECT 278.395 25.290 279.095 98.575 ;
   LAYER M4 ;
    RECT 276.295 25.290 276.995 98.575 ;
   LAYER M4 ;
    RECT 275.245 25.400 275.945 98.575 ;
   LAYER M4 ;
    RECT 274.195 25.290 274.895 98.575 ;
   LAYER M4 ;
    RECT 272.095 25.290 272.795 98.575 ;
   LAYER M4 ;
    RECT 269.995 25.290 270.695 98.575 ;
   LAYER M4 ;
    RECT 267.895 25.290 268.595 98.575 ;
   LAYER M4 ;
    RECT 265.795 25.290 266.495 98.575 ;
   LAYER M4 ;
    RECT 263.695 25.290 264.395 98.575 ;
   LAYER M4 ;
    RECT 261.595 25.290 262.295 98.575 ;
   LAYER M4 ;
    RECT 259.495 25.290 260.195 98.575 ;
   LAYER M4 ;
    RECT 258.445 25.400 259.145 98.575 ;
   LAYER M4 ;
    RECT 257.395 25.290 258.095 98.575 ;
   LAYER M4 ;
    RECT 255.295 25.290 255.995 98.575 ;
   LAYER M4 ;
    RECT 253.195 25.290 253.895 98.575 ;
   LAYER M4 ;
    RECT 251.095 25.290 251.795 98.575 ;
   LAYER M4 ;
    RECT 248.995 25.290 249.695 98.575 ;
   LAYER M4 ;
    RECT 246.895 25.290 247.595 98.575 ;
   LAYER M4 ;
    RECT 244.795 25.290 245.495 98.575 ;
   LAYER M4 ;
    RECT 242.695 25.290 243.395 98.575 ;
   LAYER M4 ;
    RECT 241.645 25.400 242.345 98.575 ;
   LAYER M4 ;
    RECT 240.595 25.290 241.295 98.575 ;
   LAYER M4 ;
    RECT 238.495 25.290 239.195 98.575 ;
   LAYER M4 ;
    RECT 236.395 25.290 237.095 98.575 ;
   LAYER M4 ;
    RECT 234.295 25.290 234.995 98.575 ;
   LAYER M4 ;
    RECT 232.195 25.290 232.895 98.575 ;
   LAYER M4 ;
    RECT 230.095 25.290 230.795 98.575 ;
   LAYER M4 ;
    RECT 227.995 25.290 228.695 98.575 ;
   LAYER M4 ;
    RECT 225.895 25.290 226.595 98.575 ;
   LAYER M4 ;
    RECT 224.845 25.400 225.545 98.575 ;
   LAYER M4 ;
    RECT 223.795 25.290 224.495 98.575 ;
   LAYER M4 ;
    RECT 221.695 25.290 222.395 98.575 ;
   LAYER M4 ;
    RECT 219.595 25.290 220.295 98.575 ;
   LAYER M4 ;
    RECT 217.495 25.290 218.195 98.575 ;
   LAYER M4 ;
    RECT 215.395 25.290 216.095 98.575 ;
   LAYER M4 ;
    RECT 213.295 25.290 213.995 98.575 ;
   LAYER M4 ;
    RECT 211.195 25.290 211.895 98.575 ;
   LAYER M4 ;
    RECT 209.095 25.290 209.795 98.575 ;
   LAYER M4 ;
    RECT 208.045 25.400 208.745 98.575 ;
   LAYER M4 ;
    RECT 206.995 25.290 207.695 98.575 ;
   LAYER M4 ;
    RECT 204.895 25.290 205.595 98.575 ;
   LAYER M4 ;
    RECT 202.795 25.290 203.495 98.575 ;
   LAYER M4 ;
    RECT 200.695 25.290 201.395 98.575 ;
   LAYER M4 ;
    RECT 198.595 25.290 199.295 98.575 ;
   LAYER M4 ;
    RECT 196.495 25.290 197.195 98.575 ;
   LAYER M4 ;
    RECT 194.395 25.290 195.095 98.575 ;
   LAYER M4 ;
    RECT 192.295 25.290 192.995 98.575 ;
   LAYER M4 ;
    RECT 191.245 25.400 191.945 98.575 ;
   LAYER M4 ;
    RECT 190.195 25.290 190.895 98.575 ;
   LAYER M4 ;
    RECT 188.095 25.290 188.795 98.575 ;
   LAYER M4 ;
    RECT 185.995 25.290 186.695 98.575 ;
   LAYER M4 ;
    RECT 183.895 25.290 184.595 98.575 ;
   LAYER M4 ;
    RECT 181.795 25.290 182.495 98.575 ;
   LAYER M4 ;
    RECT 179.695 25.290 180.395 98.575 ;
   LAYER M4 ;
    RECT 177.595 25.290 178.295 98.575 ;
   LAYER M4 ;
    RECT 175.495 25.290 176.195 98.575 ;
   LAYER M4 ;
    RECT 174.445 25.400 175.145 98.575 ;
   LAYER M4 ;
    RECT 173.395 25.290 174.095 98.575 ;
   LAYER M4 ;
    RECT 171.295 25.290 171.995 98.575 ;
   LAYER M4 ;
    RECT 169.195 25.290 169.895 98.575 ;
   LAYER M4 ;
    RECT 167.095 25.360 167.795 98.575 ;
   LAYER M4 ;
    RECT 164.995 25.360 165.695 98.575 ;
   LAYER M4 ;
    RECT 163.310 25.360 163.690 98.575 ;
   LAYER M4 ;
    RECT 160.815 25.360 161.215 98.575 ;
   LAYER M4 ;
    RECT 159.345 25.360 159.845 98.575 ;
   LAYER M4 ;
    RECT 157.295 25.360 158.355 98.575 ;
   LAYER M4 ;
    RECT 154.390 25.360 154.790 98.575 ;
   LAYER M4 ;
    RECT 151.745 25.360 152.345 98.575 ;
   LAYER M4 ;
    RECT 150.075 25.360 150.720 98.575 ;
   LAYER M4 ;
    RECT 146.820 25.360 147.620 98.575 ;
   LAYER M4 ;
    RECT 145.825 25.360 146.225 98.575 ;
   LAYER M4 ;
    RECT 144.220 25.360 144.620 98.575 ;
   LAYER M4 ;
    RECT 142.005 25.360 142.810 98.575 ;
   LAYER M4 ;
    RECT 140.695 25.360 141.495 98.575 ;
   LAYER M4 ;
    RECT 138.275 25.360 138.895 98.575 ;
   LAYER M4 ;
    RECT 135.990 25.360 136.630 98.575 ;
   LAYER M4 ;
    RECT 134.555 25.290 135.255 98.575 ;
   LAYER M4 ;
    RECT 132.455 25.290 133.155 98.575 ;
   LAYER M4 ;
    RECT 130.355 25.290 131.055 98.575 ;
   LAYER M4 ;
    RECT 128.255 25.290 128.955 98.575 ;
   LAYER M4 ;
    RECT 126.155 25.290 126.855 98.575 ;
   LAYER M4 ;
    RECT 125.105 25.400 125.805 98.575 ;
   LAYER M4 ;
    RECT 124.055 25.290 124.755 98.575 ;
   LAYER M4 ;
    RECT 121.955 25.290 122.655 98.575 ;
   LAYER M4 ;
    RECT 119.855 25.290 120.555 98.575 ;
   LAYER M4 ;
    RECT 117.755 25.290 118.455 98.575 ;
   LAYER M4 ;
    RECT 115.655 25.290 116.355 98.575 ;
   LAYER M4 ;
    RECT 113.555 25.290 114.255 98.575 ;
   LAYER M4 ;
    RECT 111.455 25.290 112.155 98.575 ;
   LAYER M4 ;
    RECT 109.355 25.290 110.055 98.575 ;
   LAYER M4 ;
    RECT 108.305 25.400 109.005 98.575 ;
   LAYER M4 ;
    RECT 107.255 25.290 107.955 98.575 ;
   LAYER M4 ;
    RECT 105.155 25.290 105.855 98.575 ;
   LAYER M4 ;
    RECT 103.055 25.290 103.755 98.575 ;
   LAYER M4 ;
    RECT 100.955 25.290 101.655 98.575 ;
   LAYER M4 ;
    RECT 98.855 25.290 99.555 98.575 ;
   LAYER M4 ;
    RECT 96.755 25.290 97.455 98.575 ;
   LAYER M4 ;
    RECT 94.655 25.290 95.355 98.575 ;
   LAYER M4 ;
    RECT 92.555 25.290 93.255 98.575 ;
   LAYER M4 ;
    RECT 91.505 25.400 92.205 98.575 ;
   LAYER M4 ;
    RECT 90.455 25.290 91.155 98.575 ;
   LAYER M4 ;
    RECT 88.355 25.290 89.055 98.575 ;
   LAYER M4 ;
    RECT 86.255 25.290 86.955 98.575 ;
   LAYER M4 ;
    RECT 84.155 25.290 84.855 98.575 ;
   LAYER M4 ;
    RECT 82.055 25.290 82.755 98.575 ;
   LAYER M4 ;
    RECT 79.955 25.290 80.655 98.575 ;
   LAYER M4 ;
    RECT 77.855 25.290 78.555 98.575 ;
   LAYER M4 ;
    RECT 75.755 25.290 76.455 98.575 ;
   LAYER M4 ;
    RECT 74.705 25.400 75.405 98.575 ;
   LAYER M4 ;
    RECT 73.655 25.290 74.355 98.575 ;
   LAYER M4 ;
    RECT 71.555 25.290 72.255 98.575 ;
   LAYER M4 ;
    RECT 69.455 25.290 70.155 98.575 ;
   LAYER M4 ;
    RECT 67.355 25.290 68.055 98.575 ;
   LAYER M4 ;
    RECT 65.255 25.290 65.955 98.575 ;
   LAYER M4 ;
    RECT 63.155 25.290 63.855 98.575 ;
   LAYER M4 ;
    RECT 61.055 25.290 61.755 98.575 ;
   LAYER M4 ;
    RECT 58.955 25.290 59.655 98.575 ;
   LAYER M4 ;
    RECT 57.905 25.400 58.605 98.575 ;
   LAYER M4 ;
    RECT 56.855 25.290 57.555 98.575 ;
   LAYER M4 ;
    RECT 54.755 25.290 55.455 98.575 ;
   LAYER M4 ;
    RECT 52.655 25.290 53.355 98.575 ;
   LAYER M4 ;
    RECT 50.555 25.290 51.255 98.575 ;
   LAYER M4 ;
    RECT 48.455 25.290 49.155 98.575 ;
   LAYER M4 ;
    RECT 46.355 25.290 47.055 98.575 ;
   LAYER M4 ;
    RECT 44.255 25.290 44.955 98.575 ;
   LAYER M4 ;
    RECT 42.155 25.290 42.855 98.575 ;
   LAYER M4 ;
    RECT 41.105 25.400 41.805 98.575 ;
   LAYER M4 ;
    RECT 40.055 25.290 40.755 98.575 ;
   LAYER M4 ;
    RECT 37.955 25.290 38.655 98.575 ;
   LAYER M4 ;
    RECT 35.855 25.290 36.555 98.575 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 98.575 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 98.575 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 98.575 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 98.575 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 98.575 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 98.575 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 98.575 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 98.575 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 98.575 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 98.575 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 98.575 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 98.575 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 98.575 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 98.575 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 98.575 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 98.575 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 98.575 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 98.575 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 98.575 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 0.495 0.760 303.920 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 303.920 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 303.920 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 303.920 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 303.920 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 303.920 11.960 ;
   LAYER M4 ;
    RECT 0.495 14.840 303.920 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 303.920 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 303.920 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 303.920 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 303.920 25.115 ;
   LAYER M4 ;
    RECT 300.445 25.290 301.145 98.575 ;
   LAYER M4 ;
    RECT 298.345 25.290 299.045 98.575 ;
   LAYER M4 ;
    RECT 296.245 25.290 296.945 98.575 ;
   LAYER M4 ;
    RECT 294.145 25.400 294.845 98.575 ;
   LAYER M4 ;
    RECT 289.945 25.290 290.645 98.575 ;
   LAYER M4 ;
    RECT 287.845 25.290 288.545 98.575 ;
   LAYER M4 ;
    RECT 285.745 25.290 286.445 98.575 ;
   LAYER M4 ;
    RECT 283.645 25.290 284.345 98.575 ;
   LAYER M4 ;
    RECT 281.545 25.290 282.245 98.575 ;
   LAYER M4 ;
    RECT 279.445 25.290 280.145 98.575 ;
   LAYER M4 ;
    RECT 277.345 25.400 278.045 98.575 ;
   LAYER M4 ;
    RECT 273.145 25.290 273.845 98.575 ;
   LAYER M4 ;
    RECT 271.045 25.290 271.745 98.575 ;
   LAYER M4 ;
    RECT 268.945 25.290 269.645 98.575 ;
   LAYER M4 ;
    RECT 266.845 25.290 267.545 98.575 ;
   LAYER M4 ;
    RECT 264.745 25.290 265.445 98.575 ;
   LAYER M4 ;
    RECT 262.645 25.290 263.345 98.575 ;
   LAYER M4 ;
    RECT 260.545 25.400 261.245 98.575 ;
   LAYER M4 ;
    RECT 256.345 25.290 257.045 98.575 ;
   LAYER M4 ;
    RECT 254.245 25.290 254.945 98.575 ;
   LAYER M4 ;
    RECT 252.145 25.290 252.845 98.575 ;
   LAYER M4 ;
    RECT 250.045 25.290 250.745 98.575 ;
   LAYER M4 ;
    RECT 247.945 25.290 248.645 98.575 ;
   LAYER M4 ;
    RECT 245.845 25.290 246.545 98.575 ;
   LAYER M4 ;
    RECT 243.745 25.400 244.445 98.575 ;
   LAYER M4 ;
    RECT 239.545 25.290 240.245 98.575 ;
   LAYER M4 ;
    RECT 237.445 25.290 238.145 98.575 ;
   LAYER M4 ;
    RECT 235.345 25.290 236.045 98.575 ;
   LAYER M4 ;
    RECT 233.245 25.290 233.945 98.575 ;
   LAYER M4 ;
    RECT 231.145 25.290 231.845 98.575 ;
   LAYER M4 ;
    RECT 229.045 25.290 229.745 98.575 ;
   LAYER M4 ;
    RECT 226.945 25.400 227.645 98.575 ;
   LAYER M4 ;
    RECT 222.745 25.290 223.445 98.575 ;
   LAYER M4 ;
    RECT 220.645 25.290 221.345 98.575 ;
   LAYER M4 ;
    RECT 218.545 25.290 219.245 98.575 ;
   LAYER M4 ;
    RECT 216.445 25.290 217.145 98.575 ;
   LAYER M4 ;
    RECT 214.345 25.290 215.045 98.575 ;
   LAYER M4 ;
    RECT 212.245 25.290 212.945 98.575 ;
   LAYER M4 ;
    RECT 210.145 25.400 210.845 98.575 ;
   LAYER M4 ;
    RECT 205.945 25.290 206.645 98.575 ;
   LAYER M4 ;
    RECT 203.845 25.290 204.545 98.575 ;
   LAYER M4 ;
    RECT 201.745 25.290 202.445 98.575 ;
   LAYER M4 ;
    RECT 199.645 25.290 200.345 98.575 ;
   LAYER M4 ;
    RECT 197.545 25.290 198.245 98.575 ;
   LAYER M4 ;
    RECT 195.445 25.290 196.145 98.575 ;
   LAYER M4 ;
    RECT 193.345 25.400 194.045 98.575 ;
   LAYER M4 ;
    RECT 189.145 25.290 189.845 98.575 ;
   LAYER M4 ;
    RECT 187.045 25.290 187.745 98.575 ;
   LAYER M4 ;
    RECT 184.945 25.290 185.645 98.575 ;
   LAYER M4 ;
    RECT 182.845 25.290 183.545 98.575 ;
   LAYER M4 ;
    RECT 180.745 25.290 181.445 98.575 ;
   LAYER M4 ;
    RECT 178.645 25.290 179.345 98.575 ;
   LAYER M4 ;
    RECT 176.545 25.400 177.245 98.575 ;
   LAYER M4 ;
    RECT 172.345 25.290 173.045 98.575 ;
   LAYER M4 ;
    RECT 170.245 25.290 170.945 98.575 ;
   LAYER M4 ;
    RECT 168.145 25.290 168.845 98.575 ;
   LAYER M4 ;
    RECT 166.045 25.360 166.745 98.575 ;
   LAYER M4 ;
    RECT 163.945 25.360 164.645 98.575 ;
   LAYER M4 ;
    RECT 162.735 25.360 163.115 98.575 ;
   LAYER M4 ;
    RECT 161.530 25.360 162.510 98.575 ;
   LAYER M4 ;
    RECT 160.100 25.360 160.500 98.575 ;
   LAYER M4 ;
    RECT 158.605 25.360 159.105 98.575 ;
   LAYER M4 ;
    RECT 155.745 25.360 156.805 98.575 ;
   LAYER M4 ;
    RECT 155.065 25.360 155.465 98.575 ;
   LAYER M4 ;
    RECT 153.050 25.360 154.110 98.575 ;
   LAYER M4 ;
    RECT 151.035 25.360 151.435 98.575 ;
   LAYER M4 ;
    RECT 148.370 25.360 149.325 98.575 ;
   LAYER M4 ;
    RECT 144.910 25.360 145.550 98.575 ;
   LAYER M4 ;
    RECT 143.310 25.360 143.900 98.575 ;
   LAYER M4 ;
    RECT 139.395 25.360 140.195 98.575 ;
   LAYER M4 ;
    RECT 137.130 25.360 137.770 98.575 ;
   LAYER M4 ;
    RECT 133.505 25.290 134.205 98.575 ;
   LAYER M4 ;
    RECT 131.405 25.290 132.105 98.575 ;
   LAYER M4 ;
    RECT 129.305 25.290 130.005 98.575 ;
   LAYER M4 ;
    RECT 127.205 25.400 127.905 98.575 ;
   LAYER M4 ;
    RECT 123.005 25.290 123.705 98.575 ;
   LAYER M4 ;
    RECT 120.905 25.290 121.605 98.575 ;
   LAYER M4 ;
    RECT 118.805 25.290 119.505 98.575 ;
   LAYER M4 ;
    RECT 116.705 25.290 117.405 98.575 ;
   LAYER M4 ;
    RECT 114.605 25.290 115.305 98.575 ;
   LAYER M4 ;
    RECT 112.505 25.290 113.205 98.575 ;
   LAYER M4 ;
    RECT 110.405 25.400 111.105 98.575 ;
   LAYER M4 ;
    RECT 106.205 25.290 106.905 98.575 ;
   LAYER M4 ;
    RECT 104.105 25.290 104.805 98.575 ;
   LAYER M4 ;
    RECT 102.005 25.290 102.705 98.575 ;
   LAYER M4 ;
    RECT 99.905 25.290 100.605 98.575 ;
   LAYER M4 ;
    RECT 97.805 25.290 98.505 98.575 ;
   LAYER M4 ;
    RECT 95.705 25.290 96.405 98.575 ;
   LAYER M4 ;
    RECT 93.605 25.400 94.305 98.575 ;
   LAYER M4 ;
    RECT 89.405 25.290 90.105 98.575 ;
   LAYER M4 ;
    RECT 87.305 25.290 88.005 98.575 ;
   LAYER M4 ;
    RECT 85.205 25.290 85.905 98.575 ;
   LAYER M4 ;
    RECT 83.105 25.290 83.805 98.575 ;
   LAYER M4 ;
    RECT 81.005 25.290 81.705 98.575 ;
   LAYER M4 ;
    RECT 78.905 25.290 79.605 98.575 ;
   LAYER M4 ;
    RECT 76.805 25.400 77.505 98.575 ;
   LAYER M4 ;
    RECT 72.605 25.290 73.305 98.575 ;
   LAYER M4 ;
    RECT 70.505 25.290 71.205 98.575 ;
   LAYER M4 ;
    RECT 68.405 25.290 69.105 98.575 ;
   LAYER M4 ;
    RECT 66.305 25.290 67.005 98.575 ;
   LAYER M4 ;
    RECT 64.205 25.290 64.905 98.575 ;
   LAYER M4 ;
    RECT 62.105 25.290 62.805 98.575 ;
   LAYER M4 ;
    RECT 60.005 25.400 60.705 98.575 ;
   LAYER M4 ;
    RECT 55.805 25.290 56.505 98.575 ;
   LAYER M4 ;
    RECT 53.705 25.290 54.405 98.575 ;
   LAYER M4 ;
    RECT 51.605 25.290 52.305 98.575 ;
   LAYER M4 ;
    RECT 49.505 25.290 50.205 98.575 ;
   LAYER M4 ;
    RECT 47.405 25.290 48.105 98.575 ;
   LAYER M4 ;
    RECT 45.305 25.290 46.005 98.575 ;
   LAYER M4 ;
    RECT 43.205 25.400 43.905 98.575 ;
   LAYER M4 ;
    RECT 39.005 25.290 39.705 98.575 ;
   LAYER M4 ;
    RECT 36.905 25.290 37.605 98.575 ;
   LAYER M4 ;
    RECT 34.805 25.290 35.505 98.575 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 98.575 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 98.575 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 98.575 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 98.575 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 98.575 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 98.575 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 98.575 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 98.575 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 98.575 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 98.575 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 98.575 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 98.575 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 98.575 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 98.575 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 304.750 99.350 ;
  LAYER M2 ;
   RECT 0.050 0.050 304.750 99.350 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 39.450 0.050 39.550 0.570 ;
  LAYER VIA2 ;
   RECT 40.850 0.050 40.950 0.570 ;
  LAYER VIA2 ;
   RECT 45.050 0.050 45.150 0.570 ;
  LAYER VIA2 ;
   RECT 46.450 0.050 46.550 0.570 ;
  LAYER VIA2 ;
   RECT 56.250 0.050 56.350 0.570 ;
  LAYER VIA2 ;
   RECT 57.650 0.050 57.750 0.570 ;
  LAYER VIA2 ;
   RECT 61.850 0.050 61.950 0.570 ;
  LAYER VIA2 ;
   RECT 63.250 0.050 63.350 0.570 ;
  LAYER VIA2 ;
   RECT 73.050 0.050 73.150 0.570 ;
  LAYER VIA2 ;
   RECT 74.450 0.050 74.550 0.570 ;
  LAYER VIA2 ;
   RECT 78.650 0.050 78.750 0.570 ;
  LAYER VIA2 ;
   RECT 80.050 0.050 80.150 0.570 ;
  LAYER VIA2 ;
   RECT 89.850 0.050 89.950 0.570 ;
  LAYER VIA2 ;
   RECT 91.250 0.050 91.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.450 0.050 95.550 0.570 ;
  LAYER VIA2 ;
   RECT 96.850 0.050 96.950 0.570 ;
  LAYER VIA2 ;
   RECT 106.650 0.050 106.750 0.570 ;
  LAYER VIA2 ;
   RECT 108.050 0.050 108.150 0.570 ;
  LAYER VIA2 ;
   RECT 112.250 0.050 112.350 0.570 ;
  LAYER VIA2 ;
   RECT 113.650 0.050 113.750 0.570 ;
  LAYER VIA2 ;
   RECT 123.450 0.050 123.550 0.570 ;
  LAYER VIA2 ;
   RECT 124.850 0.050 124.950 0.570 ;
  LAYER VIA2 ;
   RECT 129.050 0.050 129.150 0.570 ;
  LAYER VIA2 ;
   RECT 130.450 0.050 130.550 0.570 ;
  LAYER VIA2 ;
   RECT 137.450 0.050 137.550 0.570 ;
  LAYER VIA2 ;
   RECT 146.050 0.050 146.150 0.570 ;
  LAYER VIA2 ;
   RECT 147.450 0.050 147.550 0.570 ;
  LAYER VIA2 ;
   RECT 148.250 0.050 148.350 0.570 ;
  LAYER VIA2 ;
   RECT 148.850 0.050 148.950 0.570 ;
  LAYER VIA2 ;
   RECT 149.450 0.050 149.550 0.570 ;
  LAYER VIA2 ;
   RECT 150.250 0.050 150.350 0.570 ;
  LAYER VIA2 ;
   RECT 151.850 0.050 151.950 0.570 ;
  LAYER VIA2 ;
   RECT 153.250 0.050 153.350 0.570 ;
  LAYER VIA2 ;
   RECT 155.850 0.050 155.950 0.570 ;
  LAYER VIA2 ;
   RECT 156.450 0.050 156.550 0.570 ;
  LAYER VIA2 ;
   RECT 160.650 0.050 160.750 0.570 ;
  LAYER VIA2 ;
   RECT 161.250 0.050 161.350 0.570 ;
  LAYER VIA2 ;
   RECT 162.050 0.050 162.150 0.570 ;
  LAYER VIA2 ;
   RECT 172.850 0.050 172.950 0.570 ;
  LAYER VIA2 ;
   RECT 174.250 0.050 174.350 0.570 ;
  LAYER VIA2 ;
   RECT 178.250 0.050 178.350 0.570 ;
  LAYER VIA2 ;
   RECT 179.650 0.050 179.750 0.570 ;
  LAYER VIA2 ;
   RECT 189.650 0.050 189.750 0.570 ;
  LAYER VIA2 ;
   RECT 191.050 0.050 191.150 0.570 ;
  LAYER VIA2 ;
   RECT 195.050 0.050 195.150 0.570 ;
  LAYER VIA2 ;
   RECT 196.450 0.050 196.550 0.570 ;
  LAYER VIA2 ;
   RECT 206.450 0.050 206.550 0.570 ;
  LAYER VIA2 ;
   RECT 207.850 0.050 207.950 0.570 ;
  LAYER VIA2 ;
   RECT 211.850 0.050 211.950 0.570 ;
  LAYER VIA2 ;
   RECT 213.250 0.050 213.350 0.570 ;
  LAYER VIA2 ;
   RECT 223.250 0.050 223.350 0.570 ;
  LAYER VIA2 ;
   RECT 224.650 0.050 224.750 0.570 ;
  LAYER VIA2 ;
   RECT 228.650 0.050 228.750 0.570 ;
  LAYER VIA2 ;
   RECT 230.050 0.050 230.150 0.570 ;
  LAYER VIA2 ;
   RECT 240.050 0.050 240.150 0.570 ;
  LAYER VIA2 ;
   RECT 241.450 0.050 241.550 0.570 ;
  LAYER VIA2 ;
   RECT 245.450 0.050 245.550 0.570 ;
  LAYER VIA2 ;
   RECT 246.850 0.050 246.950 0.570 ;
  LAYER VIA2 ;
   RECT 256.850 0.050 256.950 0.570 ;
  LAYER VIA2 ;
   RECT 258.250 0.050 258.350 0.570 ;
  LAYER VIA2 ;
   RECT 262.250 0.050 262.350 0.570 ;
  LAYER VIA2 ;
   RECT 263.650 0.050 263.750 0.570 ;
  LAYER VIA2 ;
   RECT 273.650 0.050 273.750 0.570 ;
  LAYER VIA2 ;
   RECT 275.050 0.050 275.150 0.570 ;
  LAYER VIA2 ;
   RECT 279.050 0.050 279.150 0.570 ;
  LAYER VIA2 ;
   RECT 280.450 0.050 280.550 0.570 ;
  LAYER VIA2 ;
   RECT 290.450 0.050 290.550 0.570 ;
  LAYER VIA2 ;
   RECT 291.850 0.050 291.950 0.570 ;
  LAYER VIA2 ;
   RECT 295.850 0.050 295.950 0.570 ;
  LAYER VIA2 ;
   RECT 297.250 0.050 297.350 0.570 ;
  LAYER VIA2 ;
   RECT 303.050 0.050 303.150 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 304.750 99.350 ;
  LAYER M4 ;
   RECT 0.050 0.050 304.750 99.350 ;
 END
END ST_SPHDL_1024x32m8_L

MACRO ST_SPHDL_1024x40m8_L
 CLASS BLOCK ;
   SIZE 372.000 BY 99.400 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 181.850 0.050 181.950 0.570 ;
   LAYER M3 ;
    RECT 181.850 0.050 181.950 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 182.450 0.050 182.550 0.570 ;
   LAYER M3 ;
    RECT 182.450 0.050 182.550 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 183.050 0.050 183.150 0.570 ;
   LAYER M3 ;
    RECT 183.050 0.050 183.150 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 189.450 0.050 189.550 0.570 ;
   LAYER M3 ;
    RECT 189.450 0.050 189.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 190.050 0.050 190.150 0.570 ;
   LAYER M3 ;
    RECT 190.050 0.050 190.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 183.850 0.050 183.950 0.570 ;
   LAYER M3 ;
    RECT 183.850 0.050 183.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 185.450 0.050 185.550 0.570 ;
   LAYER M3 ;
    RECT 185.450 0.050 185.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN A[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 179.650 0.050 179.750 0.570 ;
   LAYER M3 ;
    RECT 179.650 0.050 179.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.916 LAYER M2 ;
  ANTENNAMAXAREACAR 13.057 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.347 LAYER M3 ;
 END A[7]
 PIN A[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 181.050 0.050 181.150 0.570 ;
   LAYER M3 ;
    RECT 181.050 0.050 181.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.924 LAYER M2 ;
  ANTENNAMAXAREACAR 13.892 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.282 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.376 LAYER M3 ;
 END A[8]
 PIN A[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 171.050 0.050 171.150 0.570 ;
   LAYER M3 ;
    RECT 171.050 0.050 171.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.251 LAYER M2 ;
  ANTENNAGATEAREA 0.251 LAYER M3 ;
  ANTENNAMAXAREACAR 3.203 LAYER M2 ;
  ANTENNAMAXAREACAR 9.213 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.586 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.511 LAYER M3 ;
 END A[9]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 194.250 0.050 194.350 0.570 ;
   LAYER M3 ;
    RECT 194.250 0.050 194.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 195.650 0.050 195.750 0.570 ;
   LAYER M3 ;
    RECT 195.650 0.050 195.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 91.250 0.050 91.350 0.570 ;
   LAYER M3 ;
    RECT 91.250 0.050 91.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[10]
 PIN D[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 95.450 0.050 95.550 0.570 ;
   LAYER M3 ;
    RECT 95.450 0.050 95.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[11]
 PIN D[12]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 108.050 0.050 108.150 0.570 ;
   LAYER M3 ;
    RECT 108.050 0.050 108.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[12]
 PIN D[13]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 112.250 0.050 112.350 0.570 ;
   LAYER M3 ;
    RECT 112.250 0.050 112.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[13]
 PIN D[14]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 124.850 0.050 124.950 0.570 ;
   LAYER M3 ;
    RECT 124.850 0.050 124.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[14]
 PIN D[15]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 129.050 0.050 129.150 0.570 ;
   LAYER M3 ;
    RECT 129.050 0.050 129.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[15]
 PIN D[16]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 141.650 0.050 141.750 0.570 ;
   LAYER M3 ;
    RECT 141.650 0.050 141.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[16]
 PIN D[17]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 145.850 0.050 145.950 0.570 ;
   LAYER M3 ;
    RECT 145.850 0.050 145.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[17]
 PIN D[18]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 158.450 0.050 158.550 0.570 ;
   LAYER M3 ;
    RECT 158.450 0.050 158.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[18]
 PIN D[19]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 162.650 0.050 162.750 0.570 ;
   LAYER M3 ;
    RECT 162.650 0.050 162.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[19]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[20]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 207.850 0.050 207.950 0.570 ;
   LAYER M3 ;
    RECT 207.850 0.050 207.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[20]
 PIN D[21]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 211.850 0.050 211.950 0.570 ;
   LAYER M3 ;
    RECT 211.850 0.050 211.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[21]
 PIN D[22]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 224.650 0.050 224.750 0.570 ;
   LAYER M3 ;
    RECT 224.650 0.050 224.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[22]
 PIN D[23]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 228.650 0.050 228.750 0.570 ;
   LAYER M3 ;
    RECT 228.650 0.050 228.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[23]
 PIN D[24]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 241.450 0.050 241.550 0.570 ;
   LAYER M3 ;
    RECT 241.450 0.050 241.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[24]
 PIN D[25]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 245.450 0.050 245.550 0.570 ;
   LAYER M3 ;
    RECT 245.450 0.050 245.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[25]
 PIN D[26]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 258.250 0.050 258.350 0.570 ;
   LAYER M3 ;
    RECT 258.250 0.050 258.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[26]
 PIN D[27]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 262.250 0.050 262.350 0.570 ;
   LAYER M3 ;
    RECT 262.250 0.050 262.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[27]
 PIN D[28]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 275.050 0.050 275.150 0.570 ;
   LAYER M3 ;
    RECT 275.050 0.050 275.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[28]
 PIN D[29]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 279.050 0.050 279.150 0.570 ;
   LAYER M3 ;
    RECT 279.050 0.050 279.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[29]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[30]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 291.850 0.050 291.950 0.570 ;
   LAYER M3 ;
    RECT 291.850 0.050 291.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[30]
 PIN D[31]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 295.850 0.050 295.950 0.570 ;
   LAYER M3 ;
    RECT 295.850 0.050 295.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[31]
 PIN D[32]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 308.650 0.050 308.750 0.570 ;
   LAYER M3 ;
    RECT 308.650 0.050 308.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[32]
 PIN D[33]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 312.650 0.050 312.750 0.570 ;
   LAYER M3 ;
    RECT 312.650 0.050 312.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[33]
 PIN D[34]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 325.450 0.050 325.550 0.570 ;
   LAYER M3 ;
    RECT 325.450 0.050 325.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[34]
 PIN D[35]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 329.450 0.050 329.550 0.570 ;
   LAYER M3 ;
    RECT 329.450 0.050 329.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[35]
 PIN D[36]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 342.250 0.050 342.350 0.570 ;
   LAYER M3 ;
    RECT 342.250 0.050 342.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[36]
 PIN D[37]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 346.250 0.050 346.350 0.570 ;
   LAYER M3 ;
    RECT 346.250 0.050 346.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[37]
 PIN D[38]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 359.050 0.050 359.150 0.570 ;
   LAYER M3 ;
    RECT 359.050 0.050 359.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[38]
 PIN D[39]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 363.050 0.050 363.150 0.570 ;
   LAYER M3 ;
    RECT 363.050 0.050 363.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[39]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 40.850 0.050 40.950 0.570 ;
   LAYER M3 ;
    RECT 40.850 0.050 40.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 45.050 0.050 45.150 0.570 ;
   LAYER M3 ;
    RECT 45.050 0.050 45.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 57.650 0.050 57.750 0.570 ;
   LAYER M3 ;
    RECT 57.650 0.050 57.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 61.850 0.050 61.950 0.570 ;
   LAYER M3 ;
    RECT 61.850 0.050 61.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN D[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 74.450 0.050 74.550 0.570 ;
   LAYER M3 ;
    RECT 74.450 0.050 74.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[8]
 PIN D[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 78.650 0.050 78.750 0.570 ;
   LAYER M3 ;
    RECT 78.650 0.050 78.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[9]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[10]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 89.850 0.050 89.950 0.570 ;
   LAYER M3 ;
    RECT 89.850 0.050 89.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[10]
 PIN Q[11]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 96.850 0.050 96.950 0.570 ;
   LAYER M3 ;
    RECT 96.850 0.050 96.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[11]
 PIN Q[12]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 106.650 0.050 106.750 0.570 ;
   LAYER M3 ;
    RECT 106.650 0.050 106.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[12]
 PIN Q[13]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 113.650 0.050 113.750 0.570 ;
   LAYER M3 ;
    RECT 113.650 0.050 113.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[13]
 PIN Q[14]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 123.450 0.050 123.550 0.570 ;
   LAYER M3 ;
    RECT 123.450 0.050 123.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[14]
 PIN Q[15]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 130.450 0.050 130.550 0.570 ;
   LAYER M3 ;
    RECT 130.450 0.050 130.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[15]
 PIN Q[16]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 140.250 0.050 140.350 0.570 ;
   LAYER M3 ;
    RECT 140.250 0.050 140.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[16]
 PIN Q[17]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 147.250 0.050 147.350 0.570 ;
   LAYER M3 ;
    RECT 147.250 0.050 147.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[17]
 PIN Q[18]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 157.050 0.050 157.150 0.570 ;
   LAYER M3 ;
    RECT 157.050 0.050 157.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[18]
 PIN Q[19]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 164.050 0.050 164.150 0.570 ;
   LAYER M3 ;
    RECT 164.050 0.050 164.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[19]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[20]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 206.450 0.050 206.550 0.570 ;
   LAYER M3 ;
    RECT 206.450 0.050 206.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[20]
 PIN Q[21]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 213.250 0.050 213.350 0.570 ;
   LAYER M3 ;
    RECT 213.250 0.050 213.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[21]
 PIN Q[22]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 223.250 0.050 223.350 0.570 ;
   LAYER M3 ;
    RECT 223.250 0.050 223.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[22]
 PIN Q[23]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 230.050 0.050 230.150 0.570 ;
   LAYER M3 ;
    RECT 230.050 0.050 230.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[23]
 PIN Q[24]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 240.050 0.050 240.150 0.570 ;
   LAYER M3 ;
    RECT 240.050 0.050 240.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[24]
 PIN Q[25]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 246.850 0.050 246.950 0.570 ;
   LAYER M3 ;
    RECT 246.850 0.050 246.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[25]
 PIN Q[26]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 256.850 0.050 256.950 0.570 ;
   LAYER M3 ;
    RECT 256.850 0.050 256.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[26]
 PIN Q[27]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 263.650 0.050 263.750 0.570 ;
   LAYER M3 ;
    RECT 263.650 0.050 263.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[27]
 PIN Q[28]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 273.650 0.050 273.750 0.570 ;
   LAYER M3 ;
    RECT 273.650 0.050 273.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[28]
 PIN Q[29]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 280.450 0.050 280.550 0.570 ;
   LAYER M3 ;
    RECT 280.450 0.050 280.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[29]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[30]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 290.450 0.050 290.550 0.570 ;
   LAYER M3 ;
    RECT 290.450 0.050 290.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[30]
 PIN Q[31]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 297.250 0.050 297.350 0.570 ;
   LAYER M3 ;
    RECT 297.250 0.050 297.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[31]
 PIN Q[32]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 307.250 0.050 307.350 0.570 ;
   LAYER M3 ;
    RECT 307.250 0.050 307.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[32]
 PIN Q[33]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 314.050 0.050 314.150 0.570 ;
   LAYER M3 ;
    RECT 314.050 0.050 314.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[33]
 PIN Q[34]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 324.050 0.050 324.150 0.570 ;
   LAYER M3 ;
    RECT 324.050 0.050 324.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[34]
 PIN Q[35]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 330.850 0.050 330.950 0.570 ;
   LAYER M3 ;
    RECT 330.850 0.050 330.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[35]
 PIN Q[36]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 340.850 0.050 340.950 0.570 ;
   LAYER M3 ;
    RECT 340.850 0.050 340.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[36]
 PIN Q[37]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 347.650 0.050 347.750 0.570 ;
   LAYER M3 ;
    RECT 347.650 0.050 347.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[37]
 PIN Q[38]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 357.650 0.050 357.750 0.570 ;
   LAYER M3 ;
    RECT 357.650 0.050 357.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[38]
 PIN Q[39]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 364.450 0.050 364.550 0.570 ;
   LAYER M3 ;
    RECT 364.450 0.050 364.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[39]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 39.450 0.050 39.550 0.570 ;
   LAYER M3 ;
    RECT 39.450 0.050 39.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 46.450 0.050 46.550 0.570 ;
   LAYER M3 ;
    RECT 46.450 0.050 46.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 56.250 0.050 56.350 0.570 ;
   LAYER M3 ;
    RECT 56.250 0.050 56.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 63.250 0.050 63.350 0.570 ;
   LAYER M3 ;
    RECT 63.250 0.050 63.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN Q[8]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 73.050 0.050 73.150 0.570 ;
   LAYER M3 ;
    RECT 73.050 0.050 73.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[8]
 PIN Q[9]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 80.050 0.050 80.150 0.570 ;
   LAYER M3 ;
    RECT 80.050 0.050 80.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[9]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 370.250 0.050 370.350 0.570 ;
   LAYER M3 ;
    RECT 370.250 0.050 370.350 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 194.850 0.050 194.950 0.570 ;
   LAYER M3 ;
    RECT 194.850 0.050 194.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 186.850 0.050 186.950 0.570 ;
   LAYER M3 ;
    RECT 186.850 0.050 186.950 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 75.755 25.290 76.455 98.575 ;
   LAYER M4 ;
    RECT 74.705 25.400 75.405 98.575 ;
   LAYER M4 ;
    RECT 73.655 25.290 74.355 98.575 ;
   LAYER M4 ;
    RECT 71.555 25.290 72.255 98.575 ;
   LAYER M4 ;
    RECT 69.455 25.290 70.155 98.575 ;
   LAYER M4 ;
    RECT 67.355 25.290 68.055 98.575 ;
   LAYER M4 ;
    RECT 65.255 25.290 65.955 98.575 ;
   LAYER M4 ;
    RECT 63.155 25.290 63.855 98.575 ;
   LAYER M4 ;
    RECT 61.055 25.290 61.755 98.575 ;
   LAYER M4 ;
    RECT 58.955 25.290 59.655 98.575 ;
   LAYER M4 ;
    RECT 57.905 25.400 58.605 98.575 ;
   LAYER M4 ;
    RECT 56.855 25.290 57.555 98.575 ;
   LAYER M4 ;
    RECT 54.755 25.290 55.455 98.575 ;
   LAYER M4 ;
    RECT 52.655 25.290 53.355 98.575 ;
   LAYER M4 ;
    RECT 50.555 25.290 51.255 98.575 ;
   LAYER M4 ;
    RECT 48.455 25.290 49.155 98.575 ;
   LAYER M4 ;
    RECT 46.355 25.290 47.055 98.575 ;
   LAYER M4 ;
    RECT 44.255 25.290 44.955 98.575 ;
   LAYER M4 ;
    RECT 42.155 25.290 42.855 98.575 ;
   LAYER M4 ;
    RECT 41.105 25.400 41.805 98.575 ;
   LAYER M4 ;
    RECT 40.055 25.290 40.755 98.575 ;
   LAYER M4 ;
    RECT 37.955 25.290 38.655 98.575 ;
   LAYER M4 ;
    RECT 35.855 25.290 36.555 98.575 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 98.575 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 98.575 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 98.575 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 98.575 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 98.575 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 98.575 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 98.575 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 98.575 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 98.575 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 98.575 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 98.575 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 98.575 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 98.575 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 98.575 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 98.575 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 98.575 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 98.575 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 98.575 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 98.575 ;
   LAYER M4 ;
    RECT 295.195 25.290 295.895 98.575 ;
   LAYER M4 ;
    RECT 293.095 25.290 293.795 98.575 ;
   LAYER M4 ;
    RECT 292.045 25.400 292.745 98.575 ;
   LAYER M4 ;
    RECT 290.995 25.290 291.695 98.575 ;
   LAYER M4 ;
    RECT 288.895 25.290 289.595 98.575 ;
   LAYER M4 ;
    RECT 286.795 25.290 287.495 98.575 ;
   LAYER M4 ;
    RECT 284.695 25.290 285.395 98.575 ;
   LAYER M4 ;
    RECT 282.595 25.290 283.295 98.575 ;
   LAYER M4 ;
    RECT 280.495 25.290 281.195 98.575 ;
   LAYER M4 ;
    RECT 278.395 25.290 279.095 98.575 ;
   LAYER M4 ;
    RECT 276.295 25.290 276.995 98.575 ;
   LAYER M4 ;
    RECT 275.245 25.400 275.945 98.575 ;
   LAYER M4 ;
    RECT 274.195 25.290 274.895 98.575 ;
   LAYER M4 ;
    RECT 272.095 25.290 272.795 98.575 ;
   LAYER M4 ;
    RECT 269.995 25.290 270.695 98.575 ;
   LAYER M4 ;
    RECT 267.895 25.290 268.595 98.575 ;
   LAYER M4 ;
    RECT 265.795 25.290 266.495 98.575 ;
   LAYER M4 ;
    RECT 263.695 25.290 264.395 98.575 ;
   LAYER M4 ;
    RECT 261.595 25.290 262.295 98.575 ;
   LAYER M4 ;
    RECT 259.495 25.290 260.195 98.575 ;
   LAYER M4 ;
    RECT 258.445 25.400 259.145 98.575 ;
   LAYER M4 ;
    RECT 257.395 25.290 258.095 98.575 ;
   LAYER M4 ;
    RECT 255.295 25.290 255.995 98.575 ;
   LAYER M4 ;
    RECT 253.195 25.290 253.895 98.575 ;
   LAYER M4 ;
    RECT 251.095 25.290 251.795 98.575 ;
   LAYER M4 ;
    RECT 248.995 25.290 249.695 98.575 ;
   LAYER M4 ;
    RECT 246.895 25.290 247.595 98.575 ;
   LAYER M4 ;
    RECT 244.795 25.290 245.495 98.575 ;
   LAYER M4 ;
    RECT 242.695 25.290 243.395 98.575 ;
   LAYER M4 ;
    RECT 241.645 25.400 242.345 98.575 ;
   LAYER M4 ;
    RECT 240.595 25.290 241.295 98.575 ;
   LAYER M4 ;
    RECT 238.495 25.290 239.195 98.575 ;
   LAYER M4 ;
    RECT 236.395 25.290 237.095 98.575 ;
   LAYER M4 ;
    RECT 234.295 25.290 234.995 98.575 ;
   LAYER M4 ;
    RECT 232.195 25.290 232.895 98.575 ;
   LAYER M4 ;
    RECT 230.095 25.290 230.795 98.575 ;
   LAYER M4 ;
    RECT 227.995 25.290 228.695 98.575 ;
   LAYER M4 ;
    RECT 225.895 25.290 226.595 98.575 ;
   LAYER M4 ;
    RECT 224.845 25.400 225.545 98.575 ;
   LAYER M4 ;
    RECT 223.795 25.290 224.495 98.575 ;
   LAYER M4 ;
    RECT 221.695 25.290 222.395 98.575 ;
   LAYER M4 ;
    RECT 219.595 25.290 220.295 98.575 ;
   LAYER M4 ;
    RECT 217.495 25.290 218.195 98.575 ;
   LAYER M4 ;
    RECT 215.395 25.290 216.095 98.575 ;
   LAYER M4 ;
    RECT 213.295 25.290 213.995 98.575 ;
   LAYER M4 ;
    RECT 211.195 25.290 211.895 98.575 ;
   LAYER M4 ;
    RECT 209.095 25.290 209.795 98.575 ;
   LAYER M4 ;
    RECT 208.045 25.400 208.745 98.575 ;
   LAYER M4 ;
    RECT 206.995 25.290 207.695 98.575 ;
   LAYER M4 ;
    RECT 204.895 25.290 205.595 98.575 ;
   LAYER M4 ;
    RECT 202.795 25.290 203.495 98.575 ;
   LAYER M4 ;
    RECT 200.695 25.360 201.395 98.575 ;
   LAYER M4 ;
    RECT 198.595 25.360 199.295 98.575 ;
   LAYER M4 ;
    RECT 196.910 25.360 197.290 98.575 ;
   LAYER M4 ;
    RECT 194.415 25.360 194.815 98.575 ;
   LAYER M4 ;
    RECT 192.945 25.360 193.445 98.575 ;
   LAYER M4 ;
    RECT 190.895 25.360 191.955 98.575 ;
   LAYER M4 ;
    RECT 187.990 25.360 188.390 98.575 ;
   LAYER M4 ;
    RECT 185.345 25.360 185.945 98.575 ;
   LAYER M4 ;
    RECT 183.675 25.360 184.320 98.575 ;
   LAYER M4 ;
    RECT 180.420 25.360 181.220 98.575 ;
   LAYER M4 ;
    RECT 179.425 25.360 179.825 98.575 ;
   LAYER M4 ;
    RECT 177.820 25.360 178.220 98.575 ;
   LAYER M4 ;
    RECT 175.605 25.360 176.410 98.575 ;
   LAYER M4 ;
    RECT 174.295 25.360 175.095 98.575 ;
   LAYER M4 ;
    RECT 171.875 25.360 172.495 98.575 ;
   LAYER M4 ;
    RECT 169.590 25.360 170.230 98.575 ;
   LAYER M4 ;
    RECT 168.155 25.290 168.855 98.575 ;
   LAYER M4 ;
    RECT 166.055 25.290 166.755 98.575 ;
   LAYER M4 ;
    RECT 163.955 25.290 164.655 98.575 ;
   LAYER M4 ;
    RECT 161.855 25.290 162.555 98.575 ;
   LAYER M4 ;
    RECT 159.755 25.290 160.455 98.575 ;
   LAYER M4 ;
    RECT 158.705 25.400 159.405 98.575 ;
   LAYER M4 ;
    RECT 157.655 25.290 158.355 98.575 ;
   LAYER M4 ;
    RECT 155.555 25.290 156.255 98.575 ;
   LAYER M4 ;
    RECT 153.455 25.290 154.155 98.575 ;
   LAYER M4 ;
    RECT 151.355 25.290 152.055 98.575 ;
   LAYER M4 ;
    RECT 149.255 25.290 149.955 98.575 ;
   LAYER M4 ;
    RECT 147.155 25.290 147.855 98.575 ;
   LAYER M4 ;
    RECT 145.055 25.290 145.755 98.575 ;
   LAYER M4 ;
    RECT 142.955 25.290 143.655 98.575 ;
   LAYER M4 ;
    RECT 141.905 25.400 142.605 98.575 ;
   LAYER M4 ;
    RECT 140.855 25.290 141.555 98.575 ;
   LAYER M4 ;
    RECT 138.755 25.290 139.455 98.575 ;
   LAYER M4 ;
    RECT 136.655 25.290 137.355 98.575 ;
   LAYER M4 ;
    RECT 134.555 25.290 135.255 98.575 ;
   LAYER M4 ;
    RECT 132.455 25.290 133.155 98.575 ;
   LAYER M4 ;
    RECT 130.355 25.290 131.055 98.575 ;
   LAYER M4 ;
    RECT 128.255 25.290 128.955 98.575 ;
   LAYER M4 ;
    RECT 126.155 25.290 126.855 98.575 ;
   LAYER M4 ;
    RECT 125.105 25.400 125.805 98.575 ;
   LAYER M4 ;
    RECT 124.055 25.290 124.755 98.575 ;
   LAYER M4 ;
    RECT 121.955 25.290 122.655 98.575 ;
   LAYER M4 ;
    RECT 119.855 25.290 120.555 98.575 ;
   LAYER M4 ;
    RECT 117.755 25.290 118.455 98.575 ;
   LAYER M4 ;
    RECT 115.655 25.290 116.355 98.575 ;
   LAYER M4 ;
    RECT 113.555 25.290 114.255 98.575 ;
   LAYER M4 ;
    RECT 111.455 25.290 112.155 98.575 ;
   LAYER M4 ;
    RECT 109.355 25.290 110.055 98.575 ;
   LAYER M4 ;
    RECT 108.305 25.400 109.005 98.575 ;
   LAYER M4 ;
    RECT 107.255 25.290 107.955 98.575 ;
   LAYER M4 ;
    RECT 105.155 25.290 105.855 98.575 ;
   LAYER M4 ;
    RECT 103.055 25.290 103.755 98.575 ;
   LAYER M4 ;
    RECT 100.955 25.290 101.655 98.575 ;
   LAYER M4 ;
    RECT 98.855 25.290 99.555 98.575 ;
   LAYER M4 ;
    RECT 96.755 25.290 97.455 98.575 ;
   LAYER M4 ;
    RECT 94.655 25.290 95.355 98.575 ;
   LAYER M4 ;
    RECT 92.555 25.290 93.255 98.575 ;
   LAYER M4 ;
    RECT 91.505 25.400 92.205 98.575 ;
   LAYER M4 ;
    RECT 90.455 25.290 91.155 98.575 ;
   LAYER M4 ;
    RECT 88.355 25.290 89.055 98.575 ;
   LAYER M4 ;
    RECT 86.255 25.290 86.955 98.575 ;
   LAYER M4 ;
    RECT 84.155 25.290 84.855 98.575 ;
   LAYER M4 ;
    RECT 82.055 25.290 82.755 98.575 ;
   LAYER M4 ;
    RECT 79.955 25.290 80.655 98.575 ;
   LAYER M4 ;
    RECT 77.855 25.290 78.555 98.575 ;
   LAYER M4 ;
    RECT 0.495 1.725 371.120 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 371.120 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 371.120 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 371.120 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 371.120 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 371.120 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 371.120 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 371.120 23.605 ;
   LAYER M4 ;
    RECT 369.735 25.290 370.115 98.575 ;
   LAYER M4 ;
    RECT 368.695 25.290 369.395 98.575 ;
   LAYER M4 ;
    RECT 366.595 25.290 367.295 98.575 ;
   LAYER M4 ;
    RECT 364.495 25.290 365.195 98.575 ;
   LAYER M4 ;
    RECT 362.395 25.290 363.095 98.575 ;
   LAYER M4 ;
    RECT 360.295 25.290 360.995 98.575 ;
   LAYER M4 ;
    RECT 359.245 25.400 359.945 98.575 ;
   LAYER M4 ;
    RECT 358.195 25.290 358.895 98.575 ;
   LAYER M4 ;
    RECT 356.095 25.290 356.795 98.575 ;
   LAYER M4 ;
    RECT 353.995 25.290 354.695 98.575 ;
   LAYER M4 ;
    RECT 351.895 25.290 352.595 98.575 ;
   LAYER M4 ;
    RECT 349.795 25.290 350.495 98.575 ;
   LAYER M4 ;
    RECT 347.695 25.290 348.395 98.575 ;
   LAYER M4 ;
    RECT 345.595 25.290 346.295 98.575 ;
   LAYER M4 ;
    RECT 343.495 25.290 344.195 98.575 ;
   LAYER M4 ;
    RECT 342.445 25.400 343.145 98.575 ;
   LAYER M4 ;
    RECT 341.395 25.290 342.095 98.575 ;
   LAYER M4 ;
    RECT 339.295 25.290 339.995 98.575 ;
   LAYER M4 ;
    RECT 337.195 25.290 337.895 98.575 ;
   LAYER M4 ;
    RECT 335.095 25.290 335.795 98.575 ;
   LAYER M4 ;
    RECT 332.995 25.290 333.695 98.575 ;
   LAYER M4 ;
    RECT 330.895 25.290 331.595 98.575 ;
   LAYER M4 ;
    RECT 328.795 25.290 329.495 98.575 ;
   LAYER M4 ;
    RECT 326.695 25.290 327.395 98.575 ;
   LAYER M4 ;
    RECT 325.645 25.400 326.345 98.575 ;
   LAYER M4 ;
    RECT 324.595 25.290 325.295 98.575 ;
   LAYER M4 ;
    RECT 322.495 25.290 323.195 98.575 ;
   LAYER M4 ;
    RECT 320.395 25.290 321.095 98.575 ;
   LAYER M4 ;
    RECT 318.295 25.290 318.995 98.575 ;
   LAYER M4 ;
    RECT 316.195 25.290 316.895 98.575 ;
   LAYER M4 ;
    RECT 314.095 25.290 314.795 98.575 ;
   LAYER M4 ;
    RECT 311.995 25.290 312.695 98.575 ;
   LAYER M4 ;
    RECT 309.895 25.290 310.595 98.575 ;
   LAYER M4 ;
    RECT 308.845 25.400 309.545 98.575 ;
   LAYER M4 ;
    RECT 307.795 25.290 308.495 98.575 ;
   LAYER M4 ;
    RECT 305.695 25.290 306.395 98.575 ;
   LAYER M4 ;
    RECT 303.595 25.290 304.295 98.575 ;
   LAYER M4 ;
    RECT 301.495 25.290 302.195 98.575 ;
   LAYER M4 ;
    RECT 299.395 25.290 300.095 98.575 ;
   LAYER M4 ;
    RECT 297.295 25.290 297.995 98.575 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 162.905 25.290 163.605 98.575 ;
   LAYER M4 ;
    RECT 160.805 25.400 161.505 98.575 ;
   LAYER M4 ;
    RECT 156.605 25.290 157.305 98.575 ;
   LAYER M4 ;
    RECT 154.505 25.290 155.205 98.575 ;
   LAYER M4 ;
    RECT 152.405 25.290 153.105 98.575 ;
   LAYER M4 ;
    RECT 150.305 25.290 151.005 98.575 ;
   LAYER M4 ;
    RECT 148.205 25.290 148.905 98.575 ;
   LAYER M4 ;
    RECT 146.105 25.290 146.805 98.575 ;
   LAYER M4 ;
    RECT 144.005 25.400 144.705 98.575 ;
   LAYER M4 ;
    RECT 139.805 25.290 140.505 98.575 ;
   LAYER M4 ;
    RECT 137.705 25.290 138.405 98.575 ;
   LAYER M4 ;
    RECT 135.605 25.290 136.305 98.575 ;
   LAYER M4 ;
    RECT 133.505 25.290 134.205 98.575 ;
   LAYER M4 ;
    RECT 131.405 25.290 132.105 98.575 ;
   LAYER M4 ;
    RECT 129.305 25.290 130.005 98.575 ;
   LAYER M4 ;
    RECT 127.205 25.400 127.905 98.575 ;
   LAYER M4 ;
    RECT 123.005 25.290 123.705 98.575 ;
   LAYER M4 ;
    RECT 120.905 25.290 121.605 98.575 ;
   LAYER M4 ;
    RECT 118.805 25.290 119.505 98.575 ;
   LAYER M4 ;
    RECT 116.705 25.290 117.405 98.575 ;
   LAYER M4 ;
    RECT 114.605 25.290 115.305 98.575 ;
   LAYER M4 ;
    RECT 112.505 25.290 113.205 98.575 ;
   LAYER M4 ;
    RECT 110.405 25.400 111.105 98.575 ;
   LAYER M4 ;
    RECT 106.205 25.290 106.905 98.575 ;
   LAYER M4 ;
    RECT 104.105 25.290 104.805 98.575 ;
   LAYER M4 ;
    RECT 102.005 25.290 102.705 98.575 ;
   LAYER M4 ;
    RECT 99.905 25.290 100.605 98.575 ;
   LAYER M4 ;
    RECT 97.805 25.290 98.505 98.575 ;
   LAYER M4 ;
    RECT 95.705 25.290 96.405 98.575 ;
   LAYER M4 ;
    RECT 93.605 25.400 94.305 98.575 ;
   LAYER M4 ;
    RECT 89.405 25.290 90.105 98.575 ;
   LAYER M4 ;
    RECT 87.305 25.290 88.005 98.575 ;
   LAYER M4 ;
    RECT 85.205 25.290 85.905 98.575 ;
   LAYER M4 ;
    RECT 83.105 25.290 83.805 98.575 ;
   LAYER M4 ;
    RECT 81.005 25.290 81.705 98.575 ;
   LAYER M4 ;
    RECT 78.905 25.290 79.605 98.575 ;
   LAYER M4 ;
    RECT 76.805 25.400 77.505 98.575 ;
   LAYER M4 ;
    RECT 72.605 25.290 73.305 98.575 ;
   LAYER M4 ;
    RECT 70.505 25.290 71.205 98.575 ;
   LAYER M4 ;
    RECT 68.405 25.290 69.105 98.575 ;
   LAYER M4 ;
    RECT 66.305 25.290 67.005 98.575 ;
   LAYER M4 ;
    RECT 64.205 25.290 64.905 98.575 ;
   LAYER M4 ;
    RECT 62.105 25.290 62.805 98.575 ;
   LAYER M4 ;
    RECT 60.005 25.400 60.705 98.575 ;
   LAYER M4 ;
    RECT 55.805 25.290 56.505 98.575 ;
   LAYER M4 ;
    RECT 53.705 25.290 54.405 98.575 ;
   LAYER M4 ;
    RECT 51.605 25.290 52.305 98.575 ;
   LAYER M4 ;
    RECT 49.505 25.290 50.205 98.575 ;
   LAYER M4 ;
    RECT 47.405 25.290 48.105 98.575 ;
   LAYER M4 ;
    RECT 45.305 25.290 46.005 98.575 ;
   LAYER M4 ;
    RECT 43.205 25.400 43.905 98.575 ;
   LAYER M4 ;
    RECT 39.005 25.290 39.705 98.575 ;
   LAYER M4 ;
    RECT 36.905 25.290 37.605 98.575 ;
   LAYER M4 ;
    RECT 34.805 25.290 35.505 98.575 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 98.575 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 98.575 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 98.575 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 98.575 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 98.575 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 98.575 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 98.575 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 98.575 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 98.575 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 98.575 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 98.575 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 98.575 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 98.575 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 98.575 ;
   LAYER M4 ;
    RECT 0.495 0.760 371.120 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 371.120 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 371.120 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 371.120 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 371.120 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 371.120 11.960 ;
   LAYER M4 ;
    RECT 0.495 14.840 371.120 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 371.120 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 371.120 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 371.120 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 371.120 25.115 ;
   LAYER M4 ;
    RECT 367.645 25.290 368.345 98.575 ;
   LAYER M4 ;
    RECT 365.545 25.290 366.245 98.575 ;
   LAYER M4 ;
    RECT 363.445 25.290 364.145 98.575 ;
   LAYER M4 ;
    RECT 361.345 25.400 362.045 98.575 ;
   LAYER M4 ;
    RECT 357.145 25.290 357.845 98.575 ;
   LAYER M4 ;
    RECT 355.045 25.290 355.745 98.575 ;
   LAYER M4 ;
    RECT 352.945 25.290 353.645 98.575 ;
   LAYER M4 ;
    RECT 350.845 25.290 351.545 98.575 ;
   LAYER M4 ;
    RECT 348.745 25.290 349.445 98.575 ;
   LAYER M4 ;
    RECT 346.645 25.290 347.345 98.575 ;
   LAYER M4 ;
    RECT 344.545 25.400 345.245 98.575 ;
   LAYER M4 ;
    RECT 340.345 25.290 341.045 98.575 ;
   LAYER M4 ;
    RECT 338.245 25.290 338.945 98.575 ;
   LAYER M4 ;
    RECT 336.145 25.290 336.845 98.575 ;
   LAYER M4 ;
    RECT 334.045 25.290 334.745 98.575 ;
   LAYER M4 ;
    RECT 331.945 25.290 332.645 98.575 ;
   LAYER M4 ;
    RECT 329.845 25.290 330.545 98.575 ;
   LAYER M4 ;
    RECT 327.745 25.400 328.445 98.575 ;
   LAYER M4 ;
    RECT 323.545 25.290 324.245 98.575 ;
   LAYER M4 ;
    RECT 321.445 25.290 322.145 98.575 ;
   LAYER M4 ;
    RECT 319.345 25.290 320.045 98.575 ;
   LAYER M4 ;
    RECT 317.245 25.290 317.945 98.575 ;
   LAYER M4 ;
    RECT 315.145 25.290 315.845 98.575 ;
   LAYER M4 ;
    RECT 313.045 25.290 313.745 98.575 ;
   LAYER M4 ;
    RECT 310.945 25.400 311.645 98.575 ;
   LAYER M4 ;
    RECT 306.745 25.290 307.445 98.575 ;
   LAYER M4 ;
    RECT 304.645 25.290 305.345 98.575 ;
   LAYER M4 ;
    RECT 302.545 25.290 303.245 98.575 ;
   LAYER M4 ;
    RECT 300.445 25.290 301.145 98.575 ;
   LAYER M4 ;
    RECT 298.345 25.290 299.045 98.575 ;
   LAYER M4 ;
    RECT 296.245 25.290 296.945 98.575 ;
   LAYER M4 ;
    RECT 294.145 25.400 294.845 98.575 ;
   LAYER M4 ;
    RECT 289.945 25.290 290.645 98.575 ;
   LAYER M4 ;
    RECT 287.845 25.290 288.545 98.575 ;
   LAYER M4 ;
    RECT 285.745 25.290 286.445 98.575 ;
   LAYER M4 ;
    RECT 283.645 25.290 284.345 98.575 ;
   LAYER M4 ;
    RECT 281.545 25.290 282.245 98.575 ;
   LAYER M4 ;
    RECT 279.445 25.290 280.145 98.575 ;
   LAYER M4 ;
    RECT 277.345 25.400 278.045 98.575 ;
   LAYER M4 ;
    RECT 273.145 25.290 273.845 98.575 ;
   LAYER M4 ;
    RECT 271.045 25.290 271.745 98.575 ;
   LAYER M4 ;
    RECT 268.945 25.290 269.645 98.575 ;
   LAYER M4 ;
    RECT 266.845 25.290 267.545 98.575 ;
   LAYER M4 ;
    RECT 264.745 25.290 265.445 98.575 ;
   LAYER M4 ;
    RECT 262.645 25.290 263.345 98.575 ;
   LAYER M4 ;
    RECT 260.545 25.400 261.245 98.575 ;
   LAYER M4 ;
    RECT 256.345 25.290 257.045 98.575 ;
   LAYER M4 ;
    RECT 254.245 25.290 254.945 98.575 ;
   LAYER M4 ;
    RECT 252.145 25.290 252.845 98.575 ;
   LAYER M4 ;
    RECT 250.045 25.290 250.745 98.575 ;
   LAYER M4 ;
    RECT 247.945 25.290 248.645 98.575 ;
   LAYER M4 ;
    RECT 245.845 25.290 246.545 98.575 ;
   LAYER M4 ;
    RECT 243.745 25.400 244.445 98.575 ;
   LAYER M4 ;
    RECT 239.545 25.290 240.245 98.575 ;
   LAYER M4 ;
    RECT 237.445 25.290 238.145 98.575 ;
   LAYER M4 ;
    RECT 235.345 25.290 236.045 98.575 ;
   LAYER M4 ;
    RECT 233.245 25.290 233.945 98.575 ;
   LAYER M4 ;
    RECT 231.145 25.290 231.845 98.575 ;
   LAYER M4 ;
    RECT 229.045 25.290 229.745 98.575 ;
   LAYER M4 ;
    RECT 226.945 25.400 227.645 98.575 ;
   LAYER M4 ;
    RECT 222.745 25.290 223.445 98.575 ;
   LAYER M4 ;
    RECT 220.645 25.290 221.345 98.575 ;
   LAYER M4 ;
    RECT 218.545 25.290 219.245 98.575 ;
   LAYER M4 ;
    RECT 216.445 25.290 217.145 98.575 ;
   LAYER M4 ;
    RECT 214.345 25.290 215.045 98.575 ;
   LAYER M4 ;
    RECT 212.245 25.290 212.945 98.575 ;
   LAYER M4 ;
    RECT 210.145 25.400 210.845 98.575 ;
   LAYER M4 ;
    RECT 205.945 25.290 206.645 98.575 ;
   LAYER M4 ;
    RECT 203.845 25.290 204.545 98.575 ;
   LAYER M4 ;
    RECT 201.745 25.290 202.445 98.575 ;
   LAYER M4 ;
    RECT 199.645 25.360 200.345 98.575 ;
   LAYER M4 ;
    RECT 197.545 25.360 198.245 98.575 ;
   LAYER M4 ;
    RECT 196.335 25.360 196.715 98.575 ;
   LAYER M4 ;
    RECT 195.130 25.360 196.110 98.575 ;
   LAYER M4 ;
    RECT 193.700 25.360 194.100 98.575 ;
   LAYER M4 ;
    RECT 192.205 25.360 192.705 98.575 ;
   LAYER M4 ;
    RECT 189.345 25.360 190.405 98.575 ;
   LAYER M4 ;
    RECT 188.665 25.360 189.065 98.575 ;
   LAYER M4 ;
    RECT 186.650 25.360 187.710 98.575 ;
   LAYER M4 ;
    RECT 184.635 25.360 185.035 98.575 ;
   LAYER M4 ;
    RECT 181.970 25.360 182.925 98.575 ;
   LAYER M4 ;
    RECT 178.510 25.360 179.150 98.575 ;
   LAYER M4 ;
    RECT 176.910 25.360 177.500 98.575 ;
   LAYER M4 ;
    RECT 172.995 25.360 173.795 98.575 ;
   LAYER M4 ;
    RECT 170.730 25.360 171.370 98.575 ;
   LAYER M4 ;
    RECT 167.105 25.290 167.805 98.575 ;
   LAYER M4 ;
    RECT 165.005 25.290 165.705 98.575 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 371.950 99.350 ;
  LAYER M2 ;
   RECT 0.050 0.050 371.950 99.350 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 39.450 0.050 39.550 0.570 ;
  LAYER VIA2 ;
   RECT 40.850 0.050 40.950 0.570 ;
  LAYER VIA2 ;
   RECT 45.050 0.050 45.150 0.570 ;
  LAYER VIA2 ;
   RECT 46.450 0.050 46.550 0.570 ;
  LAYER VIA2 ;
   RECT 56.250 0.050 56.350 0.570 ;
  LAYER VIA2 ;
   RECT 57.650 0.050 57.750 0.570 ;
  LAYER VIA2 ;
   RECT 61.850 0.050 61.950 0.570 ;
  LAYER VIA2 ;
   RECT 63.250 0.050 63.350 0.570 ;
  LAYER VIA2 ;
   RECT 73.050 0.050 73.150 0.570 ;
  LAYER VIA2 ;
   RECT 74.450 0.050 74.550 0.570 ;
  LAYER VIA2 ;
   RECT 78.650 0.050 78.750 0.570 ;
  LAYER VIA2 ;
   RECT 80.050 0.050 80.150 0.570 ;
  LAYER VIA2 ;
   RECT 89.850 0.050 89.950 0.570 ;
  LAYER VIA2 ;
   RECT 91.250 0.050 91.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.450 0.050 95.550 0.570 ;
  LAYER VIA2 ;
   RECT 96.850 0.050 96.950 0.570 ;
  LAYER VIA2 ;
   RECT 106.650 0.050 106.750 0.570 ;
  LAYER VIA2 ;
   RECT 108.050 0.050 108.150 0.570 ;
  LAYER VIA2 ;
   RECT 112.250 0.050 112.350 0.570 ;
  LAYER VIA2 ;
   RECT 113.650 0.050 113.750 0.570 ;
  LAYER VIA2 ;
   RECT 123.450 0.050 123.550 0.570 ;
  LAYER VIA2 ;
   RECT 124.850 0.050 124.950 0.570 ;
  LAYER VIA2 ;
   RECT 129.050 0.050 129.150 0.570 ;
  LAYER VIA2 ;
   RECT 130.450 0.050 130.550 0.570 ;
  LAYER VIA2 ;
   RECT 140.250 0.050 140.350 0.570 ;
  LAYER VIA2 ;
   RECT 141.650 0.050 141.750 0.570 ;
  LAYER VIA2 ;
   RECT 145.850 0.050 145.950 0.570 ;
  LAYER VIA2 ;
   RECT 147.250 0.050 147.350 0.570 ;
  LAYER VIA2 ;
   RECT 157.050 0.050 157.150 0.570 ;
  LAYER VIA2 ;
   RECT 158.450 0.050 158.550 0.570 ;
  LAYER VIA2 ;
   RECT 162.650 0.050 162.750 0.570 ;
  LAYER VIA2 ;
   RECT 164.050 0.050 164.150 0.570 ;
  LAYER VIA2 ;
   RECT 171.050 0.050 171.150 0.570 ;
  LAYER VIA2 ;
   RECT 179.650 0.050 179.750 0.570 ;
  LAYER VIA2 ;
   RECT 181.050 0.050 181.150 0.570 ;
  LAYER VIA2 ;
   RECT 181.850 0.050 181.950 0.570 ;
  LAYER VIA2 ;
   RECT 182.450 0.050 182.550 0.570 ;
  LAYER VIA2 ;
   RECT 183.050 0.050 183.150 0.570 ;
  LAYER VIA2 ;
   RECT 183.850 0.050 183.950 0.570 ;
  LAYER VIA2 ;
   RECT 185.450 0.050 185.550 0.570 ;
  LAYER VIA2 ;
   RECT 186.850 0.050 186.950 0.570 ;
  LAYER VIA2 ;
   RECT 189.450 0.050 189.550 0.570 ;
  LAYER VIA2 ;
   RECT 190.050 0.050 190.150 0.570 ;
  LAYER VIA2 ;
   RECT 194.250 0.050 194.350 0.570 ;
  LAYER VIA2 ;
   RECT 194.850 0.050 194.950 0.570 ;
  LAYER VIA2 ;
   RECT 195.650 0.050 195.750 0.570 ;
  LAYER VIA2 ;
   RECT 206.450 0.050 206.550 0.570 ;
  LAYER VIA2 ;
   RECT 207.850 0.050 207.950 0.570 ;
  LAYER VIA2 ;
   RECT 211.850 0.050 211.950 0.570 ;
  LAYER VIA2 ;
   RECT 213.250 0.050 213.350 0.570 ;
  LAYER VIA2 ;
   RECT 223.250 0.050 223.350 0.570 ;
  LAYER VIA2 ;
   RECT 224.650 0.050 224.750 0.570 ;
  LAYER VIA2 ;
   RECT 228.650 0.050 228.750 0.570 ;
  LAYER VIA2 ;
   RECT 230.050 0.050 230.150 0.570 ;
  LAYER VIA2 ;
   RECT 240.050 0.050 240.150 0.570 ;
  LAYER VIA2 ;
   RECT 241.450 0.050 241.550 0.570 ;
  LAYER VIA2 ;
   RECT 245.450 0.050 245.550 0.570 ;
  LAYER VIA2 ;
   RECT 246.850 0.050 246.950 0.570 ;
  LAYER VIA2 ;
   RECT 256.850 0.050 256.950 0.570 ;
  LAYER VIA2 ;
   RECT 258.250 0.050 258.350 0.570 ;
  LAYER VIA2 ;
   RECT 262.250 0.050 262.350 0.570 ;
  LAYER VIA2 ;
   RECT 263.650 0.050 263.750 0.570 ;
  LAYER VIA2 ;
   RECT 273.650 0.050 273.750 0.570 ;
  LAYER VIA2 ;
   RECT 275.050 0.050 275.150 0.570 ;
  LAYER VIA2 ;
   RECT 279.050 0.050 279.150 0.570 ;
  LAYER VIA2 ;
   RECT 280.450 0.050 280.550 0.570 ;
  LAYER VIA2 ;
   RECT 290.450 0.050 290.550 0.570 ;
  LAYER VIA2 ;
   RECT 291.850 0.050 291.950 0.570 ;
  LAYER VIA2 ;
   RECT 295.850 0.050 295.950 0.570 ;
  LAYER VIA2 ;
   RECT 297.250 0.050 297.350 0.570 ;
  LAYER VIA2 ;
   RECT 307.250 0.050 307.350 0.570 ;
  LAYER VIA2 ;
   RECT 308.650 0.050 308.750 0.570 ;
  LAYER VIA2 ;
   RECT 312.650 0.050 312.750 0.570 ;
  LAYER VIA2 ;
   RECT 314.050 0.050 314.150 0.570 ;
  LAYER VIA2 ;
   RECT 324.050 0.050 324.150 0.570 ;
  LAYER VIA2 ;
   RECT 325.450 0.050 325.550 0.570 ;
  LAYER VIA2 ;
   RECT 329.450 0.050 329.550 0.570 ;
  LAYER VIA2 ;
   RECT 330.850 0.050 330.950 0.570 ;
  LAYER VIA2 ;
   RECT 340.850 0.050 340.950 0.570 ;
  LAYER VIA2 ;
   RECT 342.250 0.050 342.350 0.570 ;
  LAYER VIA2 ;
   RECT 346.250 0.050 346.350 0.570 ;
  LAYER VIA2 ;
   RECT 347.650 0.050 347.750 0.570 ;
  LAYER VIA2 ;
   RECT 357.650 0.050 357.750 0.570 ;
  LAYER VIA2 ;
   RECT 359.050 0.050 359.150 0.570 ;
  LAYER VIA2 ;
   RECT 363.050 0.050 363.150 0.570 ;
  LAYER VIA2 ;
   RECT 364.450 0.050 364.550 0.570 ;
  LAYER VIA2 ;
   RECT 370.250 0.050 370.350 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 371.950 99.350 ;
  LAYER M4 ;
   RECT 0.050 0.050 371.950 99.350 ;
 END
END ST_SPHDL_1024x40m8_L

MACRO ST_SPHDL_128x32m8_L
 CLASS BLOCK ;
   SIZE 304.800 BY 41.000 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.250 0.050 148.350 0.570 ;
   LAYER M3 ;
    RECT 148.250 0.050 148.350 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.850 0.050 148.950 0.570 ;
   LAYER M3 ;
    RECT 148.850 0.050 148.950 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 149.450 0.050 149.550 0.570 ;
   LAYER M3 ;
    RECT 149.450 0.050 149.550 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 155.850 0.050 155.950 0.570 ;
   LAYER M3 ;
    RECT 155.850 0.050 155.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 156.450 0.050 156.550 0.570 ;
   LAYER M3 ;
    RECT 156.450 0.050 156.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 150.250 0.050 150.350 0.570 ;
   LAYER M3 ;
    RECT 150.250 0.050 150.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 151.850 0.050 151.950 0.570 ;
   LAYER M3 ;
    RECT 151.850 0.050 151.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 160.650 0.050 160.750 0.570 ;
   LAYER M3 ;
    RECT 160.650 0.050 160.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 162.050 0.050 162.150 0.570 ;
   LAYER M3 ;
    RECT 162.050 0.050 162.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 91.250 0.050 91.350 0.570 ;
   LAYER M3 ;
    RECT 91.250 0.050 91.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[10]
 PIN D[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 95.450 0.050 95.550 0.570 ;
   LAYER M3 ;
    RECT 95.450 0.050 95.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[11]
 PIN D[12]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 108.050 0.050 108.150 0.570 ;
   LAYER M3 ;
    RECT 108.050 0.050 108.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[12]
 PIN D[13]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 112.250 0.050 112.350 0.570 ;
   LAYER M3 ;
    RECT 112.250 0.050 112.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[13]
 PIN D[14]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 124.850 0.050 124.950 0.570 ;
   LAYER M3 ;
    RECT 124.850 0.050 124.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[14]
 PIN D[15]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 129.050 0.050 129.150 0.570 ;
   LAYER M3 ;
    RECT 129.050 0.050 129.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[15]
 PIN D[16]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 174.250 0.050 174.350 0.570 ;
   LAYER M3 ;
    RECT 174.250 0.050 174.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[16]
 PIN D[17]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 178.250 0.050 178.350 0.570 ;
   LAYER M3 ;
    RECT 178.250 0.050 178.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[17]
 PIN D[18]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 191.050 0.050 191.150 0.570 ;
   LAYER M3 ;
    RECT 191.050 0.050 191.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[18]
 PIN D[19]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 195.050 0.050 195.150 0.570 ;
   LAYER M3 ;
    RECT 195.050 0.050 195.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[19]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[20]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 207.850 0.050 207.950 0.570 ;
   LAYER M3 ;
    RECT 207.850 0.050 207.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[20]
 PIN D[21]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 211.850 0.050 211.950 0.570 ;
   LAYER M3 ;
    RECT 211.850 0.050 211.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[21]
 PIN D[22]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 224.650 0.050 224.750 0.570 ;
   LAYER M3 ;
    RECT 224.650 0.050 224.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[22]
 PIN D[23]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 228.650 0.050 228.750 0.570 ;
   LAYER M3 ;
    RECT 228.650 0.050 228.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[23]
 PIN D[24]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 241.450 0.050 241.550 0.570 ;
   LAYER M3 ;
    RECT 241.450 0.050 241.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[24]
 PIN D[25]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 245.450 0.050 245.550 0.570 ;
   LAYER M3 ;
    RECT 245.450 0.050 245.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[25]
 PIN D[26]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 258.250 0.050 258.350 0.570 ;
   LAYER M3 ;
    RECT 258.250 0.050 258.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[26]
 PIN D[27]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 262.250 0.050 262.350 0.570 ;
   LAYER M3 ;
    RECT 262.250 0.050 262.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[27]
 PIN D[28]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 275.050 0.050 275.150 0.570 ;
   LAYER M3 ;
    RECT 275.050 0.050 275.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[28]
 PIN D[29]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 279.050 0.050 279.150 0.570 ;
   LAYER M3 ;
    RECT 279.050 0.050 279.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[29]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[30]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 291.850 0.050 291.950 0.570 ;
   LAYER M3 ;
    RECT 291.850 0.050 291.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[30]
 PIN D[31]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 295.850 0.050 295.950 0.570 ;
   LAYER M3 ;
    RECT 295.850 0.050 295.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[31]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 40.850 0.050 40.950 0.570 ;
   LAYER M3 ;
    RECT 40.850 0.050 40.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 45.050 0.050 45.150 0.570 ;
   LAYER M3 ;
    RECT 45.050 0.050 45.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 57.650 0.050 57.750 0.570 ;
   LAYER M3 ;
    RECT 57.650 0.050 57.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 61.850 0.050 61.950 0.570 ;
   LAYER M3 ;
    RECT 61.850 0.050 61.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN D[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 74.450 0.050 74.550 0.570 ;
   LAYER M3 ;
    RECT 74.450 0.050 74.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[8]
 PIN D[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 78.650 0.050 78.750 0.570 ;
   LAYER M3 ;
    RECT 78.650 0.050 78.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[9]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[10]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 89.850 0.050 89.950 0.570 ;
   LAYER M3 ;
    RECT 89.850 0.050 89.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[10]
 PIN Q[11]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 96.850 0.050 96.950 0.570 ;
   LAYER M3 ;
    RECT 96.850 0.050 96.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[11]
 PIN Q[12]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 106.650 0.050 106.750 0.570 ;
   LAYER M3 ;
    RECT 106.650 0.050 106.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[12]
 PIN Q[13]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 113.650 0.050 113.750 0.570 ;
   LAYER M3 ;
    RECT 113.650 0.050 113.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[13]
 PIN Q[14]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 123.450 0.050 123.550 0.570 ;
   LAYER M3 ;
    RECT 123.450 0.050 123.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[14]
 PIN Q[15]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 130.450 0.050 130.550 0.570 ;
   LAYER M3 ;
    RECT 130.450 0.050 130.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[15]
 PIN Q[16]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 172.850 0.050 172.950 0.570 ;
   LAYER M3 ;
    RECT 172.850 0.050 172.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[16]
 PIN Q[17]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 179.650 0.050 179.750 0.570 ;
   LAYER M3 ;
    RECT 179.650 0.050 179.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[17]
 PIN Q[18]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 189.650 0.050 189.750 0.570 ;
   LAYER M3 ;
    RECT 189.650 0.050 189.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[18]
 PIN Q[19]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 196.450 0.050 196.550 0.570 ;
   LAYER M3 ;
    RECT 196.450 0.050 196.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[19]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[20]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 206.450 0.050 206.550 0.570 ;
   LAYER M3 ;
    RECT 206.450 0.050 206.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[20]
 PIN Q[21]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 213.250 0.050 213.350 0.570 ;
   LAYER M3 ;
    RECT 213.250 0.050 213.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[21]
 PIN Q[22]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 223.250 0.050 223.350 0.570 ;
   LAYER M3 ;
    RECT 223.250 0.050 223.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[22]
 PIN Q[23]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 230.050 0.050 230.150 0.570 ;
   LAYER M3 ;
    RECT 230.050 0.050 230.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[23]
 PIN Q[24]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 240.050 0.050 240.150 0.570 ;
   LAYER M3 ;
    RECT 240.050 0.050 240.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[24]
 PIN Q[25]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 246.850 0.050 246.950 0.570 ;
   LAYER M3 ;
    RECT 246.850 0.050 246.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[25]
 PIN Q[26]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 256.850 0.050 256.950 0.570 ;
   LAYER M3 ;
    RECT 256.850 0.050 256.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[26]
 PIN Q[27]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 263.650 0.050 263.750 0.570 ;
   LAYER M3 ;
    RECT 263.650 0.050 263.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[27]
 PIN Q[28]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 273.650 0.050 273.750 0.570 ;
   LAYER M3 ;
    RECT 273.650 0.050 273.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[28]
 PIN Q[29]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 280.450 0.050 280.550 0.570 ;
   LAYER M3 ;
    RECT 280.450 0.050 280.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[29]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[30]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 290.450 0.050 290.550 0.570 ;
   LAYER M3 ;
    RECT 290.450 0.050 290.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[30]
 PIN Q[31]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 297.250 0.050 297.350 0.570 ;
   LAYER M3 ;
    RECT 297.250 0.050 297.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[31]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 39.450 0.050 39.550 0.570 ;
   LAYER M3 ;
    RECT 39.450 0.050 39.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 46.450 0.050 46.550 0.570 ;
   LAYER M3 ;
    RECT 46.450 0.050 46.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 56.250 0.050 56.350 0.570 ;
   LAYER M3 ;
    RECT 56.250 0.050 56.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 63.250 0.050 63.350 0.570 ;
   LAYER M3 ;
    RECT 63.250 0.050 63.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN Q[8]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 73.050 0.050 73.150 0.570 ;
   LAYER M3 ;
    RECT 73.050 0.050 73.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[8]
 PIN Q[9]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 80.050 0.050 80.150 0.570 ;
   LAYER M3 ;
    RECT 80.050 0.050 80.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[9]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 303.050 0.050 303.150 0.570 ;
   LAYER M3 ;
    RECT 303.050 0.050 303.150 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 161.250 0.050 161.350 0.570 ;
   LAYER M3 ;
    RECT 161.250 0.050 161.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 153.250 0.050 153.350 0.570 ;
   LAYER M3 ;
    RECT 153.250 0.050 153.350 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 146.820 25.360 147.620 40.775 ;
   LAYER M4 ;
    RECT 145.825 25.360 146.225 40.775 ;
   LAYER M4 ;
    RECT 144.220 25.360 144.620 40.775 ;
   LAYER M4 ;
    RECT 142.005 25.360 142.810 40.775 ;
   LAYER M4 ;
    RECT 140.695 25.360 141.495 40.775 ;
   LAYER M4 ;
    RECT 138.275 25.360 138.895 40.775 ;
   LAYER M4 ;
    RECT 135.990 25.360 136.630 40.775 ;
   LAYER M4 ;
    RECT 134.555 25.290 135.255 40.775 ;
   LAYER M4 ;
    RECT 132.455 25.290 133.155 40.775 ;
   LAYER M4 ;
    RECT 130.355 25.290 131.055 40.775 ;
   LAYER M4 ;
    RECT 128.255 25.290 128.955 40.775 ;
   LAYER M4 ;
    RECT 126.155 25.290 126.855 40.775 ;
   LAYER M4 ;
    RECT 125.105 25.400 125.805 40.775 ;
   LAYER M4 ;
    RECT 124.055 25.290 124.755 40.775 ;
   LAYER M4 ;
    RECT 121.955 25.290 122.655 40.775 ;
   LAYER M4 ;
    RECT 119.855 25.290 120.555 40.775 ;
   LAYER M4 ;
    RECT 117.755 25.290 118.455 40.775 ;
   LAYER M4 ;
    RECT 115.655 25.290 116.355 40.775 ;
   LAYER M4 ;
    RECT 113.555 25.290 114.255 40.775 ;
   LAYER M4 ;
    RECT 111.455 25.290 112.155 40.775 ;
   LAYER M4 ;
    RECT 109.355 25.290 110.055 40.775 ;
   LAYER M4 ;
    RECT 108.305 25.400 109.005 40.775 ;
   LAYER M4 ;
    RECT 107.255 25.290 107.955 40.775 ;
   LAYER M4 ;
    RECT 105.155 25.290 105.855 40.775 ;
   LAYER M4 ;
    RECT 103.055 25.290 103.755 40.775 ;
   LAYER M4 ;
    RECT 100.955 25.290 101.655 40.775 ;
   LAYER M4 ;
    RECT 98.855 25.290 99.555 40.775 ;
   LAYER M4 ;
    RECT 96.755 25.290 97.455 40.775 ;
   LAYER M4 ;
    RECT 94.655 25.290 95.355 40.775 ;
   LAYER M4 ;
    RECT 92.555 25.290 93.255 40.775 ;
   LAYER M4 ;
    RECT 91.505 25.400 92.205 40.775 ;
   LAYER M4 ;
    RECT 90.455 25.290 91.155 40.775 ;
   LAYER M4 ;
    RECT 88.355 25.290 89.055 40.775 ;
   LAYER M4 ;
    RECT 86.255 25.290 86.955 40.775 ;
   LAYER M4 ;
    RECT 84.155 25.290 84.855 40.775 ;
   LAYER M4 ;
    RECT 82.055 25.290 82.755 40.775 ;
   LAYER M4 ;
    RECT 79.955 25.290 80.655 40.775 ;
   LAYER M4 ;
    RECT 77.855 25.290 78.555 40.775 ;
   LAYER M4 ;
    RECT 75.755 25.290 76.455 40.775 ;
   LAYER M4 ;
    RECT 74.705 25.400 75.405 40.775 ;
   LAYER M4 ;
    RECT 73.655 25.290 74.355 40.775 ;
   LAYER M4 ;
    RECT 71.555 25.290 72.255 40.775 ;
   LAYER M4 ;
    RECT 69.455 25.290 70.155 40.775 ;
   LAYER M4 ;
    RECT 67.355 25.290 68.055 40.775 ;
   LAYER M4 ;
    RECT 65.255 25.290 65.955 40.775 ;
   LAYER M4 ;
    RECT 63.155 25.290 63.855 40.775 ;
   LAYER M4 ;
    RECT 61.055 25.290 61.755 40.775 ;
   LAYER M4 ;
    RECT 58.955 25.290 59.655 40.775 ;
   LAYER M4 ;
    RECT 57.905 25.400 58.605 40.775 ;
   LAYER M4 ;
    RECT 56.855 25.290 57.555 40.775 ;
   LAYER M4 ;
    RECT 54.755 25.290 55.455 40.775 ;
   LAYER M4 ;
    RECT 52.655 25.290 53.355 40.775 ;
   LAYER M4 ;
    RECT 50.555 25.290 51.255 40.775 ;
   LAYER M4 ;
    RECT 48.455 25.290 49.155 40.775 ;
   LAYER M4 ;
    RECT 46.355 25.290 47.055 40.775 ;
   LAYER M4 ;
    RECT 44.255 25.290 44.955 40.775 ;
   LAYER M4 ;
    RECT 42.155 25.290 42.855 40.775 ;
   LAYER M4 ;
    RECT 41.105 25.400 41.805 40.775 ;
   LAYER M4 ;
    RECT 40.055 25.290 40.755 40.775 ;
   LAYER M4 ;
    RECT 37.955 25.290 38.655 40.775 ;
   LAYER M4 ;
    RECT 35.855 25.290 36.555 40.775 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 40.775 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 40.775 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 40.775 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 40.775 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 40.775 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 40.775 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 40.775 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 40.775 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 40.775 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 40.775 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 40.775 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 40.775 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 40.775 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 40.775 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 40.775 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 40.775 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 40.775 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 40.775 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 40.775 ;
   LAYER M4 ;
    RECT 0.495 1.725 303.920 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 303.920 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 303.920 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 303.920 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 303.920 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 303.920 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 303.920 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 303.920 23.605 ;
   LAYER M4 ;
    RECT 302.535 25.290 302.915 40.775 ;
   LAYER M4 ;
    RECT 301.495 25.290 302.195 40.775 ;
   LAYER M4 ;
    RECT 299.395 25.290 300.095 40.775 ;
   LAYER M4 ;
    RECT 297.295 25.290 297.995 40.775 ;
   LAYER M4 ;
    RECT 295.195 25.290 295.895 40.775 ;
   LAYER M4 ;
    RECT 293.095 25.290 293.795 40.775 ;
   LAYER M4 ;
    RECT 292.045 25.400 292.745 40.775 ;
   LAYER M4 ;
    RECT 290.995 25.290 291.695 40.775 ;
   LAYER M4 ;
    RECT 288.895 25.290 289.595 40.775 ;
   LAYER M4 ;
    RECT 286.795 25.290 287.495 40.775 ;
   LAYER M4 ;
    RECT 284.695 25.290 285.395 40.775 ;
   LAYER M4 ;
    RECT 282.595 25.290 283.295 40.775 ;
   LAYER M4 ;
    RECT 280.495 25.290 281.195 40.775 ;
   LAYER M4 ;
    RECT 278.395 25.290 279.095 40.775 ;
   LAYER M4 ;
    RECT 276.295 25.290 276.995 40.775 ;
   LAYER M4 ;
    RECT 275.245 25.400 275.945 40.775 ;
   LAYER M4 ;
    RECT 274.195 25.290 274.895 40.775 ;
   LAYER M4 ;
    RECT 272.095 25.290 272.795 40.775 ;
   LAYER M4 ;
    RECT 269.995 25.290 270.695 40.775 ;
   LAYER M4 ;
    RECT 267.895 25.290 268.595 40.775 ;
   LAYER M4 ;
    RECT 265.795 25.290 266.495 40.775 ;
   LAYER M4 ;
    RECT 263.695 25.290 264.395 40.775 ;
   LAYER M4 ;
    RECT 261.595 25.290 262.295 40.775 ;
   LAYER M4 ;
    RECT 259.495 25.290 260.195 40.775 ;
   LAYER M4 ;
    RECT 258.445 25.400 259.145 40.775 ;
   LAYER M4 ;
    RECT 257.395 25.290 258.095 40.775 ;
   LAYER M4 ;
    RECT 255.295 25.290 255.995 40.775 ;
   LAYER M4 ;
    RECT 253.195 25.290 253.895 40.775 ;
   LAYER M4 ;
    RECT 251.095 25.290 251.795 40.775 ;
   LAYER M4 ;
    RECT 248.995 25.290 249.695 40.775 ;
   LAYER M4 ;
    RECT 246.895 25.290 247.595 40.775 ;
   LAYER M4 ;
    RECT 244.795 25.290 245.495 40.775 ;
   LAYER M4 ;
    RECT 242.695 25.290 243.395 40.775 ;
   LAYER M4 ;
    RECT 241.645 25.400 242.345 40.775 ;
   LAYER M4 ;
    RECT 240.595 25.290 241.295 40.775 ;
   LAYER M4 ;
    RECT 238.495 25.290 239.195 40.775 ;
   LAYER M4 ;
    RECT 236.395 25.290 237.095 40.775 ;
   LAYER M4 ;
    RECT 234.295 25.290 234.995 40.775 ;
   LAYER M4 ;
    RECT 232.195 25.290 232.895 40.775 ;
   LAYER M4 ;
    RECT 230.095 25.290 230.795 40.775 ;
   LAYER M4 ;
    RECT 227.995 25.290 228.695 40.775 ;
   LAYER M4 ;
    RECT 225.895 25.290 226.595 40.775 ;
   LAYER M4 ;
    RECT 224.845 25.400 225.545 40.775 ;
   LAYER M4 ;
    RECT 223.795 25.290 224.495 40.775 ;
   LAYER M4 ;
    RECT 221.695 25.290 222.395 40.775 ;
   LAYER M4 ;
    RECT 219.595 25.290 220.295 40.775 ;
   LAYER M4 ;
    RECT 217.495 25.290 218.195 40.775 ;
   LAYER M4 ;
    RECT 215.395 25.290 216.095 40.775 ;
   LAYER M4 ;
    RECT 213.295 25.290 213.995 40.775 ;
   LAYER M4 ;
    RECT 211.195 25.290 211.895 40.775 ;
   LAYER M4 ;
    RECT 209.095 25.290 209.795 40.775 ;
   LAYER M4 ;
    RECT 208.045 25.400 208.745 40.775 ;
   LAYER M4 ;
    RECT 206.995 25.290 207.695 40.775 ;
   LAYER M4 ;
    RECT 204.895 25.290 205.595 40.775 ;
   LAYER M4 ;
    RECT 202.795 25.290 203.495 40.775 ;
   LAYER M4 ;
    RECT 200.695 25.290 201.395 40.775 ;
   LAYER M4 ;
    RECT 198.595 25.290 199.295 40.775 ;
   LAYER M4 ;
    RECT 196.495 25.290 197.195 40.775 ;
   LAYER M4 ;
    RECT 194.395 25.290 195.095 40.775 ;
   LAYER M4 ;
    RECT 192.295 25.290 192.995 40.775 ;
   LAYER M4 ;
    RECT 191.245 25.400 191.945 40.775 ;
   LAYER M4 ;
    RECT 190.195 25.290 190.895 40.775 ;
   LAYER M4 ;
    RECT 188.095 25.290 188.795 40.775 ;
   LAYER M4 ;
    RECT 185.995 25.290 186.695 40.775 ;
   LAYER M4 ;
    RECT 183.895 25.290 184.595 40.775 ;
   LAYER M4 ;
    RECT 181.795 25.290 182.495 40.775 ;
   LAYER M4 ;
    RECT 179.695 25.290 180.395 40.775 ;
   LAYER M4 ;
    RECT 177.595 25.290 178.295 40.775 ;
   LAYER M4 ;
    RECT 175.495 25.290 176.195 40.775 ;
   LAYER M4 ;
    RECT 174.445 25.400 175.145 40.775 ;
   LAYER M4 ;
    RECT 173.395 25.290 174.095 40.775 ;
   LAYER M4 ;
    RECT 171.295 25.290 171.995 40.775 ;
   LAYER M4 ;
    RECT 169.195 25.290 169.895 40.775 ;
   LAYER M4 ;
    RECT 167.095 25.360 167.795 40.775 ;
   LAYER M4 ;
    RECT 164.995 25.360 165.695 40.775 ;
   LAYER M4 ;
    RECT 163.310 25.360 163.690 40.775 ;
   LAYER M4 ;
    RECT 160.815 25.360 161.215 40.775 ;
   LAYER M4 ;
    RECT 159.345 25.360 159.845 40.775 ;
   LAYER M4 ;
    RECT 157.295 25.360 158.355 40.775 ;
   LAYER M4 ;
    RECT 154.390 25.360 154.790 40.775 ;
   LAYER M4 ;
    RECT 151.745 25.360 152.345 40.775 ;
   LAYER M4 ;
    RECT 150.075 25.360 150.720 40.775 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 62.105 25.290 62.805 40.775 ;
   LAYER M4 ;
    RECT 60.005 25.400 60.705 40.775 ;
   LAYER M4 ;
    RECT 55.805 25.290 56.505 40.775 ;
   LAYER M4 ;
    RECT 53.705 25.290 54.405 40.775 ;
   LAYER M4 ;
    RECT 51.605 25.290 52.305 40.775 ;
   LAYER M4 ;
    RECT 49.505 25.290 50.205 40.775 ;
   LAYER M4 ;
    RECT 47.405 25.290 48.105 40.775 ;
   LAYER M4 ;
    RECT 45.305 25.290 46.005 40.775 ;
   LAYER M4 ;
    RECT 43.205 25.400 43.905 40.775 ;
   LAYER M4 ;
    RECT 39.005 25.290 39.705 40.775 ;
   LAYER M4 ;
    RECT 36.905 25.290 37.605 40.775 ;
   LAYER M4 ;
    RECT 34.805 25.290 35.505 40.775 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 40.775 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 40.775 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 40.775 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 40.775 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 40.775 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 40.775 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 40.775 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 40.775 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 40.775 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 40.775 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 40.775 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 40.775 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 40.775 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 40.775 ;
   LAYER M4 ;
    RECT 0.495 0.760 303.920 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 303.920 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 303.920 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 303.920 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 303.920 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 303.920 11.960 ;
   LAYER M4 ;
    RECT 0.495 14.840 303.920 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 303.920 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 303.920 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 303.920 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 303.920 25.115 ;
   LAYER M4 ;
    RECT 300.445 25.290 301.145 40.775 ;
   LAYER M4 ;
    RECT 298.345 25.290 299.045 40.775 ;
   LAYER M4 ;
    RECT 296.245 25.290 296.945 40.775 ;
   LAYER M4 ;
    RECT 294.145 25.400 294.845 40.775 ;
   LAYER M4 ;
    RECT 289.945 25.290 290.645 40.775 ;
   LAYER M4 ;
    RECT 287.845 25.290 288.545 40.775 ;
   LAYER M4 ;
    RECT 285.745 25.290 286.445 40.775 ;
   LAYER M4 ;
    RECT 283.645 25.290 284.345 40.775 ;
   LAYER M4 ;
    RECT 281.545 25.290 282.245 40.775 ;
   LAYER M4 ;
    RECT 279.445 25.290 280.145 40.775 ;
   LAYER M4 ;
    RECT 277.345 25.400 278.045 40.775 ;
   LAYER M4 ;
    RECT 273.145 25.290 273.845 40.775 ;
   LAYER M4 ;
    RECT 271.045 25.290 271.745 40.775 ;
   LAYER M4 ;
    RECT 268.945 25.290 269.645 40.775 ;
   LAYER M4 ;
    RECT 266.845 25.290 267.545 40.775 ;
   LAYER M4 ;
    RECT 264.745 25.290 265.445 40.775 ;
   LAYER M4 ;
    RECT 262.645 25.290 263.345 40.775 ;
   LAYER M4 ;
    RECT 260.545 25.400 261.245 40.775 ;
   LAYER M4 ;
    RECT 256.345 25.290 257.045 40.775 ;
   LAYER M4 ;
    RECT 254.245 25.290 254.945 40.775 ;
   LAYER M4 ;
    RECT 252.145 25.290 252.845 40.775 ;
   LAYER M4 ;
    RECT 250.045 25.290 250.745 40.775 ;
   LAYER M4 ;
    RECT 247.945 25.290 248.645 40.775 ;
   LAYER M4 ;
    RECT 245.845 25.290 246.545 40.775 ;
   LAYER M4 ;
    RECT 243.745 25.400 244.445 40.775 ;
   LAYER M4 ;
    RECT 239.545 25.290 240.245 40.775 ;
   LAYER M4 ;
    RECT 237.445 25.290 238.145 40.775 ;
   LAYER M4 ;
    RECT 235.345 25.290 236.045 40.775 ;
   LAYER M4 ;
    RECT 233.245 25.290 233.945 40.775 ;
   LAYER M4 ;
    RECT 231.145 25.290 231.845 40.775 ;
   LAYER M4 ;
    RECT 229.045 25.290 229.745 40.775 ;
   LAYER M4 ;
    RECT 226.945 25.400 227.645 40.775 ;
   LAYER M4 ;
    RECT 222.745 25.290 223.445 40.775 ;
   LAYER M4 ;
    RECT 220.645 25.290 221.345 40.775 ;
   LAYER M4 ;
    RECT 218.545 25.290 219.245 40.775 ;
   LAYER M4 ;
    RECT 216.445 25.290 217.145 40.775 ;
   LAYER M4 ;
    RECT 214.345 25.290 215.045 40.775 ;
   LAYER M4 ;
    RECT 212.245 25.290 212.945 40.775 ;
   LAYER M4 ;
    RECT 210.145 25.400 210.845 40.775 ;
   LAYER M4 ;
    RECT 205.945 25.290 206.645 40.775 ;
   LAYER M4 ;
    RECT 203.845 25.290 204.545 40.775 ;
   LAYER M4 ;
    RECT 201.745 25.290 202.445 40.775 ;
   LAYER M4 ;
    RECT 199.645 25.290 200.345 40.775 ;
   LAYER M4 ;
    RECT 197.545 25.290 198.245 40.775 ;
   LAYER M4 ;
    RECT 195.445 25.290 196.145 40.775 ;
   LAYER M4 ;
    RECT 193.345 25.400 194.045 40.775 ;
   LAYER M4 ;
    RECT 189.145 25.290 189.845 40.775 ;
   LAYER M4 ;
    RECT 187.045 25.290 187.745 40.775 ;
   LAYER M4 ;
    RECT 184.945 25.290 185.645 40.775 ;
   LAYER M4 ;
    RECT 182.845 25.290 183.545 40.775 ;
   LAYER M4 ;
    RECT 180.745 25.290 181.445 40.775 ;
   LAYER M4 ;
    RECT 178.645 25.290 179.345 40.775 ;
   LAYER M4 ;
    RECT 176.545 25.400 177.245 40.775 ;
   LAYER M4 ;
    RECT 172.345 25.290 173.045 40.775 ;
   LAYER M4 ;
    RECT 170.245 25.290 170.945 40.775 ;
   LAYER M4 ;
    RECT 168.145 25.290 168.845 40.775 ;
   LAYER M4 ;
    RECT 166.045 25.360 166.745 40.775 ;
   LAYER M4 ;
    RECT 163.945 25.360 164.645 40.775 ;
   LAYER M4 ;
    RECT 162.735 25.360 163.115 40.775 ;
   LAYER M4 ;
    RECT 161.530 25.360 162.510 40.775 ;
   LAYER M4 ;
    RECT 160.100 25.360 160.500 40.775 ;
   LAYER M4 ;
    RECT 158.605 25.360 159.105 40.775 ;
   LAYER M4 ;
    RECT 155.745 25.360 156.805 40.775 ;
   LAYER M4 ;
    RECT 155.065 25.360 155.465 40.775 ;
   LAYER M4 ;
    RECT 153.050 25.360 154.110 40.775 ;
   LAYER M4 ;
    RECT 151.035 25.360 151.435 40.775 ;
   LAYER M4 ;
    RECT 148.370 25.360 149.325 40.775 ;
   LAYER M4 ;
    RECT 144.910 25.360 145.550 40.775 ;
   LAYER M4 ;
    RECT 143.310 25.360 143.900 40.775 ;
   LAYER M4 ;
    RECT 139.395 25.360 140.195 40.775 ;
   LAYER M4 ;
    RECT 137.130 25.360 137.770 40.775 ;
   LAYER M4 ;
    RECT 133.505 25.290 134.205 40.775 ;
   LAYER M4 ;
    RECT 131.405 25.290 132.105 40.775 ;
   LAYER M4 ;
    RECT 129.305 25.290 130.005 40.775 ;
   LAYER M4 ;
    RECT 127.205 25.400 127.905 40.775 ;
   LAYER M4 ;
    RECT 123.005 25.290 123.705 40.775 ;
   LAYER M4 ;
    RECT 120.905 25.290 121.605 40.775 ;
   LAYER M4 ;
    RECT 118.805 25.290 119.505 40.775 ;
   LAYER M4 ;
    RECT 116.705 25.290 117.405 40.775 ;
   LAYER M4 ;
    RECT 114.605 25.290 115.305 40.775 ;
   LAYER M4 ;
    RECT 112.505 25.290 113.205 40.775 ;
   LAYER M4 ;
    RECT 110.405 25.400 111.105 40.775 ;
   LAYER M4 ;
    RECT 106.205 25.290 106.905 40.775 ;
   LAYER M4 ;
    RECT 104.105 25.290 104.805 40.775 ;
   LAYER M4 ;
    RECT 102.005 25.290 102.705 40.775 ;
   LAYER M4 ;
    RECT 99.905 25.290 100.605 40.775 ;
   LAYER M4 ;
    RECT 97.805 25.290 98.505 40.775 ;
   LAYER M4 ;
    RECT 95.705 25.290 96.405 40.775 ;
   LAYER M4 ;
    RECT 93.605 25.400 94.305 40.775 ;
   LAYER M4 ;
    RECT 89.405 25.290 90.105 40.775 ;
   LAYER M4 ;
    RECT 87.305 25.290 88.005 40.775 ;
   LAYER M4 ;
    RECT 85.205 25.290 85.905 40.775 ;
   LAYER M4 ;
    RECT 83.105 25.290 83.805 40.775 ;
   LAYER M4 ;
    RECT 81.005 25.290 81.705 40.775 ;
   LAYER M4 ;
    RECT 78.905 25.290 79.605 40.775 ;
   LAYER M4 ;
    RECT 76.805 25.400 77.505 40.775 ;
   LAYER M4 ;
    RECT 72.605 25.290 73.305 40.775 ;
   LAYER M4 ;
    RECT 70.505 25.290 71.205 40.775 ;
   LAYER M4 ;
    RECT 68.405 25.290 69.105 40.775 ;
   LAYER M4 ;
    RECT 66.305 25.290 67.005 40.775 ;
   LAYER M4 ;
    RECT 64.205 25.290 64.905 40.775 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 304.750 37.950 ;
  LAYER M2 ;
   RECT 0.050 0.050 304.750 37.950 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 39.450 0.050 39.550 0.570 ;
  LAYER VIA2 ;
   RECT 40.850 0.050 40.950 0.570 ;
  LAYER VIA2 ;
   RECT 45.050 0.050 45.150 0.570 ;
  LAYER VIA2 ;
   RECT 46.450 0.050 46.550 0.570 ;
  LAYER VIA2 ;
   RECT 56.250 0.050 56.350 0.570 ;
  LAYER VIA2 ;
   RECT 57.650 0.050 57.750 0.570 ;
  LAYER VIA2 ;
   RECT 61.850 0.050 61.950 0.570 ;
  LAYER VIA2 ;
   RECT 63.250 0.050 63.350 0.570 ;
  LAYER VIA2 ;
   RECT 73.050 0.050 73.150 0.570 ;
  LAYER VIA2 ;
   RECT 74.450 0.050 74.550 0.570 ;
  LAYER VIA2 ;
   RECT 78.650 0.050 78.750 0.570 ;
  LAYER VIA2 ;
   RECT 80.050 0.050 80.150 0.570 ;
  LAYER VIA2 ;
   RECT 89.850 0.050 89.950 0.570 ;
  LAYER VIA2 ;
   RECT 91.250 0.050 91.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.450 0.050 95.550 0.570 ;
  LAYER VIA2 ;
   RECT 96.850 0.050 96.950 0.570 ;
  LAYER VIA2 ;
   RECT 106.650 0.050 106.750 0.570 ;
  LAYER VIA2 ;
   RECT 108.050 0.050 108.150 0.570 ;
  LAYER VIA2 ;
   RECT 112.250 0.050 112.350 0.570 ;
  LAYER VIA2 ;
   RECT 113.650 0.050 113.750 0.570 ;
  LAYER VIA2 ;
   RECT 123.450 0.050 123.550 0.570 ;
  LAYER VIA2 ;
   RECT 124.850 0.050 124.950 0.570 ;
  LAYER VIA2 ;
   RECT 129.050 0.050 129.150 0.570 ;
  LAYER VIA2 ;
   RECT 130.450 0.050 130.550 0.570 ;
  LAYER VIA2 ;
   RECT 148.250 0.050 148.350 0.570 ;
  LAYER VIA2 ;
   RECT 148.850 0.050 148.950 0.570 ;
  LAYER VIA2 ;
   RECT 149.450 0.050 149.550 0.570 ;
  LAYER VIA2 ;
   RECT 150.250 0.050 150.350 0.570 ;
  LAYER VIA2 ;
   RECT 151.850 0.050 151.950 0.570 ;
  LAYER VIA2 ;
   RECT 153.250 0.050 153.350 0.570 ;
  LAYER VIA2 ;
   RECT 155.850 0.050 155.950 0.570 ;
  LAYER VIA2 ;
   RECT 156.450 0.050 156.550 0.570 ;
  LAYER VIA2 ;
   RECT 160.650 0.050 160.750 0.570 ;
  LAYER VIA2 ;
   RECT 161.250 0.050 161.350 0.570 ;
  LAYER VIA2 ;
   RECT 162.050 0.050 162.150 0.570 ;
  LAYER VIA2 ;
   RECT 172.850 0.050 172.950 0.570 ;
  LAYER VIA2 ;
   RECT 174.250 0.050 174.350 0.570 ;
  LAYER VIA2 ;
   RECT 178.250 0.050 178.350 0.570 ;
  LAYER VIA2 ;
   RECT 179.650 0.050 179.750 0.570 ;
  LAYER VIA2 ;
   RECT 189.650 0.050 189.750 0.570 ;
  LAYER VIA2 ;
   RECT 191.050 0.050 191.150 0.570 ;
  LAYER VIA2 ;
   RECT 195.050 0.050 195.150 0.570 ;
  LAYER VIA2 ;
   RECT 196.450 0.050 196.550 0.570 ;
  LAYER VIA2 ;
   RECT 206.450 0.050 206.550 0.570 ;
  LAYER VIA2 ;
   RECT 207.850 0.050 207.950 0.570 ;
  LAYER VIA2 ;
   RECT 211.850 0.050 211.950 0.570 ;
  LAYER VIA2 ;
   RECT 213.250 0.050 213.350 0.570 ;
  LAYER VIA2 ;
   RECT 223.250 0.050 223.350 0.570 ;
  LAYER VIA2 ;
   RECT 224.650 0.050 224.750 0.570 ;
  LAYER VIA2 ;
   RECT 228.650 0.050 228.750 0.570 ;
  LAYER VIA2 ;
   RECT 230.050 0.050 230.150 0.570 ;
  LAYER VIA2 ;
   RECT 240.050 0.050 240.150 0.570 ;
  LAYER VIA2 ;
   RECT 241.450 0.050 241.550 0.570 ;
  LAYER VIA2 ;
   RECT 245.450 0.050 245.550 0.570 ;
  LAYER VIA2 ;
   RECT 246.850 0.050 246.950 0.570 ;
  LAYER VIA2 ;
   RECT 256.850 0.050 256.950 0.570 ;
  LAYER VIA2 ;
   RECT 258.250 0.050 258.350 0.570 ;
  LAYER VIA2 ;
   RECT 262.250 0.050 262.350 0.570 ;
  LAYER VIA2 ;
   RECT 263.650 0.050 263.750 0.570 ;
  LAYER VIA2 ;
   RECT 273.650 0.050 273.750 0.570 ;
  LAYER VIA2 ;
   RECT 275.050 0.050 275.150 0.570 ;
  LAYER VIA2 ;
   RECT 279.050 0.050 279.150 0.570 ;
  LAYER VIA2 ;
   RECT 280.450 0.050 280.550 0.570 ;
  LAYER VIA2 ;
   RECT 290.450 0.050 290.550 0.570 ;
  LAYER VIA2 ;
   RECT 291.850 0.050 291.950 0.570 ;
  LAYER VIA2 ;
   RECT 295.850 0.050 295.950 0.570 ;
  LAYER VIA2 ;
   RECT 297.250 0.050 297.350 0.570 ;
  LAYER VIA2 ;
   RECT 303.050 0.050 303.150 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 304.750 37.950 ;
  LAYER M4 ;
   RECT 0.050 0.050 304.750 40.825 ;
 END
END ST_SPHDL_128x32m8_L

MACRO ST_SPHDL_128x8m8_L
 CLASS BLOCK ;
   SIZE 103.200 BY 41.000 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 47.450 0.050 47.550 0.570 ;
   LAYER M3 ;
    RECT 47.450 0.050 47.550 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 48.050 0.050 48.150 0.570 ;
   LAYER M3 ;
    RECT 48.050 0.050 48.150 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 48.650 0.050 48.750 0.570 ;
   LAYER M3 ;
    RECT 48.650 0.050 48.750 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 55.050 0.050 55.150 0.570 ;
   LAYER M3 ;
    RECT 55.050 0.050 55.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 55.650 0.050 55.750 0.570 ;
   LAYER M3 ;
    RECT 55.650 0.050 55.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 49.450 0.050 49.550 0.570 ;
   LAYER M3 ;
    RECT 49.450 0.050 49.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 51.050 0.050 51.150 0.570 ;
   LAYER M3 ;
    RECT 51.050 0.050 51.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 59.850 0.050 59.950 0.570 ;
   LAYER M3 ;
    RECT 59.850 0.050 59.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 61.250 0.050 61.350 0.570 ;
   LAYER M3 ;
    RECT 61.250 0.050 61.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 73.450 0.050 73.550 0.570 ;
   LAYER M3 ;
    RECT 73.450 0.050 73.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 77.450 0.050 77.550 0.570 ;
   LAYER M3 ;
    RECT 77.450 0.050 77.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 90.250 0.050 90.350 0.570 ;
   LAYER M3 ;
    RECT 90.250 0.050 90.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 94.250 0.050 94.350 0.570 ;
   LAYER M3 ;
    RECT 94.250 0.050 94.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 72.050 0.050 72.150 0.570 ;
   LAYER M3 ;
    RECT 72.050 0.050 72.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 78.850 0.050 78.950 0.570 ;
   LAYER M3 ;
    RECT 78.850 0.050 78.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 88.850 0.050 88.950 0.570 ;
   LAYER M3 ;
    RECT 88.850 0.050 88.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 95.650 0.050 95.750 0.570 ;
   LAYER M3 ;
    RECT 95.650 0.050 95.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 101.450 0.050 101.550 0.570 ;
   LAYER M3 ;
    RECT 101.450 0.050 101.550 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 60.450 0.050 60.550 0.570 ;
   LAYER M3 ;
    RECT 60.450 0.050 60.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 52.450 0.050 52.550 0.570 ;
   LAYER M3 ;
    RECT 52.450 0.050 52.550 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 0.495 1.725 102.320 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 102.320 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 102.320 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 102.320 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 102.320 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 102.320 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 102.320 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 102.320 23.605 ;
   LAYER M4 ;
    RECT 100.935 25.290 101.315 40.775 ;
   LAYER M4 ;
    RECT 99.895 25.290 100.595 40.775 ;
   LAYER M4 ;
    RECT 97.795 25.290 98.495 40.775 ;
   LAYER M4 ;
    RECT 95.695 25.290 96.395 40.775 ;
   LAYER M4 ;
    RECT 93.595 25.290 94.295 40.775 ;
   LAYER M4 ;
    RECT 91.495 25.290 92.195 40.775 ;
   LAYER M4 ;
    RECT 90.445 25.400 91.145 40.775 ;
   LAYER M4 ;
    RECT 89.395 25.290 90.095 40.775 ;
   LAYER M4 ;
    RECT 87.295 25.290 87.995 40.775 ;
   LAYER M4 ;
    RECT 85.195 25.290 85.895 40.775 ;
   LAYER M4 ;
    RECT 83.095 25.290 83.795 40.775 ;
   LAYER M4 ;
    RECT 80.995 25.290 81.695 40.775 ;
   LAYER M4 ;
    RECT 78.895 25.290 79.595 40.775 ;
   LAYER M4 ;
    RECT 76.795 25.290 77.495 40.775 ;
   LAYER M4 ;
    RECT 74.695 25.290 75.395 40.775 ;
   LAYER M4 ;
    RECT 73.645 25.400 74.345 40.775 ;
   LAYER M4 ;
    RECT 72.595 25.290 73.295 40.775 ;
   LAYER M4 ;
    RECT 70.495 25.290 71.195 40.775 ;
   LAYER M4 ;
    RECT 68.395 25.290 69.095 40.775 ;
   LAYER M4 ;
    RECT 66.295 25.360 66.995 40.775 ;
   LAYER M4 ;
    RECT 64.195 25.360 64.895 40.775 ;
   LAYER M4 ;
    RECT 62.510 25.360 62.890 40.775 ;
   LAYER M4 ;
    RECT 60.015 25.360 60.415 40.775 ;
   LAYER M4 ;
    RECT 58.545 25.360 59.045 40.775 ;
   LAYER M4 ;
    RECT 56.495 25.360 57.555 40.775 ;
   LAYER M4 ;
    RECT 53.590 25.360 53.990 40.775 ;
   LAYER M4 ;
    RECT 50.945 25.360 51.545 40.775 ;
   LAYER M4 ;
    RECT 49.275 25.360 49.920 40.775 ;
   LAYER M4 ;
    RECT 46.020 25.360 46.820 40.775 ;
   LAYER M4 ;
    RECT 45.025 25.360 45.425 40.775 ;
   LAYER M4 ;
    RECT 43.420 25.360 43.820 40.775 ;
   LAYER M4 ;
    RECT 41.205 25.360 42.010 40.775 ;
   LAYER M4 ;
    RECT 39.895 25.360 40.695 40.775 ;
   LAYER M4 ;
    RECT 37.475 25.360 38.095 40.775 ;
   LAYER M4 ;
    RECT 35.190 25.360 35.830 40.775 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 40.775 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 40.775 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 40.775 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 40.775 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 40.775 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 40.775 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 40.775 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 40.775 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 40.775 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 40.775 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 40.775 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 40.775 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 40.775 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 40.775 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 40.775 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 40.775 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 40.775 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 40.775 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 40.775 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 0.495 0.760 102.320 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 102.320 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 102.320 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 102.320 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 102.320 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 102.320 11.960 ;
   LAYER M4 ;
    RECT 0.495 14.840 102.320 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 102.320 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 102.320 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 102.320 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 102.320 25.115 ;
   LAYER M4 ;
    RECT 98.845 25.290 99.545 40.775 ;
   LAYER M4 ;
    RECT 96.745 25.290 97.445 40.775 ;
   LAYER M4 ;
    RECT 94.645 25.290 95.345 40.775 ;
   LAYER M4 ;
    RECT 92.545 25.400 93.245 40.775 ;
   LAYER M4 ;
    RECT 88.345 25.290 89.045 40.775 ;
   LAYER M4 ;
    RECT 86.245 25.290 86.945 40.775 ;
   LAYER M4 ;
    RECT 84.145 25.290 84.845 40.775 ;
   LAYER M4 ;
    RECT 82.045 25.290 82.745 40.775 ;
   LAYER M4 ;
    RECT 79.945 25.290 80.645 40.775 ;
   LAYER M4 ;
    RECT 77.845 25.290 78.545 40.775 ;
   LAYER M4 ;
    RECT 75.745 25.400 76.445 40.775 ;
   LAYER M4 ;
    RECT 71.545 25.290 72.245 40.775 ;
   LAYER M4 ;
    RECT 69.445 25.290 70.145 40.775 ;
   LAYER M4 ;
    RECT 67.345 25.290 68.045 40.775 ;
   LAYER M4 ;
    RECT 65.245 25.360 65.945 40.775 ;
   LAYER M4 ;
    RECT 63.145 25.360 63.845 40.775 ;
   LAYER M4 ;
    RECT 61.935 25.360 62.315 40.775 ;
   LAYER M4 ;
    RECT 60.730 25.360 61.710 40.775 ;
   LAYER M4 ;
    RECT 59.300 25.360 59.700 40.775 ;
   LAYER M4 ;
    RECT 57.805 25.360 58.305 40.775 ;
   LAYER M4 ;
    RECT 54.945 25.360 56.005 40.775 ;
   LAYER M4 ;
    RECT 54.265 25.360 54.665 40.775 ;
   LAYER M4 ;
    RECT 52.250 25.360 53.310 40.775 ;
   LAYER M4 ;
    RECT 50.235 25.360 50.635 40.775 ;
   LAYER M4 ;
    RECT 47.570 25.360 48.525 40.775 ;
   LAYER M4 ;
    RECT 44.110 25.360 44.750 40.775 ;
   LAYER M4 ;
    RECT 42.510 25.360 43.100 40.775 ;
   LAYER M4 ;
    RECT 38.595 25.360 39.395 40.775 ;
   LAYER M4 ;
    RECT 36.330 25.360 36.970 40.775 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 40.775 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 40.775 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 40.775 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 40.775 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 40.775 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 40.775 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 40.775 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 40.775 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 40.775 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 40.775 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 40.775 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 40.775 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 40.775 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 40.775 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 103.150 37.950 ;
  LAYER M2 ;
   RECT 0.050 0.050 103.150 37.950 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 47.450 0.050 47.550 0.570 ;
  LAYER VIA2 ;
   RECT 48.050 0.050 48.150 0.570 ;
  LAYER VIA2 ;
   RECT 48.650 0.050 48.750 0.570 ;
  LAYER VIA2 ;
   RECT 49.450 0.050 49.550 0.570 ;
  LAYER VIA2 ;
   RECT 51.050 0.050 51.150 0.570 ;
  LAYER VIA2 ;
   RECT 52.450 0.050 52.550 0.570 ;
  LAYER VIA2 ;
   RECT 55.050 0.050 55.150 0.570 ;
  LAYER VIA2 ;
   RECT 55.650 0.050 55.750 0.570 ;
  LAYER VIA2 ;
   RECT 59.850 0.050 59.950 0.570 ;
  LAYER VIA2 ;
   RECT 60.450 0.050 60.550 0.570 ;
  LAYER VIA2 ;
   RECT 61.250 0.050 61.350 0.570 ;
  LAYER VIA2 ;
   RECT 72.050 0.050 72.150 0.570 ;
  LAYER VIA2 ;
   RECT 73.450 0.050 73.550 0.570 ;
  LAYER VIA2 ;
   RECT 77.450 0.050 77.550 0.570 ;
  LAYER VIA2 ;
   RECT 78.850 0.050 78.950 0.570 ;
  LAYER VIA2 ;
   RECT 88.850 0.050 88.950 0.570 ;
  LAYER VIA2 ;
   RECT 90.250 0.050 90.350 0.570 ;
  LAYER VIA2 ;
   RECT 94.250 0.050 94.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.650 0.050 95.750 0.570 ;
  LAYER VIA2 ;
   RECT 101.450 0.050 101.550 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 103.150 37.950 ;
  LAYER M4 ;
   RECT 0.050 0.050 103.150 40.825 ;
 END
END ST_SPHDL_128x8m8_L

MACRO ST_SPHDL_352x12m8_L
 CLASS BLOCK ;
   SIZE 136.800 BY 53.200 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 64.250 0.050 64.350 0.570 ;
   LAYER M3 ;
    RECT 64.250 0.050 64.350 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 64.850 0.050 64.950 0.570 ;
   LAYER M3 ;
    RECT 64.850 0.050 64.950 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 65.450 0.050 65.550 0.570 ;
   LAYER M3 ;
    RECT 65.450 0.050 65.550 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 71.850 0.050 71.950 0.570 ;
   LAYER M3 ;
    RECT 71.850 0.050 71.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 72.450 0.050 72.550 0.570 ;
   LAYER M3 ;
    RECT 72.450 0.050 72.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 66.250 0.050 66.350 0.570 ;
   LAYER M3 ;
    RECT 66.250 0.050 66.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 67.850 0.050 67.950 0.570 ;
   LAYER M3 ;
    RECT 67.850 0.050 67.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN A[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 62.050 0.050 62.150 0.570 ;
   LAYER M3 ;
    RECT 62.050 0.050 62.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.916 LAYER M2 ;
  ANTENNAMAXAREACAR 13.057 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.347 LAYER M3 ;
 END A[7]
 PIN A[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 63.450 0.050 63.550 0.570 ;
   LAYER M3 ;
    RECT 63.450 0.050 63.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.924 LAYER M2 ;
  ANTENNAMAXAREACAR 13.892 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.282 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.376 LAYER M3 ;
 END A[8]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 76.650 0.050 76.750 0.570 ;
   LAYER M3 ;
    RECT 76.650 0.050 76.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 78.050 0.050 78.150 0.570 ;
   LAYER M3 ;
    RECT 78.050 0.050 78.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 123.850 0.050 123.950 0.570 ;
   LAYER M3 ;
    RECT 123.850 0.050 123.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[10]
 PIN D[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 127.850 0.050 127.950 0.570 ;
   LAYER M3 ;
    RECT 127.850 0.050 127.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[11]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 40.850 0.050 40.950 0.570 ;
   LAYER M3 ;
    RECT 40.850 0.050 40.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 45.050 0.050 45.150 0.570 ;
   LAYER M3 ;
    RECT 45.050 0.050 45.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 90.250 0.050 90.350 0.570 ;
   LAYER M3 ;
    RECT 90.250 0.050 90.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 94.250 0.050 94.350 0.570 ;
   LAYER M3 ;
    RECT 94.250 0.050 94.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN D[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 107.050 0.050 107.150 0.570 ;
   LAYER M3 ;
    RECT 107.050 0.050 107.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[8]
 PIN D[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 111.050 0.050 111.150 0.570 ;
   LAYER M3 ;
    RECT 111.050 0.050 111.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[9]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[10]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 122.450 0.050 122.550 0.570 ;
   LAYER M3 ;
    RECT 122.450 0.050 122.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[10]
 PIN Q[11]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 129.250 0.050 129.350 0.570 ;
   LAYER M3 ;
    RECT 129.250 0.050 129.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[11]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 39.450 0.050 39.550 0.570 ;
   LAYER M3 ;
    RECT 39.450 0.050 39.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 46.450 0.050 46.550 0.570 ;
   LAYER M3 ;
    RECT 46.450 0.050 46.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 88.850 0.050 88.950 0.570 ;
   LAYER M3 ;
    RECT 88.850 0.050 88.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 95.650 0.050 95.750 0.570 ;
   LAYER M3 ;
    RECT 95.650 0.050 95.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN Q[8]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 105.650 0.050 105.750 0.570 ;
   LAYER M3 ;
    RECT 105.650 0.050 105.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[8]
 PIN Q[9]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 112.450 0.050 112.550 0.570 ;
   LAYER M3 ;
    RECT 112.450 0.050 112.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[9]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 135.050 0.050 135.150 0.570 ;
   LAYER M3 ;
    RECT 135.050 0.050 135.150 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 77.250 0.050 77.350 0.570 ;
   LAYER M3 ;
    RECT 77.250 0.050 77.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 69.250 0.050 69.350 0.570 ;
   LAYER M3 ;
    RECT 69.250 0.050 69.350 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 0.495 1.725 135.920 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 135.920 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 135.920 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 135.920 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 135.920 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 135.920 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 135.920 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 135.920 23.605 ;
   LAYER M4 ;
    RECT 134.535 25.290 134.915 52.355 ;
   LAYER M4 ;
    RECT 133.495 25.290 134.195 52.355 ;
   LAYER M4 ;
    RECT 131.395 25.290 132.095 52.355 ;
   LAYER M4 ;
    RECT 129.295 25.290 129.995 52.355 ;
   LAYER M4 ;
    RECT 127.195 25.290 127.895 52.355 ;
   LAYER M4 ;
    RECT 125.095 25.290 125.795 52.355 ;
   LAYER M4 ;
    RECT 124.045 25.400 124.745 52.355 ;
   LAYER M4 ;
    RECT 122.995 25.290 123.695 52.355 ;
   LAYER M4 ;
    RECT 120.895 25.290 121.595 52.355 ;
   LAYER M4 ;
    RECT 118.795 25.290 119.495 52.355 ;
   LAYER M4 ;
    RECT 116.695 25.290 117.395 52.355 ;
   LAYER M4 ;
    RECT 114.595 25.290 115.295 52.355 ;
   LAYER M4 ;
    RECT 112.495 25.290 113.195 52.355 ;
   LAYER M4 ;
    RECT 110.395 25.290 111.095 52.355 ;
   LAYER M4 ;
    RECT 108.295 25.290 108.995 52.355 ;
   LAYER M4 ;
    RECT 107.245 25.400 107.945 52.355 ;
   LAYER M4 ;
    RECT 106.195 25.290 106.895 52.355 ;
   LAYER M4 ;
    RECT 104.095 25.290 104.795 52.355 ;
   LAYER M4 ;
    RECT 101.995 25.290 102.695 52.355 ;
   LAYER M4 ;
    RECT 99.895 25.290 100.595 52.355 ;
   LAYER M4 ;
    RECT 97.795 25.290 98.495 52.355 ;
   LAYER M4 ;
    RECT 95.695 25.290 96.395 52.355 ;
   LAYER M4 ;
    RECT 93.595 25.290 94.295 52.355 ;
   LAYER M4 ;
    RECT 91.495 25.290 92.195 52.355 ;
   LAYER M4 ;
    RECT 90.445 25.400 91.145 52.355 ;
   LAYER M4 ;
    RECT 89.395 25.290 90.095 52.355 ;
   LAYER M4 ;
    RECT 87.295 25.290 87.995 52.355 ;
   LAYER M4 ;
    RECT 85.195 25.290 85.895 52.355 ;
   LAYER M4 ;
    RECT 83.095 25.360 83.795 52.355 ;
   LAYER M4 ;
    RECT 80.995 25.360 81.695 52.355 ;
   LAYER M4 ;
    RECT 79.310 25.360 79.690 52.355 ;
   LAYER M4 ;
    RECT 76.815 25.360 77.215 52.355 ;
   LAYER M4 ;
    RECT 75.345 25.360 75.845 52.355 ;
   LAYER M4 ;
    RECT 73.295 25.360 74.355 52.355 ;
   LAYER M4 ;
    RECT 70.390 25.360 70.790 52.355 ;
   LAYER M4 ;
    RECT 67.745 25.360 68.345 52.355 ;
   LAYER M4 ;
    RECT 66.075 25.360 66.720 52.355 ;
   LAYER M4 ;
    RECT 62.820 25.360 63.620 52.355 ;
   LAYER M4 ;
    RECT 61.825 25.360 62.225 52.355 ;
   LAYER M4 ;
    RECT 60.220 25.360 60.620 52.355 ;
   LAYER M4 ;
    RECT 58.005 25.360 58.810 52.355 ;
   LAYER M4 ;
    RECT 56.695 25.360 57.495 52.355 ;
   LAYER M4 ;
    RECT 54.275 25.360 54.895 52.355 ;
   LAYER M4 ;
    RECT 51.990 25.360 52.630 52.355 ;
   LAYER M4 ;
    RECT 50.555 25.290 51.255 52.355 ;
   LAYER M4 ;
    RECT 48.455 25.290 49.155 52.355 ;
   LAYER M4 ;
    RECT 46.355 25.290 47.055 52.355 ;
   LAYER M4 ;
    RECT 44.255 25.290 44.955 52.355 ;
   LAYER M4 ;
    RECT 42.155 25.290 42.855 52.355 ;
   LAYER M4 ;
    RECT 41.105 25.400 41.805 52.355 ;
   LAYER M4 ;
    RECT 40.055 25.290 40.755 52.355 ;
   LAYER M4 ;
    RECT 37.955 25.290 38.655 52.355 ;
   LAYER M4 ;
    RECT 35.855 25.290 36.555 52.355 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 52.355 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 52.355 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 52.355 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 52.355 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 52.355 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 52.355 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 52.355 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 52.355 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 52.355 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 52.355 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 52.355 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 52.355 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 52.355 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 52.355 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 52.355 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 52.355 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 52.355 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 52.355 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 52.355 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 0.495 0.760 135.920 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 135.920 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 135.920 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 135.920 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 135.920 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 135.920 11.960 ;
   LAYER M4 ;
    RECT 0.495 14.840 135.920 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 135.920 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 135.920 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 135.920 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 135.920 25.115 ;
   LAYER M4 ;
    RECT 132.445 25.290 133.145 52.355 ;
   LAYER M4 ;
    RECT 130.345 25.290 131.045 52.355 ;
   LAYER M4 ;
    RECT 128.245 25.290 128.945 52.355 ;
   LAYER M4 ;
    RECT 126.145 25.400 126.845 52.355 ;
   LAYER M4 ;
    RECT 121.945 25.290 122.645 52.355 ;
   LAYER M4 ;
    RECT 119.845 25.290 120.545 52.355 ;
   LAYER M4 ;
    RECT 117.745 25.290 118.445 52.355 ;
   LAYER M4 ;
    RECT 115.645 25.290 116.345 52.355 ;
   LAYER M4 ;
    RECT 113.545 25.290 114.245 52.355 ;
   LAYER M4 ;
    RECT 111.445 25.290 112.145 52.355 ;
   LAYER M4 ;
    RECT 109.345 25.400 110.045 52.355 ;
   LAYER M4 ;
    RECT 105.145 25.290 105.845 52.355 ;
   LAYER M4 ;
    RECT 103.045 25.290 103.745 52.355 ;
   LAYER M4 ;
    RECT 100.945 25.290 101.645 52.355 ;
   LAYER M4 ;
    RECT 98.845 25.290 99.545 52.355 ;
   LAYER M4 ;
    RECT 96.745 25.290 97.445 52.355 ;
   LAYER M4 ;
    RECT 94.645 25.290 95.345 52.355 ;
   LAYER M4 ;
    RECT 92.545 25.400 93.245 52.355 ;
   LAYER M4 ;
    RECT 88.345 25.290 89.045 52.355 ;
   LAYER M4 ;
    RECT 86.245 25.290 86.945 52.355 ;
   LAYER M4 ;
    RECT 84.145 25.290 84.845 52.355 ;
   LAYER M4 ;
    RECT 82.045 25.360 82.745 52.355 ;
   LAYER M4 ;
    RECT 79.945 25.360 80.645 52.355 ;
   LAYER M4 ;
    RECT 78.735 25.360 79.115 52.355 ;
   LAYER M4 ;
    RECT 77.530 25.360 78.510 52.355 ;
   LAYER M4 ;
    RECT 76.100 25.360 76.500 52.355 ;
   LAYER M4 ;
    RECT 74.605 25.360 75.105 52.355 ;
   LAYER M4 ;
    RECT 71.745 25.360 72.805 52.355 ;
   LAYER M4 ;
    RECT 71.065 25.360 71.465 52.355 ;
   LAYER M4 ;
    RECT 69.050 25.360 70.110 52.355 ;
   LAYER M4 ;
    RECT 67.035 25.360 67.435 52.355 ;
   LAYER M4 ;
    RECT 64.370 25.360 65.325 52.355 ;
   LAYER M4 ;
    RECT 60.910 25.360 61.550 52.355 ;
   LAYER M4 ;
    RECT 59.310 25.360 59.900 52.355 ;
   LAYER M4 ;
    RECT 55.395 25.360 56.195 52.355 ;
   LAYER M4 ;
    RECT 53.130 25.360 53.770 52.355 ;
   LAYER M4 ;
    RECT 49.505 25.290 50.205 52.355 ;
   LAYER M4 ;
    RECT 47.405 25.290 48.105 52.355 ;
   LAYER M4 ;
    RECT 45.305 25.290 46.005 52.355 ;
   LAYER M4 ;
    RECT 43.205 25.400 43.905 52.355 ;
   LAYER M4 ;
    RECT 39.005 25.290 39.705 52.355 ;
   LAYER M4 ;
    RECT 36.905 25.290 37.605 52.355 ;
   LAYER M4 ;
    RECT 34.805 25.290 35.505 52.355 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 52.355 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 52.355 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 52.355 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 52.355 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 52.355 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 52.355 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 52.355 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 52.355 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 52.355 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 52.355 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 52.355 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 52.355 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 52.355 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 52.355 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 136.750 53.150 ;
  LAYER M2 ;
   RECT 0.050 0.050 136.750 53.150 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 39.450 0.050 39.550 0.570 ;
  LAYER VIA2 ;
   RECT 40.850 0.050 40.950 0.570 ;
  LAYER VIA2 ;
   RECT 45.050 0.050 45.150 0.570 ;
  LAYER VIA2 ;
   RECT 46.450 0.050 46.550 0.570 ;
  LAYER VIA2 ;
   RECT 62.050 0.050 62.150 0.570 ;
  LAYER VIA2 ;
   RECT 63.450 0.050 63.550 0.570 ;
  LAYER VIA2 ;
   RECT 64.250 0.050 64.350 0.570 ;
  LAYER VIA2 ;
   RECT 64.850 0.050 64.950 0.570 ;
  LAYER VIA2 ;
   RECT 65.450 0.050 65.550 0.570 ;
  LAYER VIA2 ;
   RECT 66.250 0.050 66.350 0.570 ;
  LAYER VIA2 ;
   RECT 67.850 0.050 67.950 0.570 ;
  LAYER VIA2 ;
   RECT 69.250 0.050 69.350 0.570 ;
  LAYER VIA2 ;
   RECT 71.850 0.050 71.950 0.570 ;
  LAYER VIA2 ;
   RECT 72.450 0.050 72.550 0.570 ;
  LAYER VIA2 ;
   RECT 76.650 0.050 76.750 0.570 ;
  LAYER VIA2 ;
   RECT 77.250 0.050 77.350 0.570 ;
  LAYER VIA2 ;
   RECT 78.050 0.050 78.150 0.570 ;
  LAYER VIA2 ;
   RECT 88.850 0.050 88.950 0.570 ;
  LAYER VIA2 ;
   RECT 90.250 0.050 90.350 0.570 ;
  LAYER VIA2 ;
   RECT 94.250 0.050 94.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.650 0.050 95.750 0.570 ;
  LAYER VIA2 ;
   RECT 105.650 0.050 105.750 0.570 ;
  LAYER VIA2 ;
   RECT 107.050 0.050 107.150 0.570 ;
  LAYER VIA2 ;
   RECT 111.050 0.050 111.150 0.570 ;
  LAYER VIA2 ;
   RECT 112.450 0.050 112.550 0.570 ;
  LAYER VIA2 ;
   RECT 122.450 0.050 122.550 0.570 ;
  LAYER VIA2 ;
   RECT 123.850 0.050 123.950 0.570 ;
  LAYER VIA2 ;
   RECT 127.850 0.050 127.950 0.570 ;
  LAYER VIA2 ;
   RECT 129.250 0.050 129.350 0.570 ;
  LAYER VIA2 ;
   RECT 135.050 0.050 135.150 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 136.750 53.150 ;
  LAYER M4 ;
   RECT 0.050 0.050 136.750 53.150 ;
 END
END ST_SPHDL_352x12m8_L

MACRO ST_SPHDL_4096x32m8_L
 CLASS BLOCK ;
   SIZE 304.800 BY 311.800 ;
 SYMMETRY R90 X Y ;
 PIN A[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.250 0.050 148.350 0.570 ;
   LAYER M3 ;
    RECT 148.250 0.050 148.350 0.570 ;
  END
  ANTENNADIFFAREA 0.066 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 7.871 LAYER M2 ;
  ANTENNAMAXAREACAR 12.314 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.575 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.013 LAYER M3 ;
 END A[0]
 PIN A[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 143.650 0.050 143.750 0.570 ;
   LAYER M3 ;
    RECT 143.650 0.050 143.750 0.570 ;
  END
  ANTENNADIFFAREA 0.090 LAYER M3 ;
  ANTENNAGATEAREA 0.252 LAYER M2 ;
  ANTENNAGATEAREA 0.252 LAYER M3 ;
  ANTENNAMAXAREACAR 0.941 LAYER M2 ;
  ANTENNAMAXAREACAR 6.310 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.301 LAYER M3 ;
 END A[10]
 PIN A[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 136.650 0.050 136.750 0.570 ;
   LAYER M3 ;
    RECT 136.650 0.050 136.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.251 LAYER M2 ;
  ANTENNAGATEAREA 0.251 LAYER M3 ;
  ANTENNAMAXAREACAR 0.362 LAYER M2 ;
  ANTENNAMAXAREACAR 5.727 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.297 LAYER M3 ;
 END A[11]
 PIN A[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 148.850 0.050 148.950 0.570 ;
   LAYER M3 ;
    RECT 148.850 0.050 148.950 0.570 ;
  END
  ANTENNADIFFAREA 0.067 LAYER M3 ;
  ANTENNAGATEAREA 0.084 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 2.374 LAYER M2 ;
  ANTENNAMAXAREACAR 7.059 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.068 LAYER M3 ;
 END A[1]
 PIN A[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 149.450 0.050 149.550 0.570 ;
   LAYER M3 ;
    RECT 149.450 0.050 149.550 0.570 ;
  END
  ANTENNADIFFAREA 0.065 LAYER M3 ;
  ANTENNAGATEAREA 0.228 LAYER M2 ;
  ANTENNAGATEAREA 0.228 LAYER M3 ;
  ANTENNAMAXAREACAR 0.451 LAYER M2 ;
  ANTENNAMAXAREACAR 4.045 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.767 LAYER M3 ;
 END A[2]
 PIN A[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 155.850 0.050 155.950 0.570 ;
   LAYER M3 ;
    RECT 155.850 0.050 155.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.100 LAYER M2 ;
  ANTENNAMAXAREACAR 13.652 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.404 LAYER M3 ;
 END A[3]
 PIN A[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 156.450 0.050 156.550 0.570 ;
   LAYER M3 ;
    RECT 156.450 0.050 156.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.066 LAYER M2 ;
  ANTENNAMAXAREACAR 12.811 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.219 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.345 LAYER M3 ;
 END A[4]
 PIN A[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 150.250 0.050 150.350 0.570 ;
   LAYER M3 ;
    RECT 150.250 0.050 150.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.864 LAYER M2 ;
  ANTENNAMAXAREACAR 14.205 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.513 LAYER M3 ;
 END A[5]
 PIN A[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 151.850 0.050 151.950 0.570 ;
   LAYER M3 ;
    RECT 151.850 0.050 151.950 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 5.158 LAYER M2 ;
  ANTENNAMAXAREACAR 15.799 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.350 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.468 LAYER M3 ;
 END A[6]
 PIN A[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 146.050 0.050 146.150 0.570 ;
   LAYER M3 ;
    RECT 146.050 0.050 146.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 2.916 LAYER M2 ;
  ANTENNAMAXAREACAR 13.057 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.347 LAYER M3 ;
 END A[7]
 PIN A[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 147.450 0.050 147.550 0.570 ;
   LAYER M3 ;
    RECT 147.450 0.050 147.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.138 LAYER M2 ;
  ANTENNAGATEAREA 0.138 LAYER M3 ;
  ANTENNAMAXAREACAR 3.924 LAYER M2 ;
  ANTENNAMAXAREACAR 13.892 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.282 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.376 LAYER M3 ;
 END A[8]
 PIN A[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 137.450 0.050 137.550 0.570 ;
   LAYER M3 ;
    RECT 137.450 0.050 137.550 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.251 LAYER M2 ;
  ANTENNAGATEAREA 0.251 LAYER M3 ;
  ANTENNAMAXAREACAR 3.203 LAYER M2 ;
  ANTENNAMAXAREACAR 9.213 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.586 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.511 LAYER M3 ;
 END A[9]
 PIN CK
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 160.650 0.050 160.750 0.570 ;
   LAYER M3 ;
    RECT 160.650 0.050 160.750 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.480 LAYER M2 ;
  ANTENNAGATEAREA 1.256 LAYER M3 ;
  ANTENNAMAXAREACAR 1.206 LAYER M2 ;
  ANTENNAMAXAREACAR 2.600 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.687 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.750 LAYER M3 ;
 END CK
 PIN CSN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 162.050 0.050 162.150 0.570 ;
   LAYER M3 ;
    RECT 162.050 0.050 162.150 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.060 LAYER M2 ;
  ANTENNAGATEAREA 0.060 LAYER M3 ;
  ANTENNAMAXAREACAR 2.470 LAYER M2 ;
  ANTENNAMAXAREACAR 26.441 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.386 LAYER M3 ;
 END CSN
 PIN D[0]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 7.250 0.050 7.350 0.570 ;
   LAYER M3 ;
    RECT 7.250 0.050 7.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[0]
 PIN D[10]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 91.250 0.050 91.350 0.570 ;
   LAYER M3 ;
    RECT 91.250 0.050 91.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[10]
 PIN D[11]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 95.450 0.050 95.550 0.570 ;
   LAYER M3 ;
    RECT 95.450 0.050 95.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[11]
 PIN D[12]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 108.050 0.050 108.150 0.570 ;
   LAYER M3 ;
    RECT 108.050 0.050 108.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[12]
 PIN D[13]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 112.250 0.050 112.350 0.570 ;
   LAYER M3 ;
    RECT 112.250 0.050 112.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[13]
 PIN D[14]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 124.850 0.050 124.950 0.570 ;
   LAYER M3 ;
    RECT 124.850 0.050 124.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[14]
 PIN D[15]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 129.050 0.050 129.150 0.570 ;
   LAYER M3 ;
    RECT 129.050 0.050 129.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[15]
 PIN D[16]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 174.250 0.050 174.350 0.570 ;
   LAYER M3 ;
    RECT 174.250 0.050 174.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[16]
 PIN D[17]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 178.250 0.050 178.350 0.570 ;
   LAYER M3 ;
    RECT 178.250 0.050 178.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[17]
 PIN D[18]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 191.050 0.050 191.150 0.570 ;
   LAYER M3 ;
    RECT 191.050 0.050 191.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[18]
 PIN D[19]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 195.050 0.050 195.150 0.570 ;
   LAYER M3 ;
    RECT 195.050 0.050 195.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[19]
 PIN D[1]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 11.450 0.050 11.550 0.570 ;
   LAYER M3 ;
    RECT 11.450 0.050 11.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[1]
 PIN D[20]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 207.850 0.050 207.950 0.570 ;
   LAYER M3 ;
    RECT 207.850 0.050 207.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[20]
 PIN D[21]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 211.850 0.050 211.950 0.570 ;
   LAYER M3 ;
    RECT 211.850 0.050 211.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[21]
 PIN D[22]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 224.650 0.050 224.750 0.570 ;
   LAYER M3 ;
    RECT 224.650 0.050 224.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[22]
 PIN D[23]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 228.650 0.050 228.750 0.570 ;
   LAYER M3 ;
    RECT 228.650 0.050 228.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[23]
 PIN D[24]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 241.450 0.050 241.550 0.570 ;
   LAYER M3 ;
    RECT 241.450 0.050 241.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[24]
 PIN D[25]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 245.450 0.050 245.550 0.570 ;
   LAYER M3 ;
    RECT 245.450 0.050 245.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[25]
 PIN D[26]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 258.250 0.050 258.350 0.570 ;
   LAYER M3 ;
    RECT 258.250 0.050 258.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[26]
 PIN D[27]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 262.250 0.050 262.350 0.570 ;
   LAYER M3 ;
    RECT 262.250 0.050 262.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[27]
 PIN D[28]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 275.050 0.050 275.150 0.570 ;
   LAYER M3 ;
    RECT 275.050 0.050 275.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[28]
 PIN D[29]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 279.050 0.050 279.150 0.570 ;
   LAYER M3 ;
    RECT 279.050 0.050 279.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[29]
 PIN D[2]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 24.050 0.050 24.150 0.570 ;
   LAYER M3 ;
    RECT 24.050 0.050 24.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[2]
 PIN D[30]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 291.850 0.050 291.950 0.570 ;
   LAYER M3 ;
    RECT 291.850 0.050 291.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[30]
 PIN D[31]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 295.850 0.050 295.950 0.570 ;
   LAYER M3 ;
    RECT 295.850 0.050 295.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[31]
 PIN D[3]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 28.250 0.050 28.350 0.570 ;
   LAYER M3 ;
    RECT 28.250 0.050 28.350 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[3]
 PIN D[4]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 40.850 0.050 40.950 0.570 ;
   LAYER M3 ;
    RECT 40.850 0.050 40.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[4]
 PIN D[5]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 45.050 0.050 45.150 0.570 ;
   LAYER M3 ;
    RECT 45.050 0.050 45.150 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[5]
 PIN D[6]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 57.650 0.050 57.750 0.570 ;
   LAYER M3 ;
    RECT 57.650 0.050 57.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[6]
 PIN D[7]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 61.850 0.050 61.950 0.570 ;
   LAYER M3 ;
    RECT 61.850 0.050 61.950 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[7]
 PIN D[8]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 74.450 0.050 74.550 0.570 ;
   LAYER M3 ;
    RECT 74.450 0.050 74.550 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[8]
 PIN D[9]
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 78.650 0.050 78.750 0.570 ;
   LAYER M3 ;
    RECT 78.650 0.050 78.750 0.570 ;
  END
  ANTENNADIFFAREA 0.076 LAYER M2 ;
  ANTENNADIFFAREA 0.076 LAYER M3 ;
  ANTENNAGATEAREA 0.027 LAYER M2 ;
  ANTENNAGATEAREA 0.027 LAYER M3 ;
  ANTENNAMAXAREACAR 13.119 LAYER M2 ;
  ANTENNAMAXAREACAR 20.819 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.020 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.298 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.156 LAYER M3 ;
 END D[9]
 PIN Q[0]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 5.850 0.050 5.950 0.570 ;
   LAYER M3 ;
    RECT 5.850 0.050 5.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[0]
 PIN Q[10]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 89.850 0.050 89.950 0.570 ;
   LAYER M3 ;
    RECT 89.850 0.050 89.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[10]
 PIN Q[11]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 96.850 0.050 96.950 0.570 ;
   LAYER M3 ;
    RECT 96.850 0.050 96.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[11]
 PIN Q[12]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 106.650 0.050 106.750 0.570 ;
   LAYER M3 ;
    RECT 106.650 0.050 106.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[12]
 PIN Q[13]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 113.650 0.050 113.750 0.570 ;
   LAYER M3 ;
    RECT 113.650 0.050 113.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[13]
 PIN Q[14]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 123.450 0.050 123.550 0.570 ;
   LAYER M3 ;
    RECT 123.450 0.050 123.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[14]
 PIN Q[15]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 130.450 0.050 130.550 0.570 ;
   LAYER M3 ;
    RECT 130.450 0.050 130.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[15]
 PIN Q[16]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 172.850 0.050 172.950 0.570 ;
   LAYER M3 ;
    RECT 172.850 0.050 172.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[16]
 PIN Q[17]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 179.650 0.050 179.750 0.570 ;
   LAYER M3 ;
    RECT 179.650 0.050 179.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[17]
 PIN Q[18]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 189.650 0.050 189.750 0.570 ;
   LAYER M3 ;
    RECT 189.650 0.050 189.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[18]
 PIN Q[19]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 196.450 0.050 196.550 0.570 ;
   LAYER M3 ;
    RECT 196.450 0.050 196.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[19]
 PIN Q[1]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 12.850 0.050 12.950 0.570 ;
   LAYER M3 ;
    RECT 12.850 0.050 12.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[1]
 PIN Q[20]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 206.450 0.050 206.550 0.570 ;
   LAYER M3 ;
    RECT 206.450 0.050 206.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[20]
 PIN Q[21]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 213.250 0.050 213.350 0.570 ;
   LAYER M3 ;
    RECT 213.250 0.050 213.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[21]
 PIN Q[22]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 223.250 0.050 223.350 0.570 ;
   LAYER M3 ;
    RECT 223.250 0.050 223.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[22]
 PIN Q[23]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 230.050 0.050 230.150 0.570 ;
   LAYER M3 ;
    RECT 230.050 0.050 230.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[23]
 PIN Q[24]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 240.050 0.050 240.150 0.570 ;
   LAYER M3 ;
    RECT 240.050 0.050 240.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[24]
 PIN Q[25]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 246.850 0.050 246.950 0.570 ;
   LAYER M3 ;
    RECT 246.850 0.050 246.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[25]
 PIN Q[26]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 256.850 0.050 256.950 0.570 ;
   LAYER M3 ;
    RECT 256.850 0.050 256.950 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[26]
 PIN Q[27]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 263.650 0.050 263.750 0.570 ;
   LAYER M3 ;
    RECT 263.650 0.050 263.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[27]
 PIN Q[28]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 273.650 0.050 273.750 0.570 ;
   LAYER M3 ;
    RECT 273.650 0.050 273.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[28]
 PIN Q[29]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 280.450 0.050 280.550 0.570 ;
   LAYER M3 ;
    RECT 280.450 0.050 280.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[29]
 PIN Q[2]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 22.650 0.050 22.750 0.570 ;
   LAYER M3 ;
    RECT 22.650 0.050 22.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[2]
 PIN Q[30]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 290.450 0.050 290.550 0.570 ;
   LAYER M3 ;
    RECT 290.450 0.050 290.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[30]
 PIN Q[31]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 297.250 0.050 297.350 0.570 ;
   LAYER M3 ;
    RECT 297.250 0.050 297.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[31]
 PIN Q[3]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 29.650 0.050 29.750 0.570 ;
   LAYER M3 ;
    RECT 29.650 0.050 29.750 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[3]
 PIN Q[4]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 39.450 0.050 39.550 0.570 ;
   LAYER M3 ;
    RECT 39.450 0.050 39.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[4]
 PIN Q[5]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 46.450 0.050 46.550 0.570 ;
   LAYER M3 ;
    RECT 46.450 0.050 46.550 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[5]
 PIN Q[6]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 56.250 0.050 56.350 0.570 ;
   LAYER M3 ;
    RECT 56.250 0.050 56.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[6]
 PIN Q[7]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 63.250 0.050 63.350 0.570 ;
   LAYER M3 ;
    RECT 63.250 0.050 63.350 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[7]
 PIN Q[8]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 73.050 0.050 73.150 0.570 ;
   LAYER M3 ;
    RECT 73.050 0.050 73.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[8]
 PIN Q[9]
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 80.050 0.050 80.150 0.570 ;
   LAYER M3 ;
    RECT 80.050 0.050 80.150 0.570 ;
  END
  ANTENNADIFFAREA 1.039 LAYER M2 ;
  ANTENNADIFFAREA 1.039 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.030 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.160 LAYER M3 ;
 END Q[9]
 PIN RY
  DIRECTION OUTPUT ;
  PORT
   LAYER M2 ;
    RECT 303.050 0.050 303.150 0.570 ;
   LAYER M3 ;
    RECT 303.050 0.050 303.150 0.570 ;
  END
  ANTENNADIFFAREA 1.191 LAYER M2 ;
  ANTENNADIFFAREA 1.191 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 1.238 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.179 LAYER M3 ;
 END RY
 PIN TBYPASS
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 161.250 0.050 161.350 0.570 ;
   LAYER M3 ;
    RECT 161.250 0.050 161.350 0.570 ;
  END
  ANTENNADIFFAREA 0.060 LAYER M3 ;
  ANTENNAGATEAREA 0.042 LAYER M2 ;
  ANTENNAGATEAREA 0.102 LAYER M3 ;
  ANTENNAMAXAREACAR 19.706 LAYER M2 ;
  ANTENNAMAXAREACAR 32.634 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.747 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 1.319 LAYER M3 ;
 END TBYPASS
 PIN WEN
  DIRECTION INPUT ;
  PORT
   LAYER M2 ;
    RECT 153.250 0.050 153.350 0.570 ;
   LAYER M3 ;
    RECT 153.250 0.050 153.350 0.570 ;
  END
  ANTENNADIFFAREA 0.070 LAYER M3 ;
  ANTENNAGATEAREA 0.036 LAYER M2 ;
  ANTENNAGATEAREA 0.036 LAYER M3 ;
  ANTENNAMAXAREACAR 6.497 LAYER M2 ;
  ANTENNAMAXAREACAR 26.803 LAYER M3 ;
  ANTENNAPARTIALCUTAREA 0.040 LAYER VIA2 ;
  ANTENNAPARTIALMETALAREA 0.163 LAYER M2 ;
  ANTENNAPARTIALMETALAREA 0.679 LAYER M3 ;
 END WEN
 PIN gnd
  DIRECTION INOUT ;
  USE GROUND ;
  PORT
   LAYER M4 ;
    RECT 128.255 25.290 128.955 311.095 ;
   LAYER M4 ;
    RECT 126.155 25.290 126.855 311.095 ;
   LAYER M4 ;
    RECT 125.105 25.400 125.805 311.095 ;
   LAYER M4 ;
    RECT 124.055 25.290 124.755 311.095 ;
   LAYER M4 ;
    RECT 121.955 25.290 122.655 311.095 ;
   LAYER M4 ;
    RECT 119.855 25.290 120.555 311.095 ;
   LAYER M4 ;
    RECT 117.755 25.290 118.455 311.095 ;
   LAYER M4 ;
    RECT 115.655 25.290 116.355 311.095 ;
   LAYER M4 ;
    RECT 113.555 25.290 114.255 311.095 ;
   LAYER M4 ;
    RECT 111.455 25.290 112.155 311.095 ;
   LAYER M4 ;
    RECT 109.355 25.290 110.055 311.095 ;
   LAYER M4 ;
    RECT 108.305 25.400 109.005 311.095 ;
   LAYER M4 ;
    RECT 107.255 25.290 107.955 311.095 ;
   LAYER M4 ;
    RECT 105.155 25.290 105.855 311.095 ;
   LAYER M4 ;
    RECT 103.055 25.290 103.755 311.095 ;
   LAYER M4 ;
    RECT 100.955 25.290 101.655 311.095 ;
   LAYER M4 ;
    RECT 98.855 25.290 99.555 311.095 ;
   LAYER M4 ;
    RECT 96.755 25.290 97.455 311.095 ;
   LAYER M4 ;
    RECT 94.655 25.290 95.355 311.095 ;
   LAYER M4 ;
    RECT 92.555 25.290 93.255 311.095 ;
   LAYER M4 ;
    RECT 91.505 25.400 92.205 311.095 ;
   LAYER M4 ;
    RECT 90.455 25.290 91.155 311.095 ;
   LAYER M4 ;
    RECT 88.355 25.290 89.055 311.095 ;
   LAYER M4 ;
    RECT 86.255 25.290 86.955 311.095 ;
   LAYER M4 ;
    RECT 84.155 25.290 84.855 311.095 ;
   LAYER M4 ;
    RECT 82.055 25.290 82.755 311.095 ;
   LAYER M4 ;
    RECT 79.955 25.290 80.655 311.095 ;
   LAYER M4 ;
    RECT 77.855 25.290 78.555 311.095 ;
   LAYER M4 ;
    RECT 75.755 25.290 76.455 311.095 ;
   LAYER M4 ;
    RECT 74.705 25.400 75.405 311.095 ;
   LAYER M4 ;
    RECT 73.655 25.290 74.355 311.095 ;
   LAYER M4 ;
    RECT 71.555 25.290 72.255 311.095 ;
   LAYER M4 ;
    RECT 69.455 25.290 70.155 311.095 ;
   LAYER M4 ;
    RECT 67.355 25.290 68.055 311.095 ;
   LAYER M4 ;
    RECT 65.255 25.290 65.955 311.095 ;
   LAYER M4 ;
    RECT 63.155 25.290 63.855 311.095 ;
   LAYER M4 ;
    RECT 61.055 25.290 61.755 311.095 ;
   LAYER M4 ;
    RECT 58.955 25.290 59.655 311.095 ;
   LAYER M4 ;
    RECT 57.905 25.400 58.605 311.095 ;
   LAYER M4 ;
    RECT 56.855 25.290 57.555 311.095 ;
   LAYER M4 ;
    RECT 54.755 25.290 55.455 311.095 ;
   LAYER M4 ;
    RECT 52.655 25.290 53.355 311.095 ;
   LAYER M4 ;
    RECT 50.555 25.290 51.255 311.095 ;
   LAYER M4 ;
    RECT 48.455 25.290 49.155 311.095 ;
   LAYER M4 ;
    RECT 46.355 25.290 47.055 311.095 ;
   LAYER M4 ;
    RECT 44.255 25.290 44.955 311.095 ;
   LAYER M4 ;
    RECT 42.155 25.290 42.855 311.095 ;
   LAYER M4 ;
    RECT 41.105 25.400 41.805 311.095 ;
   LAYER M4 ;
    RECT 40.055 25.290 40.755 311.095 ;
   LAYER M4 ;
    RECT 37.955 25.290 38.655 311.095 ;
   LAYER M4 ;
    RECT 35.855 25.290 36.555 311.095 ;
   LAYER M4 ;
    RECT 33.755 25.290 34.455 311.095 ;
   LAYER M4 ;
    RECT 31.655 25.290 32.355 311.095 ;
   LAYER M4 ;
    RECT 29.555 25.290 30.255 311.095 ;
   LAYER M4 ;
    RECT 27.455 25.290 28.155 311.095 ;
   LAYER M4 ;
    RECT 25.355 25.290 26.055 311.095 ;
   LAYER M4 ;
    RECT 24.305 25.400 25.005 311.095 ;
   LAYER M4 ;
    RECT 23.255 25.290 23.955 311.095 ;
   LAYER M4 ;
    RECT 21.155 25.290 21.855 311.095 ;
   LAYER M4 ;
    RECT 19.055 25.290 19.755 311.095 ;
   LAYER M4 ;
    RECT 16.955 25.290 17.655 311.095 ;
   LAYER M4 ;
    RECT 14.855 25.290 15.555 311.095 ;
   LAYER M4 ;
    RECT 12.755 25.290 13.455 311.095 ;
   LAYER M4 ;
    RECT 10.655 25.290 11.355 311.095 ;
   LAYER M4 ;
    RECT 8.555 25.290 9.255 311.095 ;
   LAYER M4 ;
    RECT 7.505 25.400 8.205 311.095 ;
   LAYER M4 ;
    RECT 6.455 25.290 7.155 311.095 ;
   LAYER M4 ;
    RECT 4.355 25.290 5.055 311.095 ;
   LAYER M4 ;
    RECT 2.255 25.290 2.955 311.095 ;
   LAYER M4 ;
    RECT 0.485 25.290 0.865 311.095 ;
   LAYER M4 ;
    RECT 0.495 1.725 303.920 2.425 ;
   LAYER M4 ;
    RECT 0.495 5.995 303.920 6.375 ;
   LAYER M4 ;
    RECT 0.495 7.305 303.920 8.555 ;
   LAYER M4 ;
    RECT 0.495 10.120 303.920 11.020 ;
   LAYER M4 ;
    RECT 0.495 15.420 303.920 16.660 ;
   LAYER M4 ;
    RECT 0.495 19.075 303.920 19.775 ;
   LAYER M4 ;
    RECT 0.495 20.805 303.920 21.225 ;
   LAYER M4 ;
    RECT 0.495 22.595 303.920 23.605 ;
   LAYER M4 ;
    RECT 302.535 25.290 302.915 311.095 ;
   LAYER M4 ;
    RECT 301.495 25.290 302.195 311.095 ;
   LAYER M4 ;
    RECT 299.395 25.290 300.095 311.095 ;
   LAYER M4 ;
    RECT 297.295 25.290 297.995 311.095 ;
   LAYER M4 ;
    RECT 295.195 25.290 295.895 311.095 ;
   LAYER M4 ;
    RECT 293.095 25.290 293.795 311.095 ;
   LAYER M4 ;
    RECT 292.045 25.400 292.745 311.095 ;
   LAYER M4 ;
    RECT 290.995 25.290 291.695 311.095 ;
   LAYER M4 ;
    RECT 288.895 25.290 289.595 311.095 ;
   LAYER M4 ;
    RECT 286.795 25.290 287.495 311.095 ;
   LAYER M4 ;
    RECT 284.695 25.290 285.395 311.095 ;
   LAYER M4 ;
    RECT 282.595 25.290 283.295 311.095 ;
   LAYER M4 ;
    RECT 280.495 25.290 281.195 311.095 ;
   LAYER M4 ;
    RECT 278.395 25.290 279.095 311.095 ;
   LAYER M4 ;
    RECT 276.295 25.290 276.995 311.095 ;
   LAYER M4 ;
    RECT 275.245 25.400 275.945 311.095 ;
   LAYER M4 ;
    RECT 274.195 25.290 274.895 311.095 ;
   LAYER M4 ;
    RECT 272.095 25.290 272.795 311.095 ;
   LAYER M4 ;
    RECT 269.995 25.290 270.695 311.095 ;
   LAYER M4 ;
    RECT 267.895 25.290 268.595 311.095 ;
   LAYER M4 ;
    RECT 265.795 25.290 266.495 311.095 ;
   LAYER M4 ;
    RECT 263.695 25.290 264.395 311.095 ;
   LAYER M4 ;
    RECT 261.595 25.290 262.295 311.095 ;
   LAYER M4 ;
    RECT 259.495 25.290 260.195 311.095 ;
   LAYER M4 ;
    RECT 258.445 25.400 259.145 311.095 ;
   LAYER M4 ;
    RECT 257.395 25.290 258.095 311.095 ;
   LAYER M4 ;
    RECT 255.295 25.290 255.995 311.095 ;
   LAYER M4 ;
    RECT 253.195 25.290 253.895 311.095 ;
   LAYER M4 ;
    RECT 251.095 25.290 251.795 311.095 ;
   LAYER M4 ;
    RECT 248.995 25.290 249.695 311.095 ;
   LAYER M4 ;
    RECT 246.895 25.290 247.595 311.095 ;
   LAYER M4 ;
    RECT 244.795 25.290 245.495 311.095 ;
   LAYER M4 ;
    RECT 242.695 25.290 243.395 311.095 ;
   LAYER M4 ;
    RECT 241.645 25.400 242.345 311.095 ;
   LAYER M4 ;
    RECT 240.595 25.290 241.295 311.095 ;
   LAYER M4 ;
    RECT 238.495 25.290 239.195 311.095 ;
   LAYER M4 ;
    RECT 236.395 25.290 237.095 311.095 ;
   LAYER M4 ;
    RECT 234.295 25.290 234.995 311.095 ;
   LAYER M4 ;
    RECT 232.195 25.290 232.895 311.095 ;
   LAYER M4 ;
    RECT 230.095 25.290 230.795 311.095 ;
   LAYER M4 ;
    RECT 227.995 25.290 228.695 311.095 ;
   LAYER M4 ;
    RECT 225.895 25.290 226.595 311.095 ;
   LAYER M4 ;
    RECT 224.845 25.400 225.545 311.095 ;
   LAYER M4 ;
    RECT 223.795 25.290 224.495 311.095 ;
   LAYER M4 ;
    RECT 221.695 25.290 222.395 311.095 ;
   LAYER M4 ;
    RECT 219.595 25.290 220.295 311.095 ;
   LAYER M4 ;
    RECT 217.495 25.290 218.195 311.095 ;
   LAYER M4 ;
    RECT 215.395 25.290 216.095 311.095 ;
   LAYER M4 ;
    RECT 213.295 25.290 213.995 311.095 ;
   LAYER M4 ;
    RECT 211.195 25.290 211.895 311.095 ;
   LAYER M4 ;
    RECT 209.095 25.290 209.795 311.095 ;
   LAYER M4 ;
    RECT 208.045 25.400 208.745 311.095 ;
   LAYER M4 ;
    RECT 206.995 25.290 207.695 311.095 ;
   LAYER M4 ;
    RECT 204.895 25.290 205.595 311.095 ;
   LAYER M4 ;
    RECT 202.795 25.290 203.495 311.095 ;
   LAYER M4 ;
    RECT 200.695 25.290 201.395 311.095 ;
   LAYER M4 ;
    RECT 198.595 25.290 199.295 311.095 ;
   LAYER M4 ;
    RECT 196.495 25.290 197.195 311.095 ;
   LAYER M4 ;
    RECT 194.395 25.290 195.095 311.095 ;
   LAYER M4 ;
    RECT 192.295 25.290 192.995 311.095 ;
   LAYER M4 ;
    RECT 191.245 25.400 191.945 311.095 ;
   LAYER M4 ;
    RECT 190.195 25.290 190.895 311.095 ;
   LAYER M4 ;
    RECT 188.095 25.290 188.795 311.095 ;
   LAYER M4 ;
    RECT 185.995 25.290 186.695 311.095 ;
   LAYER M4 ;
    RECT 183.895 25.290 184.595 311.095 ;
   LAYER M4 ;
    RECT 181.795 25.290 182.495 311.095 ;
   LAYER M4 ;
    RECT 179.695 25.290 180.395 311.095 ;
   LAYER M4 ;
    RECT 177.595 25.290 178.295 311.095 ;
   LAYER M4 ;
    RECT 175.495 25.290 176.195 311.095 ;
   LAYER M4 ;
    RECT 174.445 25.400 175.145 311.095 ;
   LAYER M4 ;
    RECT 173.395 25.290 174.095 311.095 ;
   LAYER M4 ;
    RECT 171.295 25.290 171.995 311.095 ;
   LAYER M4 ;
    RECT 169.195 25.290 169.895 311.095 ;
   LAYER M4 ;
    RECT 167.095 25.360 167.795 311.095 ;
   LAYER M4 ;
    RECT 164.995 25.360 165.695 311.095 ;
   LAYER M4 ;
    RECT 163.310 25.360 163.690 311.095 ;
   LAYER M4 ;
    RECT 160.815 25.360 161.215 311.095 ;
   LAYER M4 ;
    RECT 159.345 25.360 159.845 311.095 ;
   LAYER M4 ;
    RECT 157.295 25.360 158.355 311.095 ;
   LAYER M4 ;
    RECT 154.390 25.360 154.790 311.095 ;
   LAYER M4 ;
    RECT 151.745 25.360 152.345 311.095 ;
   LAYER M4 ;
    RECT 150.075 25.360 150.720 311.095 ;
   LAYER M4 ;
    RECT 146.820 25.360 147.620 311.095 ;
   LAYER M4 ;
    RECT 145.825 25.360 146.225 311.095 ;
   LAYER M4 ;
    RECT 144.220 25.360 144.620 311.095 ;
   LAYER M4 ;
    RECT 142.005 25.360 142.810 311.095 ;
   LAYER M4 ;
    RECT 140.695 25.360 141.495 311.095 ;
   LAYER M4 ;
    RECT 138.275 25.360 138.895 311.095 ;
   LAYER M4 ;
    RECT 135.990 25.360 136.630 311.095 ;
   LAYER M4 ;
    RECT 134.555 25.290 135.255 311.095 ;
   LAYER M4 ;
    RECT 132.455 25.290 133.155 311.095 ;
   LAYER M4 ;
    RECT 130.355 25.290 131.055 311.095 ;
  END
 END gnd
 PIN vdd
  DIRECTION INOUT ;
  USE POWER ;
  PORT
   LAYER M4 ;
    RECT 36.905 25.290 37.605 311.095 ;
   LAYER M4 ;
    RECT 34.805 25.290 35.505 311.095 ;
   LAYER M4 ;
    RECT 32.705 25.290 33.405 311.095 ;
   LAYER M4 ;
    RECT 30.605 25.290 31.305 311.095 ;
   LAYER M4 ;
    RECT 28.505 25.290 29.205 311.095 ;
   LAYER M4 ;
    RECT 26.405 25.400 27.105 311.095 ;
   LAYER M4 ;
    RECT 22.205 25.290 22.905 311.095 ;
   LAYER M4 ;
    RECT 20.105 25.290 20.805 311.095 ;
   LAYER M4 ;
    RECT 18.005 25.290 18.705 311.095 ;
   LAYER M4 ;
    RECT 15.905 25.290 16.605 311.095 ;
   LAYER M4 ;
    RECT 13.805 25.290 14.505 311.095 ;
   LAYER M4 ;
    RECT 11.705 25.290 12.405 311.095 ;
   LAYER M4 ;
    RECT 9.605 25.400 10.305 311.095 ;
   LAYER M4 ;
    RECT 5.405 25.290 6.105 311.095 ;
   LAYER M4 ;
    RECT 3.305 25.290 4.005 311.095 ;
   LAYER M4 ;
    RECT 1.205 25.290 1.905 311.095 ;
   LAYER M4 ;
    RECT 0.495 14.840 303.920 15.020 ;
   LAYER M4 ;
    RECT 0.495 17.425 303.920 18.695 ;
   LAYER M4 ;
    RECT 0.495 20.085 303.920 20.505 ;
   LAYER M4 ;
    RECT 0.495 21.550 303.920 22.250 ;
   LAYER M4 ;
    RECT 0.495 24.105 303.920 25.115 ;
   LAYER M4 ;
    RECT 300.445 25.290 301.145 311.095 ;
   LAYER M4 ;
    RECT 298.345 25.290 299.045 311.095 ;
   LAYER M4 ;
    RECT 296.245 25.290 296.945 311.095 ;
   LAYER M4 ;
    RECT 294.145 25.400 294.845 311.095 ;
   LAYER M4 ;
    RECT 289.945 25.290 290.645 311.095 ;
   LAYER M4 ;
    RECT 287.845 25.290 288.545 311.095 ;
   LAYER M4 ;
    RECT 285.745 25.290 286.445 311.095 ;
   LAYER M4 ;
    RECT 283.645 25.290 284.345 311.095 ;
   LAYER M4 ;
    RECT 281.545 25.290 282.245 311.095 ;
   LAYER M4 ;
    RECT 279.445 25.290 280.145 311.095 ;
   LAYER M4 ;
    RECT 277.345 25.400 278.045 311.095 ;
   LAYER M4 ;
    RECT 273.145 25.290 273.845 311.095 ;
   LAYER M4 ;
    RECT 271.045 25.290 271.745 311.095 ;
   LAYER M4 ;
    RECT 268.945 25.290 269.645 311.095 ;
   LAYER M4 ;
    RECT 266.845 25.290 267.545 311.095 ;
   LAYER M4 ;
    RECT 264.745 25.290 265.445 311.095 ;
   LAYER M4 ;
    RECT 262.645 25.290 263.345 311.095 ;
   LAYER M4 ;
    RECT 260.545 25.400 261.245 311.095 ;
   LAYER M4 ;
    RECT 256.345 25.290 257.045 311.095 ;
   LAYER M4 ;
    RECT 254.245 25.290 254.945 311.095 ;
   LAYER M4 ;
    RECT 252.145 25.290 252.845 311.095 ;
   LAYER M4 ;
    RECT 250.045 25.290 250.745 311.095 ;
   LAYER M4 ;
    RECT 247.945 25.290 248.645 311.095 ;
   LAYER M4 ;
    RECT 245.845 25.290 246.545 311.095 ;
   LAYER M4 ;
    RECT 243.745 25.400 244.445 311.095 ;
   LAYER M4 ;
    RECT 239.545 25.290 240.245 311.095 ;
   LAYER M4 ;
    RECT 237.445 25.290 238.145 311.095 ;
   LAYER M4 ;
    RECT 235.345 25.290 236.045 311.095 ;
   LAYER M4 ;
    RECT 233.245 25.290 233.945 311.095 ;
   LAYER M4 ;
    RECT 231.145 25.290 231.845 311.095 ;
   LAYER M4 ;
    RECT 229.045 25.290 229.745 311.095 ;
   LAYER M4 ;
    RECT 226.945 25.400 227.645 311.095 ;
   LAYER M4 ;
    RECT 222.745 25.290 223.445 311.095 ;
   LAYER M4 ;
    RECT 220.645 25.290 221.345 311.095 ;
   LAYER M4 ;
    RECT 218.545 25.290 219.245 311.095 ;
   LAYER M4 ;
    RECT 216.445 25.290 217.145 311.095 ;
   LAYER M4 ;
    RECT 214.345 25.290 215.045 311.095 ;
   LAYER M4 ;
    RECT 212.245 25.290 212.945 311.095 ;
   LAYER M4 ;
    RECT 210.145 25.400 210.845 311.095 ;
   LAYER M4 ;
    RECT 205.945 25.290 206.645 311.095 ;
   LAYER M4 ;
    RECT 203.845 25.290 204.545 311.095 ;
   LAYER M4 ;
    RECT 201.745 25.290 202.445 311.095 ;
   LAYER M4 ;
    RECT 199.645 25.290 200.345 311.095 ;
   LAYER M4 ;
    RECT 197.545 25.290 198.245 311.095 ;
   LAYER M4 ;
    RECT 195.445 25.290 196.145 311.095 ;
   LAYER M4 ;
    RECT 193.345 25.400 194.045 311.095 ;
   LAYER M4 ;
    RECT 189.145 25.290 189.845 311.095 ;
   LAYER M4 ;
    RECT 187.045 25.290 187.745 311.095 ;
   LAYER M4 ;
    RECT 184.945 25.290 185.645 311.095 ;
   LAYER M4 ;
    RECT 182.845 25.290 183.545 311.095 ;
   LAYER M4 ;
    RECT 180.745 25.290 181.445 311.095 ;
   LAYER M4 ;
    RECT 178.645 25.290 179.345 311.095 ;
   LAYER M4 ;
    RECT 176.545 25.400 177.245 311.095 ;
   LAYER M4 ;
    RECT 172.345 25.290 173.045 311.095 ;
   LAYER M4 ;
    RECT 170.245 25.290 170.945 311.095 ;
   LAYER M4 ;
    RECT 168.145 25.290 168.845 311.095 ;
   LAYER M4 ;
    RECT 166.045 25.360 166.745 311.095 ;
   LAYER M4 ;
    RECT 163.945 25.360 164.645 311.095 ;
   LAYER M4 ;
    RECT 162.735 25.360 163.115 311.095 ;
   LAYER M4 ;
    RECT 161.530 25.360 162.510 311.095 ;
   LAYER M4 ;
    RECT 160.100 25.360 160.500 311.095 ;
   LAYER M4 ;
    RECT 158.605 25.360 159.105 311.095 ;
   LAYER M4 ;
    RECT 155.745 25.360 156.805 311.095 ;
   LAYER M4 ;
    RECT 155.065 25.360 155.465 311.095 ;
   LAYER M4 ;
    RECT 153.050 25.360 154.110 311.095 ;
   LAYER M4 ;
    RECT 151.035 25.360 151.435 311.095 ;
   LAYER M4 ;
    RECT 148.370 25.360 149.325 311.095 ;
   LAYER M4 ;
    RECT 144.910 25.360 145.550 311.095 ;
   LAYER M4 ;
    RECT 143.310 25.360 143.900 311.095 ;
   LAYER M4 ;
    RECT 139.395 25.360 140.195 311.095 ;
   LAYER M4 ;
    RECT 137.130 25.360 137.770 311.095 ;
   LAYER M4 ;
    RECT 133.505 25.290 134.205 311.095 ;
   LAYER M4 ;
    RECT 131.405 25.290 132.105 311.095 ;
   LAYER M4 ;
    RECT 129.305 25.290 130.005 311.095 ;
   LAYER M4 ;
    RECT 127.205 25.400 127.905 311.095 ;
   LAYER M4 ;
    RECT 123.005 25.290 123.705 311.095 ;
   LAYER M4 ;
    RECT 120.905 25.290 121.605 311.095 ;
   LAYER M4 ;
    RECT 118.805 25.290 119.505 311.095 ;
   LAYER M4 ;
    RECT 116.705 25.290 117.405 311.095 ;
   LAYER M4 ;
    RECT 114.605 25.290 115.305 311.095 ;
   LAYER M4 ;
    RECT 112.505 25.290 113.205 311.095 ;
   LAYER M4 ;
    RECT 110.405 25.400 111.105 311.095 ;
   LAYER M4 ;
    RECT 106.205 25.290 106.905 311.095 ;
   LAYER M4 ;
    RECT 104.105 25.290 104.805 311.095 ;
   LAYER M4 ;
    RECT 102.005 25.290 102.705 311.095 ;
   LAYER M4 ;
    RECT 99.905 25.290 100.605 311.095 ;
   LAYER M4 ;
    RECT 97.805 25.290 98.505 311.095 ;
   LAYER M4 ;
    RECT 95.705 25.290 96.405 311.095 ;
   LAYER M4 ;
    RECT 93.605 25.400 94.305 311.095 ;
   LAYER M4 ;
    RECT 89.405 25.290 90.105 311.095 ;
   LAYER M4 ;
    RECT 87.305 25.290 88.005 311.095 ;
   LAYER M4 ;
    RECT 85.205 25.290 85.905 311.095 ;
   LAYER M4 ;
    RECT 83.105 25.290 83.805 311.095 ;
   LAYER M4 ;
    RECT 81.005 25.290 81.705 311.095 ;
   LAYER M4 ;
    RECT 78.905 25.290 79.605 311.095 ;
   LAYER M4 ;
    RECT 76.805 25.400 77.505 311.095 ;
   LAYER M4 ;
    RECT 72.605 25.290 73.305 311.095 ;
   LAYER M4 ;
    RECT 70.505 25.290 71.205 311.095 ;
   LAYER M4 ;
    RECT 68.405 25.290 69.105 311.095 ;
   LAYER M4 ;
    RECT 66.305 25.290 67.005 311.095 ;
   LAYER M4 ;
    RECT 64.205 25.290 64.905 311.095 ;
   LAYER M4 ;
    RECT 62.105 25.290 62.805 311.095 ;
   LAYER M4 ;
    RECT 60.005 25.400 60.705 311.095 ;
   LAYER M4 ;
    RECT 55.805 25.290 56.505 311.095 ;
   LAYER M4 ;
    RECT 53.705 25.290 54.405 311.095 ;
   LAYER M4 ;
    RECT 51.605 25.290 52.305 311.095 ;
   LAYER M4 ;
    RECT 49.505 25.290 50.205 311.095 ;
   LAYER M4 ;
    RECT 47.405 25.290 48.105 311.095 ;
   LAYER M4 ;
    RECT 45.305 25.290 46.005 311.095 ;
   LAYER M4 ;
    RECT 43.205 25.400 43.905 311.095 ;
   LAYER M4 ;
    RECT 39.005 25.290 39.705 311.095 ;
   LAYER M4 ;
    RECT 0.495 0.760 303.920 1.140 ;
   LAYER M4 ;
    RECT 0.495 3.075 303.920 3.455 ;
   LAYER M4 ;
    RECT 0.495 4.095 303.920 5.095 ;
   LAYER M4 ;
    RECT 0.495 6.605 303.920 6.985 ;
   LAYER M4 ;
    RECT 0.495 8.980 303.920 9.680 ;
   LAYER M4 ;
    RECT 0.495 11.780 303.920 11.960 ;
  END
 END vdd
 OBS
  LAYER M1 ;
   RECT 0.050 0.050 304.750 311.750 ;
  LAYER M2 ;
   RECT 0.050 0.050 304.750 311.750 ;
  LAYER VIA2 ;
   RECT 5.850 0.050 5.950 0.570 ;
  LAYER VIA2 ;
   RECT 7.250 0.050 7.350 0.570 ;
  LAYER VIA2 ;
   RECT 11.450 0.050 11.550 0.570 ;
  LAYER VIA2 ;
   RECT 12.850 0.050 12.950 0.570 ;
  LAYER VIA2 ;
   RECT 22.650 0.050 22.750 0.570 ;
  LAYER VIA2 ;
   RECT 24.050 0.050 24.150 0.570 ;
  LAYER VIA2 ;
   RECT 28.250 0.050 28.350 0.570 ;
  LAYER VIA2 ;
   RECT 29.650 0.050 29.750 0.570 ;
  LAYER VIA2 ;
   RECT 39.450 0.050 39.550 0.570 ;
  LAYER VIA2 ;
   RECT 40.850 0.050 40.950 0.570 ;
  LAYER VIA2 ;
   RECT 45.050 0.050 45.150 0.570 ;
  LAYER VIA2 ;
   RECT 46.450 0.050 46.550 0.570 ;
  LAYER VIA2 ;
   RECT 56.250 0.050 56.350 0.570 ;
  LAYER VIA2 ;
   RECT 57.650 0.050 57.750 0.570 ;
  LAYER VIA2 ;
   RECT 61.850 0.050 61.950 0.570 ;
  LAYER VIA2 ;
   RECT 63.250 0.050 63.350 0.570 ;
  LAYER VIA2 ;
   RECT 73.050 0.050 73.150 0.570 ;
  LAYER VIA2 ;
   RECT 74.450 0.050 74.550 0.570 ;
  LAYER VIA2 ;
   RECT 78.650 0.050 78.750 0.570 ;
  LAYER VIA2 ;
   RECT 80.050 0.050 80.150 0.570 ;
  LAYER VIA2 ;
   RECT 89.850 0.050 89.950 0.570 ;
  LAYER VIA2 ;
   RECT 91.250 0.050 91.350 0.570 ;
  LAYER VIA2 ;
   RECT 95.450 0.050 95.550 0.570 ;
  LAYER VIA2 ;
   RECT 96.850 0.050 96.950 0.570 ;
  LAYER VIA2 ;
   RECT 106.650 0.050 106.750 0.570 ;
  LAYER VIA2 ;
   RECT 108.050 0.050 108.150 0.570 ;
  LAYER VIA2 ;
   RECT 112.250 0.050 112.350 0.570 ;
  LAYER VIA2 ;
   RECT 113.650 0.050 113.750 0.570 ;
  LAYER VIA2 ;
   RECT 123.450 0.050 123.550 0.570 ;
  LAYER VIA2 ;
   RECT 124.850 0.050 124.950 0.570 ;
  LAYER VIA2 ;
   RECT 129.050 0.050 129.150 0.570 ;
  LAYER VIA2 ;
   RECT 130.450 0.050 130.550 0.570 ;
  LAYER VIA2 ;
   RECT 136.650 0.050 136.750 0.570 ;
  LAYER VIA2 ;
   RECT 137.450 0.050 137.550 0.570 ;
  LAYER VIA2 ;
   RECT 143.650 0.050 143.750 0.570 ;
  LAYER VIA2 ;
   RECT 146.050 0.050 146.150 0.570 ;
  LAYER VIA2 ;
   RECT 147.450 0.050 147.550 0.570 ;
  LAYER VIA2 ;
   RECT 148.250 0.050 148.350 0.570 ;
  LAYER VIA2 ;
   RECT 148.850 0.050 148.950 0.570 ;
  LAYER VIA2 ;
   RECT 149.450 0.050 149.550 0.570 ;
  LAYER VIA2 ;
   RECT 150.250 0.050 150.350 0.570 ;
  LAYER VIA2 ;
   RECT 151.850 0.050 151.950 0.570 ;
  LAYER VIA2 ;
   RECT 153.250 0.050 153.350 0.570 ;
  LAYER VIA2 ;
   RECT 155.850 0.050 155.950 0.570 ;
  LAYER VIA2 ;
   RECT 156.450 0.050 156.550 0.570 ;
  LAYER VIA2 ;
   RECT 160.650 0.050 160.750 0.570 ;
  LAYER VIA2 ;
   RECT 161.250 0.050 161.350 0.570 ;
  LAYER VIA2 ;
   RECT 162.050 0.050 162.150 0.570 ;
  LAYER VIA2 ;
   RECT 172.850 0.050 172.950 0.570 ;
  LAYER VIA2 ;
   RECT 174.250 0.050 174.350 0.570 ;
  LAYER VIA2 ;
   RECT 178.250 0.050 178.350 0.570 ;
  LAYER VIA2 ;
   RECT 179.650 0.050 179.750 0.570 ;
  LAYER VIA2 ;
   RECT 189.650 0.050 189.750 0.570 ;
  LAYER VIA2 ;
   RECT 191.050 0.050 191.150 0.570 ;
  LAYER VIA2 ;
   RECT 195.050 0.050 195.150 0.570 ;
  LAYER VIA2 ;
   RECT 196.450 0.050 196.550 0.570 ;
  LAYER VIA2 ;
   RECT 206.450 0.050 206.550 0.570 ;
  LAYER VIA2 ;
   RECT 207.850 0.050 207.950 0.570 ;
  LAYER VIA2 ;
   RECT 211.850 0.050 211.950 0.570 ;
  LAYER VIA2 ;
   RECT 213.250 0.050 213.350 0.570 ;
  LAYER VIA2 ;
   RECT 223.250 0.050 223.350 0.570 ;
  LAYER VIA2 ;
   RECT 224.650 0.050 224.750 0.570 ;
  LAYER VIA2 ;
   RECT 228.650 0.050 228.750 0.570 ;
  LAYER VIA2 ;
   RECT 230.050 0.050 230.150 0.570 ;
  LAYER VIA2 ;
   RECT 240.050 0.050 240.150 0.570 ;
  LAYER VIA2 ;
   RECT 241.450 0.050 241.550 0.570 ;
  LAYER VIA2 ;
   RECT 245.450 0.050 245.550 0.570 ;
  LAYER VIA2 ;
   RECT 246.850 0.050 246.950 0.570 ;
  LAYER VIA2 ;
   RECT 256.850 0.050 256.950 0.570 ;
  LAYER VIA2 ;
   RECT 258.250 0.050 258.350 0.570 ;
  LAYER VIA2 ;
   RECT 262.250 0.050 262.350 0.570 ;
  LAYER VIA2 ;
   RECT 263.650 0.050 263.750 0.570 ;
  LAYER VIA2 ;
   RECT 273.650 0.050 273.750 0.570 ;
  LAYER VIA2 ;
   RECT 275.050 0.050 275.150 0.570 ;
  LAYER VIA2 ;
   RECT 279.050 0.050 279.150 0.570 ;
  LAYER VIA2 ;
   RECT 280.450 0.050 280.550 0.570 ;
  LAYER VIA2 ;
   RECT 290.450 0.050 290.550 0.570 ;
  LAYER VIA2 ;
   RECT 291.850 0.050 291.950 0.570 ;
  LAYER VIA2 ;
   RECT 295.850 0.050 295.950 0.570 ;
  LAYER VIA2 ;
   RECT 297.250 0.050 297.350 0.570 ;
  LAYER VIA2 ;
   RECT 303.050 0.050 303.150 0.570 ;
  LAYER M3 ;
   RECT 0.050 0.050 304.750 311.750 ;
  LAYER M4 ;
   RECT 0.050 0.050 304.750 311.750 ;
 END
END ST_SPHDL_4096x32m8_L

END LIBRARY
