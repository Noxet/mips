
module regfile ( clk, rst_n, .regfile_i({\regfile_i[ADRREAD0][4] , 
        \regfile_i[ADRREAD0][3] , \regfile_i[ADRREAD0][2] , 
        \regfile_i[ADRREAD0][1] , \regfile_i[ADRREAD0][0] , 
        \regfile_i[ADRREAD1][4] , \regfile_i[ADRREAD1][3] , 
        \regfile_i[ADRREAD1][2] , \regfile_i[ADRREAD1][1] , 
        \regfile_i[ADRREAD1][0] , \regfile_i[ADRWRITE][4] , 
        \regfile_i[ADRWRITE][3] , \regfile_i[ADRWRITE][2] , 
        \regfile_i[ADRWRITE][1] , \regfile_i[ADRWRITE][0] , 
        \regfile_i[WRITE_DATA][31] , \regfile_i[WRITE_DATA][30] , 
        \regfile_i[WRITE_DATA][29] , \regfile_i[WRITE_DATA][28] , 
        \regfile_i[WRITE_DATA][27] , \regfile_i[WRITE_DATA][26] , 
        \regfile_i[WRITE_DATA][25] , \regfile_i[WRITE_DATA][24] , 
        \regfile_i[WRITE_DATA][23] , \regfile_i[WRITE_DATA][22] , 
        \regfile_i[WRITE_DATA][21] , \regfile_i[WRITE_DATA][20] , 
        \regfile_i[WRITE_DATA][19] , \regfile_i[WRITE_DATA][18] , 
        \regfile_i[WRITE_DATA][17] , \regfile_i[WRITE_DATA][16] , 
        \regfile_i[WRITE_DATA][15] , \regfile_i[WRITE_DATA][14] , 
        \regfile_i[WRITE_DATA][13] , \regfile_i[WRITE_DATA][12] , 
        \regfile_i[WRITE_DATA][11] , \regfile_i[WRITE_DATA][10] , 
        \regfile_i[WRITE_DATA][9] , \regfile_i[WRITE_DATA][8] , 
        \regfile_i[WRITE_DATA][7] , \regfile_i[WRITE_DATA][6] , 
        \regfile_i[WRITE_DATA][5] , \regfile_i[WRITE_DATA][4] , 
        \regfile_i[WRITE_DATA][3] , \regfile_i[WRITE_DATA][2] , 
        \regfile_i[WRITE_DATA][1] , \regfile_i[WRITE_DATA][0] , 
        \regfile_i[FORWARD_A] , \regfile_i[FORWARD_B] , \regfile_i[WR_EN] }), 
    .regfile_o({\regfile_o[READ_DATA0][31] , \regfile_o[READ_DATA0][30] , 
        \regfile_o[READ_DATA0][29] , \regfile_o[READ_DATA0][28] , 
        \regfile_o[READ_DATA0][27] , \regfile_o[READ_DATA0][26] , 
        \regfile_o[READ_DATA0][25] , \regfile_o[READ_DATA0][24] , 
        \regfile_o[READ_DATA0][23] , \regfile_o[READ_DATA0][22] , 
        \regfile_o[READ_DATA0][21] , \regfile_o[READ_DATA0][20] , 
        \regfile_o[READ_DATA0][19] , \regfile_o[READ_DATA0][18] , 
        \regfile_o[READ_DATA0][17] , \regfile_o[READ_DATA0][16] , 
        \regfile_o[READ_DATA0][15] , \regfile_o[READ_DATA0][14] , 
        \regfile_o[READ_DATA0][13] , \regfile_o[READ_DATA0][12] , 
        \regfile_o[READ_DATA0][11] , \regfile_o[READ_DATA0][10] , 
        \regfile_o[READ_DATA0][9] , \regfile_o[READ_DATA0][8] , 
        \regfile_o[READ_DATA0][7] , \regfile_o[READ_DATA0][6] , 
        \regfile_o[READ_DATA0][5] , \regfile_o[READ_DATA0][4] , 
        \regfile_o[READ_DATA0][3] , \regfile_o[READ_DATA0][2] , 
        \regfile_o[READ_DATA0][1] , \regfile_o[READ_DATA0][0] , 
        \regfile_o[READ_DATA1][31] , \regfile_o[READ_DATA1][30] , 
        \regfile_o[READ_DATA1][29] , \regfile_o[READ_DATA1][28] , 
        \regfile_o[READ_DATA1][27] , \regfile_o[READ_DATA1][26] , 
        \regfile_o[READ_DATA1][25] , \regfile_o[READ_DATA1][24] , 
        \regfile_o[READ_DATA1][23] , \regfile_o[READ_DATA1][22] , 
        \regfile_o[READ_DATA1][21] , \regfile_o[READ_DATA1][20] , 
        \regfile_o[READ_DATA1][19] , \regfile_o[READ_DATA1][18] , 
        \regfile_o[READ_DATA1][17] , \regfile_o[READ_DATA1][16] , 
        \regfile_o[READ_DATA1][15] , \regfile_o[READ_DATA1][14] , 
        \regfile_o[READ_DATA1][13] , \regfile_o[READ_DATA1][12] , 
        \regfile_o[READ_DATA1][11] , \regfile_o[READ_DATA1][10] , 
        \regfile_o[READ_DATA1][9] , \regfile_o[READ_DATA1][8] , 
        \regfile_o[READ_DATA1][7] , \regfile_o[READ_DATA1][6] , 
        \regfile_o[READ_DATA1][5] , \regfile_o[READ_DATA1][4] , 
        \regfile_o[READ_DATA1][3] , \regfile_o[READ_DATA1][2] , 
        \regfile_o[READ_DATA1][1] , \regfile_o[READ_DATA1][0] }) );
  input clk, rst_n, \regfile_i[ADRREAD0][4] , \regfile_i[ADRREAD0][3] ,
         \regfile_i[ADRREAD0][2] , \regfile_i[ADRREAD0][1] ,
         \regfile_i[ADRREAD0][0] , \regfile_i[ADRREAD1][4] ,
         \regfile_i[ADRREAD1][3] , \regfile_i[ADRREAD1][2] ,
         \regfile_i[ADRREAD1][1] , \regfile_i[ADRREAD1][0] ,
         \regfile_i[ADRWRITE][4] , \regfile_i[ADRWRITE][3] ,
         \regfile_i[ADRWRITE][2] , \regfile_i[ADRWRITE][1] ,
         \regfile_i[ADRWRITE][0] , \regfile_i[WRITE_DATA][31] ,
         \regfile_i[WRITE_DATA][30] , \regfile_i[WRITE_DATA][29] ,
         \regfile_i[WRITE_DATA][28] , \regfile_i[WRITE_DATA][27] ,
         \regfile_i[WRITE_DATA][26] , \regfile_i[WRITE_DATA][25] ,
         \regfile_i[WRITE_DATA][24] , \regfile_i[WRITE_DATA][23] ,
         \regfile_i[WRITE_DATA][22] , \regfile_i[WRITE_DATA][21] ,
         \regfile_i[WRITE_DATA][20] , \regfile_i[WRITE_DATA][19] ,
         \regfile_i[WRITE_DATA][18] , \regfile_i[WRITE_DATA][17] ,
         \regfile_i[WRITE_DATA][16] , \regfile_i[WRITE_DATA][15] ,
         \regfile_i[WRITE_DATA][14] , \regfile_i[WRITE_DATA][13] ,
         \regfile_i[WRITE_DATA][12] , \regfile_i[WRITE_DATA][11] ,
         \regfile_i[WRITE_DATA][10] , \regfile_i[WRITE_DATA][9] ,
         \regfile_i[WRITE_DATA][8] , \regfile_i[WRITE_DATA][7] ,
         \regfile_i[WRITE_DATA][6] , \regfile_i[WRITE_DATA][5] ,
         \regfile_i[WRITE_DATA][4] , \regfile_i[WRITE_DATA][3] ,
         \regfile_i[WRITE_DATA][2] , \regfile_i[WRITE_DATA][1] ,
         \regfile_i[WRITE_DATA][0] , \regfile_i[FORWARD_A] ,
         \regfile_i[FORWARD_B] , \regfile_i[WR_EN] ;
  output \regfile_o[READ_DATA0][31] , \regfile_o[READ_DATA0][30] ,
         \regfile_o[READ_DATA0][29] , \regfile_o[READ_DATA0][28] ,
         \regfile_o[READ_DATA0][27] , \regfile_o[READ_DATA0][26] ,
         \regfile_o[READ_DATA0][25] , \regfile_o[READ_DATA0][24] ,
         \regfile_o[READ_DATA0][23] , \regfile_o[READ_DATA0][22] ,
         \regfile_o[READ_DATA0][21] , \regfile_o[READ_DATA0][20] ,
         \regfile_o[READ_DATA0][19] , \regfile_o[READ_DATA0][18] ,
         \regfile_o[READ_DATA0][17] , \regfile_o[READ_DATA0][16] ,
         \regfile_o[READ_DATA0][15] , \regfile_o[READ_DATA0][14] ,
         \regfile_o[READ_DATA0][13] , \regfile_o[READ_DATA0][12] ,
         \regfile_o[READ_DATA0][11] , \regfile_o[READ_DATA0][10] ,
         \regfile_o[READ_DATA0][9] , \regfile_o[READ_DATA0][8] ,
         \regfile_o[READ_DATA0][7] , \regfile_o[READ_DATA0][6] ,
         \regfile_o[READ_DATA0][5] , \regfile_o[READ_DATA0][4] ,
         \regfile_o[READ_DATA0][3] , \regfile_o[READ_DATA0][2] ,
         \regfile_o[READ_DATA0][1] , \regfile_o[READ_DATA0][0] ,
         \regfile_o[READ_DATA1][31] , \regfile_o[READ_DATA1][30] ,
         \regfile_o[READ_DATA1][29] , \regfile_o[READ_DATA1][28] ,
         \regfile_o[READ_DATA1][27] , \regfile_o[READ_DATA1][26] ,
         \regfile_o[READ_DATA1][25] , \regfile_o[READ_DATA1][24] ,
         \regfile_o[READ_DATA1][23] , \regfile_o[READ_DATA1][22] ,
         \regfile_o[READ_DATA1][21] , \regfile_o[READ_DATA1][20] ,
         \regfile_o[READ_DATA1][19] , \regfile_o[READ_DATA1][18] ,
         \regfile_o[READ_DATA1][17] , \regfile_o[READ_DATA1][16] ,
         \regfile_o[READ_DATA1][15] , \regfile_o[READ_DATA1][14] ,
         \regfile_o[READ_DATA1][13] , \regfile_o[READ_DATA1][12] ,
         \regfile_o[READ_DATA1][11] , \regfile_o[READ_DATA1][10] ,
         \regfile_o[READ_DATA1][9] , \regfile_o[READ_DATA1][8] ,
         \regfile_o[READ_DATA1][7] , \regfile_o[READ_DATA1][6] ,
         \regfile_o[READ_DATA1][5] , \regfile_o[READ_DATA1][4] ,
         \regfile_o[READ_DATA1][3] , \regfile_o[READ_DATA1][2] ,
         \regfile_o[READ_DATA1][1] , \regfile_o[READ_DATA1][0] ;
  wire   \registers[31][31] , \registers[31][30] , \registers[31][29] ,
         \registers[31][28] , \registers[31][27] , \registers[31][26] ,
         \registers[31][25] , \registers[31][24] , \registers[31][23] ,
         \registers[31][22] , \registers[31][21] , \registers[31][20] ,
         \registers[31][19] , \registers[31][18] , \registers[31][17] ,
         \registers[31][16] , \registers[31][15] , \registers[31][14] ,
         \registers[31][13] , \registers[31][12] , \registers[31][11] ,
         \registers[31][10] , \registers[31][9] , \registers[31][8] ,
         \registers[31][7] , \registers[31][6] , \registers[31][5] ,
         \registers[31][4] , \registers[31][3] , \registers[31][2] ,
         \registers[31][1] , \registers[31][0] , \registers[30][31] ,
         \registers[30][30] , \registers[30][29] , \registers[30][28] ,
         \registers[30][27] , \registers[30][26] , \registers[30][25] ,
         \registers[30][24] , \registers[30][23] , \registers[30][22] ,
         \registers[30][21] , \registers[30][20] , \registers[30][19] ,
         \registers[30][18] , \registers[30][17] , \registers[30][16] ,
         \registers[30][15] , \registers[30][14] , \registers[30][13] ,
         \registers[30][12] , \registers[30][11] , \registers[30][10] ,
         \registers[30][9] , \registers[30][8] , \registers[30][7] ,
         \registers[30][6] , \registers[30][5] , \registers[30][4] ,
         \registers[30][3] , \registers[30][2] , \registers[30][1] ,
         \registers[30][0] , \registers[25][31] , \registers[25][30] ,
         \registers[25][29] , \registers[25][28] , \registers[25][27] ,
         \registers[25][26] , \registers[25][25] , \registers[25][24] ,
         \registers[25][23] , \registers[25][22] , \registers[25][21] ,
         \registers[25][20] , \registers[25][19] , \registers[25][18] ,
         \registers[25][17] , \registers[25][16] , \registers[25][15] ,
         \registers[25][14] , \registers[25][13] , \registers[25][12] ,
         \registers[25][11] , \registers[25][10] , \registers[25][9] ,
         \registers[25][8] , \registers[25][7] , \registers[25][6] ,
         \registers[25][5] , \registers[25][4] , \registers[25][3] ,
         \registers[25][2] , \registers[25][1] , \registers[25][0] ,
         \registers[24][31] , \registers[24][30] , \registers[24][29] ,
         \registers[24][28] , \registers[24][27] , \registers[24][26] ,
         \registers[24][25] , \registers[24][24] , \registers[24][23] ,
         \registers[24][22] , \registers[24][21] , \registers[24][20] ,
         \registers[24][19] , \registers[24][18] , \registers[24][17] ,
         \registers[24][16] , \registers[24][15] , \registers[24][14] ,
         \registers[24][13] , \registers[24][12] , \registers[24][11] ,
         \registers[24][10] , \registers[24][9] , \registers[24][8] ,
         \registers[24][7] , \registers[24][6] , \registers[24][5] ,
         \registers[24][4] , \registers[24][3] , \registers[24][2] ,
         \registers[24][1] , \registers[24][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[22][31] , \registers[22][30] ,
         \registers[22][29] , \registers[22][28] , \registers[22][27] ,
         \registers[22][26] , \registers[22][25] , \registers[22][24] ,
         \registers[22][23] , \registers[22][22] , \registers[22][21] ,
         \registers[22][20] , \registers[22][19] , \registers[22][18] ,
         \registers[22][17] , \registers[22][16] , \registers[22][15] ,
         \registers[22][14] , \registers[22][13] , \registers[22][12] ,
         \registers[22][11] , \registers[22][10] , \registers[22][9] ,
         \registers[22][8] , \registers[22][7] , \registers[22][6] ,
         \registers[22][5] , \registers[22][4] , \registers[22][3] ,
         \registers[22][2] , \registers[22][1] , \registers[22][0] ,
         \registers[21][31] , \registers[21][30] , \registers[21][29] ,
         \registers[21][28] , \registers[21][27] , \registers[21][26] ,
         \registers[21][25] , \registers[21][24] , \registers[21][23] ,
         \registers[21][22] , \registers[21][21] , \registers[21][20] ,
         \registers[21][19] , \registers[21][18] , \registers[21][17] ,
         \registers[21][16] , \registers[21][15] , \registers[21][14] ,
         \registers[21][13] , \registers[21][12] , \registers[21][11] ,
         \registers[21][10] , \registers[21][9] , \registers[21][8] ,
         \registers[21][7] , \registers[21][6] , \registers[21][5] ,
         \registers[21][4] , \registers[21][3] , \registers[21][2] ,
         \registers[21][1] , \registers[21][0] , \registers[20][31] ,
         \registers[20][30] , \registers[20][29] , \registers[20][28] ,
         \registers[20][27] , \registers[20][26] , \registers[20][25] ,
         \registers[20][24] , \registers[20][23] , \registers[20][22] ,
         \registers[20][21] , \registers[20][20] , \registers[20][19] ,
         \registers[20][18] , \registers[20][17] , \registers[20][16] ,
         \registers[20][15] , \registers[20][14] , \registers[20][13] ,
         \registers[20][12] , \registers[20][11] , \registers[20][10] ,
         \registers[20][9] , \registers[20][8] , \registers[20][7] ,
         \registers[20][6] , \registers[20][5] , \registers[20][4] ,
         \registers[20][3] , \registers[20][2] , \registers[20][1] ,
         \registers[20][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[18][31] , \registers[18][30] , \registers[18][29] ,
         \registers[18][28] , \registers[18][27] , \registers[18][26] ,
         \registers[18][25] , \registers[18][24] , \registers[18][23] ,
         \registers[18][22] , \registers[18][21] , \registers[18][20] ,
         \registers[18][19] , \registers[18][18] , \registers[18][17] ,
         \registers[18][16] , \registers[18][15] , \registers[18][14] ,
         \registers[18][13] , \registers[18][12] , \registers[18][11] ,
         \registers[18][10] , \registers[18][9] , \registers[18][8] ,
         \registers[18][7] , \registers[18][6] , \registers[18][5] ,
         \registers[18][4] , \registers[18][3] , \registers[18][2] ,
         \registers[18][1] , \registers[18][0] , \registers[17][31] ,
         \registers[17][30] , \registers[17][29] , \registers[17][28] ,
         \registers[17][27] , \registers[17][26] , \registers[17][25] ,
         \registers[17][24] , \registers[17][23] , \registers[17][22] ,
         \registers[17][21] , \registers[17][20] , \registers[17][19] ,
         \registers[17][18] , \registers[17][17] , \registers[17][16] ,
         \registers[17][15] , \registers[17][14] , \registers[17][13] ,
         \registers[17][12] , \registers[17][11] , \registers[17][10] ,
         \registers[17][9] , \registers[17][8] , \registers[17][7] ,
         \registers[17][6] , \registers[17][5] , \registers[17][4] ,
         \registers[17][3] , \registers[17][2] , \registers[17][1] ,
         \registers[17][0] , \registers[16][31] , \registers[16][30] ,
         \registers[16][29] , \registers[16][28] , \registers[16][27] ,
         \registers[16][26] , \registers[16][25] , \registers[16][24] ,
         \registers[16][23] , \registers[16][22] , \registers[16][21] ,
         \registers[16][20] , \registers[16][19] , \registers[16][18] ,
         \registers[16][17] , \registers[16][16] , \registers[16][15] ,
         \registers[16][14] , \registers[16][13] , \registers[16][12] ,
         \registers[16][11] , \registers[16][10] , \registers[16][9] ,
         \registers[16][8] , \registers[16][7] , \registers[16][6] ,
         \registers[16][5] , \registers[16][4] , \registers[16][3] ,
         \registers[16][2] , \registers[16][1] , \registers[16][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[12][31] ,
         \registers[12][30] , \registers[12][29] , \registers[12][28] ,
         \registers[12][27] , \registers[12][26] , \registers[12][25] ,
         \registers[12][24] , \registers[12][23] , \registers[12][22] ,
         \registers[12][21] , \registers[12][20] , \registers[12][19] ,
         \registers[12][18] , \registers[12][17] , \registers[12][16] ,
         \registers[12][15] , \registers[12][14] , \registers[12][13] ,
         \registers[12][12] , \registers[12][11] , \registers[12][10] ,
         \registers[12][9] , \registers[12][8] , \registers[12][7] ,
         \registers[12][6] , \registers[12][5] , \registers[12][4] ,
         \registers[12][3] , \registers[12][2] , \registers[12][1] ,
         \registers[12][0] , \registers[11][31] , \registers[11][30] ,
         \registers[11][29] , \registers[11][28] , \registers[11][27] ,
         \registers[11][26] , \registers[11][25] , \registers[11][24] ,
         \registers[11][23] , \registers[11][22] , \registers[11][21] ,
         \registers[11][20] , \registers[11][19] , \registers[11][18] ,
         \registers[11][17] , \registers[11][16] , \registers[11][15] ,
         \registers[11][14] , \registers[11][13] , \registers[11][12] ,
         \registers[11][11] , \registers[11][10] , \registers[11][9] ,
         \registers[11][8] , \registers[11][7] , \registers[11][6] ,
         \registers[11][5] , \registers[11][4] , \registers[11][3] ,
         \registers[11][2] , \registers[11][1] , \registers[11][0] ,
         \registers[10][31] , \registers[10][30] , \registers[10][29] ,
         \registers[10][28] , \registers[10][27] , \registers[10][26] ,
         \registers[10][25] , \registers[10][24] , \registers[10][23] ,
         \registers[10][22] , \registers[10][21] , \registers[10][20] ,
         \registers[10][19] , \registers[10][18] , \registers[10][17] ,
         \registers[10][16] , \registers[10][15] , \registers[10][14] ,
         \registers[10][13] , \registers[10][12] , \registers[10][11] ,
         \registers[10][10] , \registers[10][9] , \registers[10][8] ,
         \registers[10][7] , \registers[10][6] , \registers[10][5] ,
         \registers[10][4] , \registers[10][3] , \registers[10][2] ,
         \registers[10][1] , \registers[10][0] , \registers[7][31] ,
         \registers[7][30] , \registers[7][29] , \registers[7][28] ,
         \registers[7][27] , \registers[7][26] , \registers[7][25] ,
         \registers[7][24] , \registers[7][23] , \registers[7][22] ,
         \registers[7][21] , \registers[7][20] , \registers[7][19] ,
         \registers[7][18] , \registers[7][17] , \registers[7][16] ,
         \registers[7][15] , \registers[7][14] , \registers[7][13] ,
         \registers[7][12] , \registers[7][11] , \registers[7][10] ,
         \registers[7][9] , \registers[7][8] , \registers[7][7] ,
         \registers[7][6] , \registers[7][5] , \registers[7][4] ,
         \registers[7][3] , \registers[7][2] , \registers[7][1] ,
         \registers[7][0] , \registers[6][31] , \registers[6][30] ,
         \registers[6][29] , \registers[6][28] , \registers[6][27] ,
         \registers[6][26] , \registers[6][25] , \registers[6][24] ,
         \registers[6][23] , \registers[6][22] , \registers[6][21] ,
         \registers[6][20] , \registers[6][19] , \registers[6][18] ,
         \registers[6][17] , \registers[6][16] , \registers[6][15] ,
         \registers[6][14] , \registers[6][13] , \registers[6][12] ,
         \registers[6][11] , \registers[6][10] , \registers[6][9] ,
         \registers[6][8] , \registers[6][7] , \registers[6][6] ,
         \registers[6][5] , \registers[6][4] , \registers[6][3] ,
         \registers[6][2] , \registers[6][1] , \registers[6][0] ,
         \registers[5][31] , \registers[5][30] , \registers[5][29] ,
         \registers[5][28] , \registers[5][27] , \registers[5][26] ,
         \registers[5][25] , \registers[5][24] , \registers[5][23] ,
         \registers[5][22] , \registers[5][21] , \registers[5][20] ,
         \registers[5][19] , \registers[5][18] , \registers[5][17] ,
         \registers[5][16] , \registers[5][15] , \registers[5][14] ,
         \registers[5][13] , \registers[5][12] , \registers[5][11] ,
         \registers[5][10] , \registers[5][9] , \registers[5][8] ,
         \registers[5][7] , \registers[5][6] , \registers[5][5] ,
         \registers[5][4] , \registers[5][3] , \registers[5][2] ,
         \registers[5][1] , \registers[5][0] , \registers[4][31] ,
         \registers[4][30] , \registers[4][29] , \registers[4][28] ,
         \registers[4][27] , \registers[4][26] , \registers[4][25] ,
         \registers[4][24] , \registers[4][23] , \registers[4][22] ,
         \registers[4][21] , \registers[4][20] , \registers[4][19] ,
         \registers[4][18] , \registers[4][17] , \registers[4][16] ,
         \registers[4][15] , \registers[4][14] , \registers[4][13] ,
         \registers[4][12] , \registers[4][11] , \registers[4][10] ,
         \registers[4][9] , \registers[4][8] , \registers[4][7] ,
         \registers[4][6] , \registers[4][5] , \registers[4][4] ,
         \registers[4][3] , \registers[4][2] , \registers[4][1] ,
         \registers[4][0] , \registers[3][31] , \registers[3][30] ,
         \registers[3][29] , \registers[3][28] , \registers[3][27] ,
         \registers[3][26] , \registers[3][25] , \registers[3][24] ,
         \registers[3][23] , \registers[3][22] , \registers[3][21] ,
         \registers[3][20] , \registers[3][19] , \registers[3][18] ,
         \registers[3][17] , \registers[3][16] , \registers[3][15] ,
         \registers[3][14] , \registers[3][13] , \registers[3][12] ,
         \registers[3][11] , \registers[3][10] , \registers[3][9] ,
         \registers[3][8] , \registers[3][7] , \registers[3][6] ,
         \registers[3][5] , \registers[3][4] , \registers[3][3] ,
         \registers[3][2] , \registers[3][1] , \registers[3][0] ,
         \registers[2][31] , \registers[2][30] , \registers[2][29] ,
         \registers[2][28] , \registers[2][27] , \registers[2][26] ,
         \registers[2][25] , \registers[2][24] , \registers[2][23] ,
         \registers[2][22] , \registers[2][21] , \registers[2][20] ,
         \registers[2][19] , \registers[2][18] , \registers[2][17] ,
         \registers[2][16] , \registers[2][15] , \registers[2][14] ,
         \registers[2][13] , \registers[2][12] , \registers[2][11] ,
         \registers[2][10] , \registers[2][9] , \registers[2][8] ,
         \registers[2][7] , \registers[2][6] , \registers[2][5] ,
         \registers[2][4] , \registers[2][3] , \registers[2][2] ,
         \registers[2][1] , \registers[2][0] , \registers[1][31] ,
         \registers[1][30] , \registers[1][29] , \registers[1][28] ,
         \registers[1][27] , \registers[1][26] , \registers[1][25] ,
         \registers[1][24] , \registers[1][23] , \registers[1][22] ,
         \registers[1][21] , \registers[1][20] , \registers[1][19] ,
         \registers[1][18] , \registers[1][17] , \registers[1][16] ,
         \registers[1][15] , \registers[1][14] , \registers[1][13] ,
         \registers[1][12] , \registers[1][11] , \registers[1][10] ,
         \registers[1][9] , \registers[1][8] , \registers[1][7] ,
         \registers[1][6] , \registers[1][5] , \registers[1][4] ,
         \registers[1][3] , \registers[1][2] , \registers[1][1] ,
         \registers[1][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n795, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2824, n2825, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2841, n2846, n2847, n2848, n2849, n2850, n2851, n2853, n2855,
         n2856, n2857, n2859, n2860, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664;

  HS65_LH_DFPRQX9 \registers_reg[31][31]  ( .D(n2425), .CP(clk), .RN(n6539), 
        .Q(\registers[31][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][30]  ( .D(n2424), .CP(clk), .RN(n6569), 
        .Q(\registers[31][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][29]  ( .D(n2423), .CP(clk), .RN(n6571), 
        .Q(\registers[31][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][28]  ( .D(n2422), .CP(clk), .RN(n6570), 
        .Q(\registers[31][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][27]  ( .D(n2421), .CP(clk), .RN(n6570), 
        .Q(\registers[31][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][26]  ( .D(n2420), .CP(clk), .RN(n6569), 
        .Q(\registers[31][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][25]  ( .D(n2419), .CP(clk), .RN(n6572), 
        .Q(\registers[31][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][24]  ( .D(n2418), .CP(clk), .RN(n6572), 
        .Q(\registers[31][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][23]  ( .D(n2417), .CP(clk), .RN(n6572), 
        .Q(\registers[31][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][22]  ( .D(n2416), .CP(clk), .RN(n6572), 
        .Q(\registers[31][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][21]  ( .D(n2415), .CP(clk), .RN(n6568), 
        .Q(\registers[31][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][20]  ( .D(n2414), .CP(clk), .RN(n6568), 
        .Q(\registers[31][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][19]  ( .D(n2413), .CP(clk), .RN(n6568), 
        .Q(\registers[31][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][18]  ( .D(n2412), .CP(clk), .RN(n6568), 
        .Q(\registers[31][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][17]  ( .D(n2411), .CP(clk), .RN(n6568), 
        .Q(\registers[31][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][16]  ( .D(n2410), .CP(clk), .RN(n6568), 
        .Q(\registers[31][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][15]  ( .D(n2409), .CP(clk), .RN(n6568), 
        .Q(\registers[31][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][14]  ( .D(n2408), .CP(clk), .RN(n6568), 
        .Q(\registers[31][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][13]  ( .D(n2407), .CP(clk), .RN(n6578), 
        .Q(\registers[31][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][12]  ( .D(n2406), .CP(clk), .RN(n6578), 
        .Q(\registers[31][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][11]  ( .D(n2405), .CP(clk), .RN(n6578), 
        .Q(\registers[31][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][10]  ( .D(n2404), .CP(clk), .RN(n6578), 
        .Q(\registers[31][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][9]  ( .D(n2403), .CP(clk), .RN(n6580), 
        .Q(\registers[31][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][8]  ( .D(n2402), .CP(clk), .RN(n6580), 
        .Q(\registers[31][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][7]  ( .D(n2401), .CP(clk), .RN(n6580), 
        .Q(\registers[31][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][6]  ( .D(n2400), .CP(clk), .RN(n6580), 
        .Q(\registers[31][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][5]  ( .D(n2399), .CP(clk), .RN(n6580), 
        .Q(\registers[31][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][4]  ( .D(n2398), .CP(clk), .RN(n6580), 
        .Q(\registers[31][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][3]  ( .D(n2397), .CP(clk), .RN(n6580), 
        .Q(\registers[31][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][2]  ( .D(n2396), .CP(clk), .RN(n6580), 
        .Q(\registers[31][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][1]  ( .D(n2395), .CP(clk), .RN(n6578), 
        .Q(\registers[31][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][0]  ( .D(n2394), .CP(clk), .RN(n6578), 
        .Q(\registers[31][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][31]  ( .D(n2393), .CP(clk), .RN(n6583), 
        .Q(\registers[30][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][30]  ( .D(n2392), .CP(clk), .RN(n6583), 
        .Q(\registers[30][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][29]  ( .D(n2391), .CP(clk), .RN(n6583), 
        .Q(\registers[30][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][28]  ( .D(n2390), .CP(clk), .RN(n6583), 
        .Q(\registers[30][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][27]  ( .D(n2389), .CP(clk), .RN(n6584), 
        .Q(\registers[30][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][26]  ( .D(n2388), .CP(clk), .RN(n6584), 
        .Q(\registers[30][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][25]  ( .D(n2387), .CP(clk), .RN(n6584), 
        .Q(\registers[30][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][24]  ( .D(n2386), .CP(clk), .RN(n6584), 
        .Q(\registers[30][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][23]  ( .D(n2385), .CP(clk), .RN(n6579), 
        .Q(\registers[30][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][22]  ( .D(n2384), .CP(clk), .RN(n6579), 
        .Q(\registers[30][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][21]  ( .D(n2383), .CP(clk), .RN(n6585), 
        .Q(\registers[30][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][20]  ( .D(n2382), .CP(clk), .RN(n6583), 
        .Q(\registers[30][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][19]  ( .D(n2381), .CP(clk), .RN(n6583), 
        .Q(\registers[30][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][18]  ( .D(n2380), .CP(clk), .RN(n6583), 
        .Q(\registers[30][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][17]  ( .D(n2379), .CP(clk), .RN(n6582), 
        .Q(\registers[30][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][16]  ( .D(n2378), .CP(clk), .RN(n6582), 
        .Q(\registers[30][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][15]  ( .D(n2377), .CP(clk), .RN(n6582), 
        .Q(\registers[30][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][14]  ( .D(n2376), .CP(clk), .RN(n6582), 
        .Q(\registers[30][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][13]  ( .D(n2375), .CP(clk), .RN(n6582), 
        .Q(\registers[30][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][12]  ( .D(n2374), .CP(clk), .RN(n6582), 
        .Q(\registers[30][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][11]  ( .D(n2373), .CP(clk), .RN(n6582), 
        .Q(\registers[30][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][10]  ( .D(n2372), .CP(clk), .RN(n6582), 
        .Q(\registers[30][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][9]  ( .D(n2371), .CP(clk), .RN(n6583), 
        .Q(\registers[30][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][8]  ( .D(n2370), .CP(clk), .RN(n6583), 
        .Q(\registers[30][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][7]  ( .D(n2369), .CP(clk), .RN(n6585), 
        .Q(\registers[30][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][6]  ( .D(n2368), .CP(clk), .RN(n6585), 
        .Q(\registers[30][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][5]  ( .D(n2367), .CP(clk), .RN(n6585), 
        .Q(\registers[30][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][4]  ( .D(n2366), .CP(clk), .RN(n6585), 
        .Q(\registers[30][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][3]  ( .D(n2365), .CP(clk), .RN(n6585), 
        .Q(\registers[30][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][2]  ( .D(n2364), .CP(clk), .RN(n6585), 
        .Q(\registers[30][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][1]  ( .D(n2363), .CP(clk), .RN(n6585), 
        .Q(\registers[30][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][0]  ( .D(n2362), .CP(clk), .RN(n6585), 
        .Q(\registers[30][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][31]  ( .D(n2233), .CP(clk), .RN(n6586), 
        .Q(\registers[25][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][30]  ( .D(n2232), .CP(clk), .RN(n6586), 
        .Q(\registers[25][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][29]  ( .D(n2231), .CP(clk), .RN(n6589), 
        .Q(\registers[25][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][28]  ( .D(n2230), .CP(clk), .RN(n6589), 
        .Q(\registers[25][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][27]  ( .D(n2229), .CP(clk), .RN(n6589), 
        .Q(\registers[25][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][26]  ( .D(n2228), .CP(clk), .RN(n6589), 
        .Q(\registers[25][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][25]  ( .D(n2227), .CP(clk), .RN(n6586), 
        .Q(\registers[25][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][24]  ( .D(n2226), .CP(clk), .RN(n6586), 
        .Q(\registers[25][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][23]  ( .D(n2225), .CP(clk), .RN(n6585), 
        .Q(\registers[25][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][22]  ( .D(n2224), .CP(clk), .RN(n6585), 
        .Q(\registers[25][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][21]  ( .D(n2223), .CP(clk), .RN(n6585), 
        .Q(\registers[25][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][20]  ( .D(n2222), .CP(clk), .RN(n6583), 
        .Q(\registers[25][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][19]  ( .D(n2221), .CP(clk), .RN(n6583), 
        .Q(\registers[25][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][18]  ( .D(n2220), .CP(clk), .RN(n6583), 
        .Q(\registers[25][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][17]  ( .D(n2219), .CP(clk), .RN(n6588), 
        .Q(\registers[25][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][16]  ( .D(n2218), .CP(clk), .RN(n6588), 
        .Q(\registers[25][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][15]  ( .D(n2217), .CP(clk), .RN(n6588), 
        .Q(\registers[25][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][14]  ( .D(n2216), .CP(clk), .RN(n6586), 
        .Q(\registers[25][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][13]  ( .D(n2215), .CP(clk), .RN(n6584), 
        .Q(\registers[25][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][12]  ( .D(n2214), .CP(clk), .RN(n6584), 
        .Q(\registers[25][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][11]  ( .D(n2213), .CP(clk), .RN(n6584), 
        .Q(\registers[25][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][10]  ( .D(n2212), .CP(clk), .RN(n6584), 
        .Q(\registers[25][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][9]  ( .D(n2211), .CP(clk), .RN(n6584), 
        .Q(\registers[25][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][8]  ( .D(n2210), .CP(clk), .RN(n6584), 
        .Q(\registers[25][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][7]  ( .D(n2209), .CP(clk), .RN(n6584), 
        .Q(\registers[25][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][6]  ( .D(n2208), .CP(clk), .RN(n6584), 
        .Q(\registers[25][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][5]  ( .D(n2207), .CP(clk), .RN(n6586), 
        .Q(\registers[25][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][4]  ( .D(n2206), .CP(clk), .RN(n6586), 
        .Q(\registers[25][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][3]  ( .D(n2205), .CP(clk), .RN(n6586), 
        .Q(\registers[25][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][2]  ( .D(n2204), .CP(clk), .RN(n6586), 
        .Q(\registers[25][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][1]  ( .D(n2203), .CP(clk), .RN(n6586), 
        .Q(\registers[25][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][0]  ( .D(n2202), .CP(clk), .RN(n6586), 
        .Q(\registers[25][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][31]  ( .D(n2201), .CP(clk), .RN(n6591), 
        .Q(\registers[24][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][30]  ( .D(n2200), .CP(clk), .RN(n6591), 
        .Q(\registers[24][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][29]  ( .D(n2199), .CP(clk), .RN(n6591), 
        .Q(\registers[24][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][28]  ( .D(n2198), .CP(clk), .RN(n6591), 
        .Q(\registers[24][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][27]  ( .D(n2197), .CP(clk), .RN(n6590), 
        .Q(\registers[24][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][26]  ( .D(n2196), .CP(clk), .RN(n6592), 
        .Q(\registers[24][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][25]  ( .D(n2195), .CP(clk), .RN(n6592), 
        .Q(\registers[24][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][24]  ( .D(n2194), .CP(clk), .RN(n6592), 
        .Q(\registers[24][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][23]  ( .D(n2193), .CP(clk), .RN(n6590), 
        .Q(\registers[24][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][22]  ( .D(n2192), .CP(clk), .RN(n6590), 
        .Q(\registers[24][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][21]  ( .D(n2191), .CP(clk), .RN(n6590), 
        .Q(\registers[24][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][20]  ( .D(n2190), .CP(clk), .RN(n6590), 
        .Q(\registers[24][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][19]  ( .D(n2189), .CP(clk), .RN(n6588), 
        .Q(\registers[24][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][18]  ( .D(n2188), .CP(clk), .RN(n6588), 
        .Q(\registers[24][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][17]  ( .D(n2187), .CP(clk), .RN(n6588), 
        .Q(\registers[24][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][16]  ( .D(n2186), .CP(clk), .RN(n6588), 
        .Q(\registers[24][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][15]  ( .D(n2185), .CP(clk), .RN(n6588), 
        .Q(\registers[24][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][14]  ( .D(n2184), .CP(clk), .RN(n6590), 
        .Q(\registers[24][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][13]  ( .D(n2183), .CP(clk), .RN(n6590), 
        .Q(\registers[24][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][12]  ( .D(n2182), .CP(clk), .RN(n6590), 
        .Q(\registers[24][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][11]  ( .D(n2181), .CP(clk), .RN(n6590), 
        .Q(\registers[24][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][10]  ( .D(n2180), .CP(clk), .RN(n6589), 
        .Q(\registers[24][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][9]  ( .D(n2179), .CP(clk), .RN(n6589), 
        .Q(\registers[24][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][8]  ( .D(n2178), .CP(clk), .RN(n6589), 
        .Q(\registers[24][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][7]  ( .D(n2177), .CP(clk), .RN(n6589), 
        .Q(\registers[24][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][6]  ( .D(n2176), .CP(clk), .RN(n6589), 
        .Q(\registers[24][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][5]  ( .D(n2175), .CP(clk), .RN(n6589), 
        .Q(\registers[24][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][4]  ( .D(n2174), .CP(clk), .RN(n6589), 
        .Q(\registers[24][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][3]  ( .D(n2173), .CP(clk), .RN(n6589), 
        .Q(\registers[24][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][2]  ( .D(n2172), .CP(clk), .RN(n6590), 
        .Q(\registers[24][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][1]  ( .D(n2171), .CP(clk), .RN(n6590), 
        .Q(\registers[24][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][0]  ( .D(n2170), .CP(clk), .RN(n6590), 
        .Q(\registers[24][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][31]  ( .D(n2169), .CP(clk), .RN(n6593), 
        .Q(\registers[23][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][30]  ( .D(n2168), .CP(clk), .RN(n6593), 
        .Q(\registers[23][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][29]  ( .D(n2167), .CP(clk), .RN(n6593), 
        .Q(\registers[23][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][28]  ( .D(n2166), .CP(clk), .RN(n6593), 
        .Q(\registers[23][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][27]  ( .D(n2165), .CP(clk), .RN(n6594), 
        .Q(\registers[23][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][26]  ( .D(n2164), .CP(clk), .RN(n6594), 
        .Q(\registers[23][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][25]  ( .D(n2163), .CP(clk), .RN(n6594), 
        .Q(\registers[23][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][24]  ( .D(n2162), .CP(clk), .RN(n6594), 
        .Q(\registers[23][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][23]  ( .D(n2161), .CP(clk), .RN(n6592), 
        .Q(\registers[23][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][22]  ( .D(n2160), .CP(clk), .RN(n6595), 
        .Q(\registers[23][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][21]  ( .D(n2159), .CP(clk), .RN(n6595), 
        .Q(\registers[23][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][20]  ( .D(n2158), .CP(clk), .RN(n6593), 
        .Q(\registers[23][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][19]  ( .D(n2157), .CP(clk), .RN(n6593), 
        .Q(\registers[23][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][18]  ( .D(n2156), .CP(clk), .RN(n6592), 
        .Q(\registers[23][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][17]  ( .D(n2155), .CP(clk), .RN(n6592), 
        .Q(\registers[23][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][16]  ( .D(n2154), .CP(clk), .RN(n6592), 
        .Q(\registers[23][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][15]  ( .D(n2153), .CP(clk), .RN(n6592), 
        .Q(\registers[23][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][14]  ( .D(n2152), .CP(clk), .RN(n6592), 
        .Q(\registers[23][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][13]  ( .D(n2151), .CP(clk), .RN(n6592), 
        .Q(\registers[23][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][12]  ( .D(n2150), .CP(clk), .RN(n6592), 
        .Q(\registers[23][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][11]  ( .D(n2149), .CP(clk), .RN(n6592), 
        .Q(\registers[23][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][10]  ( .D(n2148), .CP(clk), .RN(n6593), 
        .Q(\registers[23][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][9]  ( .D(n2147), .CP(clk), .RN(n6593), 
        .Q(\registers[23][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][8]  ( .D(n2146), .CP(clk), .RN(n6593), 
        .Q(\registers[23][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][7]  ( .D(n2145), .CP(clk), .RN(n6591), 
        .Q(\registers[23][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][6]  ( .D(n2144), .CP(clk), .RN(n6591), 
        .Q(\registers[23][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][5]  ( .D(n2143), .CP(clk), .RN(n6591), 
        .Q(\registers[23][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][4]  ( .D(n2142), .CP(clk), .RN(n6591), 
        .Q(\registers[23][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][3]  ( .D(n2141), .CP(clk), .RN(n6591), 
        .Q(\registers[23][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][2]  ( .D(n2140), .CP(clk), .RN(n6591), 
        .Q(\registers[23][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][1]  ( .D(n2139), .CP(clk), .RN(n6591), 
        .Q(\registers[23][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][0]  ( .D(n2138), .CP(clk), .RN(n6591), 
        .Q(\registers[23][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][31]  ( .D(n2137), .CP(clk), .RN(n6596), 
        .Q(\registers[22][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][30]  ( .D(n2136), .CP(clk), .RN(n6597), 
        .Q(\registers[22][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][29]  ( .D(n2135), .CP(clk), .RN(n6597), 
        .Q(\registers[22][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][28]  ( .D(n2134), .CP(clk), .RN(n6597), 
        .Q(\registers[22][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][27]  ( .D(n2133), .CP(clk), .RN(n6597), 
        .Q(\registers[22][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][26]  ( .D(n2132), .CP(clk), .RN(n6596), 
        .Q(\registers[22][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][25]  ( .D(n2131), .CP(clk), .RN(n6596), 
        .Q(\registers[22][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][24]  ( .D(n2130), .CP(clk), .RN(n6596), 
        .Q(\registers[22][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][23]  ( .D(n2129), .CP(clk), .RN(n6595), 
        .Q(\registers[22][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][22]  ( .D(n2128), .CP(clk), .RN(n6595), 
        .Q(\registers[22][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][21]  ( .D(n2127), .CP(clk), .RN(n6593), 
        .Q(\registers[22][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][20]  ( .D(n2126), .CP(clk), .RN(n6593), 
        .Q(\registers[22][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][19]  ( .D(n2125), .CP(clk), .RN(n6593), 
        .Q(\registers[22][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][18]  ( .D(n2124), .CP(clk), .RN(n6597), 
        .Q(\registers[22][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][17]  ( .D(n2123), .CP(clk), .RN(n6597), 
        .Q(\registers[22][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][16]  ( .D(n2122), .CP(clk), .RN(n6597), 
        .Q(\registers[22][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][15]  ( .D(n2121), .CP(clk), .RN(n6594), 
        .Q(\registers[22][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][14]  ( .D(n2120), .CP(clk), .RN(n6594), 
        .Q(\registers[22][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][13]  ( .D(n2119), .CP(clk), .RN(n6594), 
        .Q(\registers[22][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][12]  ( .D(n2118), .CP(clk), .RN(n6594), 
        .Q(\registers[22][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][11]  ( .D(n2117), .CP(clk), .RN(n6594), 
        .Q(\registers[22][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][10]  ( .D(n2116), .CP(clk), .RN(n6594), 
        .Q(\registers[22][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][9]  ( .D(n2115), .CP(clk), .RN(n6594), 
        .Q(\registers[22][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][8]  ( .D(n2114), .CP(clk), .RN(n6594), 
        .Q(\registers[22][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][7]  ( .D(n2113), .CP(clk), .RN(n6586), 
        .Q(\registers[22][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][6]  ( .D(n2112), .CP(clk), .RN(n6538), 
        .Q(\registers[22][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][5]  ( .D(n2111), .CP(clk), .RN(n6538), 
        .Q(\registers[22][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][4]  ( .D(n2110), .CP(clk), .RN(n6538), 
        .Q(\registers[22][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][3]  ( .D(n2109), .CP(clk), .RN(n6538), 
        .Q(\registers[22][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][2]  ( .D(n2108), .CP(clk), .RN(n6538), 
        .Q(\registers[22][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][1]  ( .D(n2107), .CP(clk), .RN(n6538), 
        .Q(\registers[22][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][0]  ( .D(n2106), .CP(clk), .RN(n6538), 
        .Q(\registers[22][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][31]  ( .D(n2105), .CP(clk), .RN(n6541), 
        .Q(\registers[21][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][30]  ( .D(n2104), .CP(clk), .RN(n6542), 
        .Q(\registers[21][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][29]  ( .D(n2103), .CP(clk), .RN(n6541), 
        .Q(\registers[21][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][28]  ( .D(n2102), .CP(clk), .RN(n6542), 
        .Q(\registers[21][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][27]  ( .D(n2101), .CP(clk), .RN(n6541), 
        .Q(\registers[21][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][26]  ( .D(n2100), .CP(clk), .RN(n6540), 
        .Q(\registers[21][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][25]  ( .D(n2099), .CP(clk), .RN(n6540), 
        .Q(\registers[21][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][24]  ( .D(n2098), .CP(clk), .RN(n6539), 
        .Q(\registers[21][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][23]  ( .D(n2097), .CP(clk), .RN(n6539), 
        .Q(\registers[21][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][22]  ( .D(n2096), .CP(clk), .RN(n6573), 
        .Q(\registers[21][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][21]  ( .D(n2095), .CP(clk), .RN(n6573), 
        .Q(\registers[21][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][20]  ( .D(n2094), .CP(clk), .RN(n6572), 
        .Q(\registers[21][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][19]  ( .D(n2093), .CP(clk), .RN(n6572), 
        .Q(\registers[21][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][18]  ( .D(n2092), .CP(clk), .RN(n6569), 
        .Q(\registers[21][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][17]  ( .D(n2091), .CP(clk), .RN(n6569), 
        .Q(\registers[21][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][16]  ( .D(n2090), .CP(clk), .RN(n6569), 
        .Q(\registers[21][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][15]  ( .D(n2089), .CP(clk), .RN(n6569), 
        .Q(\registers[21][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][14]  ( .D(n2088), .CP(clk), .RN(n6569), 
        .Q(\registers[21][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][13]  ( .D(n2087), .CP(clk), .RN(n6569), 
        .Q(\registers[21][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][12]  ( .D(n2086), .CP(clk), .RN(n6569), 
        .Q(\registers[21][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][11]  ( .D(n2085), .CP(clk), .RN(n6569), 
        .Q(\registers[21][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][10]  ( .D(n2084), .CP(clk), .RN(n6572), 
        .Q(\registers[21][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][9]  ( .D(n2083), .CP(clk), .RN(n6572), 
        .Q(\registers[21][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][8]  ( .D(n2082), .CP(clk), .RN(n6572), 
        .Q(\registers[21][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][7]  ( .D(n2081), .CP(clk), .RN(n6570), 
        .Q(\registers[21][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][6]  ( .D(n2080), .CP(clk), .RN(n6570), 
        .Q(\registers[21][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][5]  ( .D(n2079), .CP(clk), .RN(n6570), 
        .Q(\registers[21][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][4]  ( .D(n2078), .CP(clk), .RN(n6570), 
        .Q(\registers[21][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][3]  ( .D(n2077), .CP(clk), .RN(n6570), 
        .Q(\registers[21][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][2]  ( .D(n2076), .CP(clk), .RN(n6570), 
        .Q(\registers[21][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][1]  ( .D(n2075), .CP(clk), .RN(n6570), 
        .Q(\registers[21][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][0]  ( .D(n2074), .CP(clk), .RN(n6570), 
        .Q(\registers[21][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][31]  ( .D(n2073), .CP(clk), .RN(n6574), 
        .Q(\registers[20][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][30]  ( .D(n2072), .CP(clk), .RN(n6571), 
        .Q(\registers[20][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][29]  ( .D(n2071), .CP(clk), .RN(n6571), 
        .Q(\registers[20][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][28]  ( .D(n2070), .CP(clk), .RN(n6571), 
        .Q(\registers[20][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][27]  ( .D(n2069), .CP(clk), .RN(n6570), 
        .Q(\registers[20][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][26]  ( .D(n2068), .CP(clk), .RN(n6570), 
        .Q(\registers[20][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][25]  ( .D(n2067), .CP(clk), .RN(n6569), 
        .Q(\registers[20][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][24]  ( .D(n2066), .CP(clk), .RN(n6569), 
        .Q(\registers[20][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][23]  ( .D(n2065), .CP(clk), .RN(n6574), 
        .Q(\registers[20][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][22]  ( .D(n2064), .CP(clk), .RN(n6574), 
        .Q(\registers[20][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][21]  ( .D(n2063), .CP(clk), .RN(n6573), 
        .Q(\registers[20][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][20]  ( .D(n2062), .CP(clk), .RN(n6574), 
        .Q(\registers[20][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][19]  ( .D(n2061), .CP(clk), .RN(n6574), 
        .Q(\registers[20][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][18]  ( .D(n2060), .CP(clk), .RN(n6573), 
        .Q(\registers[20][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][17]  ( .D(n2059), .CP(clk), .RN(n6573), 
        .Q(\registers[20][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][16]  ( .D(n2058), .CP(clk), .RN(n6573), 
        .Q(\registers[20][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][15]  ( .D(n2057), .CP(clk), .RN(n6573), 
        .Q(\registers[20][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][14]  ( .D(n2056), .CP(clk), .RN(n6573), 
        .Q(\registers[20][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][13]  ( .D(n2055), .CP(clk), .RN(n6573), 
        .Q(\registers[20][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][12]  ( .D(n2054), .CP(clk), .RN(n6573), 
        .Q(\registers[20][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][11]  ( .D(n2053), .CP(clk), .RN(n6573), 
        .Q(\registers[20][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][10]  ( .D(n2052), .CP(clk), .RN(n6574), 
        .Q(\registers[20][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][9]  ( .D(n2051), .CP(clk), .RN(n6574), 
        .Q(\registers[20][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][8]  ( .D(n2050), .CP(clk), .RN(n6574), 
        .Q(\registers[20][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][7]  ( .D(n2049), .CP(clk), .RN(n6576), 
        .Q(\registers[20][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][6]  ( .D(n2048), .CP(clk), .RN(n6576), 
        .Q(\registers[20][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][5]  ( .D(n2047), .CP(clk), .RN(n6576), 
        .Q(\registers[20][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][4]  ( .D(n2046), .CP(clk), .RN(n6576), 
        .Q(\registers[20][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][3]  ( .D(n2045), .CP(clk), .RN(n6576), 
        .Q(\registers[20][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][2]  ( .D(n2044), .CP(clk), .RN(n6576), 
        .Q(\registers[20][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][1]  ( .D(n2043), .CP(clk), .RN(n6576), 
        .Q(\registers[20][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][0]  ( .D(n2042), .CP(clk), .RN(n6576), 
        .Q(\registers[20][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][31]  ( .D(n2041), .CP(clk), .RN(n6588), 
        .Q(\registers[19][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][30]  ( .D(n2040), .CP(clk), .RN(n6588), 
        .Q(\registers[19][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][29]  ( .D(n2039), .CP(clk), .RN(n6588), 
        .Q(\registers[19][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][28]  ( .D(n2038), .CP(clk), .RN(n6588), 
        .Q(\registers[19][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][27]  ( .D(n2037), .CP(clk), .RN(n6578), 
        .Q(\registers[19][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][26]  ( .D(n2036), .CP(clk), .RN(n6577), 
        .Q(\registers[19][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][25]  ( .D(n2035), .CP(clk), .RN(n6577), 
        .Q(\registers[19][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][24]  ( .D(n2034), .CP(clk), .RN(n6577), 
        .Q(\registers[19][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][23]  ( .D(n2033), .CP(clk), .RN(n6577), 
        .Q(\registers[19][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][22]  ( .D(n2032), .CP(clk), .RN(n6577), 
        .Q(\registers[19][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][21]  ( .D(n2031), .CP(clk), .RN(n6577), 
        .Q(\registers[19][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][20]  ( .D(n2030), .CP(clk), .RN(n6577), 
        .Q(\registers[19][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][19]  ( .D(n2029), .CP(clk), .RN(n6587), 
        .Q(\registers[19][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][18]  ( .D(n2028), .CP(clk), .RN(n6587), 
        .Q(\registers[19][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][17]  ( .D(n2027), .CP(clk), .RN(n6587), 
        .Q(\registers[19][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][16]  ( .D(n2026), .CP(clk), .RN(n6587), 
        .Q(\registers[19][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][15]  ( .D(n2025), .CP(clk), .RN(n6587), 
        .Q(\registers[19][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][14]  ( .D(n2024), .CP(clk), .RN(n6587), 
        .Q(\registers[19][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][13]  ( .D(n2023), .CP(clk), .RN(n6587), 
        .Q(\registers[19][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][12]  ( .D(n2022), .CP(clk), .RN(n6587), 
        .Q(\registers[19][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][11]  ( .D(n2021), .CP(clk), .RN(n6587), 
        .Q(\registers[19][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][10]  ( .D(n2020), .CP(clk), .RN(n6587), 
        .Q(\registers[19][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][9]  ( .D(n2019), .CP(clk), .RN(n6587), 
        .Q(\registers[19][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][8]  ( .D(n2018), .CP(clk), .RN(n6587), 
        .Q(\registers[19][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][7]  ( .D(n2017), .CP(clk), .RN(n6571), 
        .Q(\registers[19][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][6]  ( .D(n2016), .CP(clk), .RN(n6571), 
        .Q(\registers[19][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][5]  ( .D(n2015), .CP(clk), .RN(n6571), 
        .Q(\registers[19][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][4]  ( .D(n2014), .CP(clk), .RN(n6571), 
        .Q(\registers[19][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][3]  ( .D(n2013), .CP(clk), .RN(n6571), 
        .Q(\registers[19][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][2]  ( .D(n2012), .CP(clk), .RN(n6571), 
        .Q(\registers[19][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][1]  ( .D(n2011), .CP(clk), .RN(n6571), 
        .Q(\registers[19][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][0]  ( .D(n2010), .CP(clk), .RN(n6571), 
        .Q(\registers[19][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][31]  ( .D(n2009), .CP(clk), .RN(n6577), 
        .Q(\registers[18][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][30]  ( .D(n2008), .CP(clk), .RN(n6577), 
        .Q(\registers[18][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][29]  ( .D(n2007), .CP(clk), .RN(n6577), 
        .Q(\registers[18][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][28]  ( .D(n2006), .CP(clk), .RN(n6578), 
        .Q(\registers[18][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][27]  ( .D(n2005), .CP(clk), .RN(n6578), 
        .Q(\registers[18][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][26]  ( .D(n2004), .CP(clk), .RN(n6578), 
        .Q(\registers[18][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][25]  ( .D(n2003), .CP(clk), .RN(n6577), 
        .Q(\registers[18][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][24]  ( .D(n2002), .CP(clk), .RN(n6577), 
        .Q(\registers[18][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][23]  ( .D(n2001), .CP(clk), .RN(n6574), 
        .Q(\registers[18][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][22]  ( .D(n2000), .CP(clk), .RN(n6574), 
        .Q(\registers[18][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][21]  ( .D(n1999), .CP(clk), .RN(n6574), 
        .Q(\registers[18][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][20]  ( .D(n1998), .CP(clk), .RN(n6573), 
        .Q(\registers[18][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][19]  ( .D(n1997), .CP(clk), .RN(n6572), 
        .Q(\registers[18][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][18]  ( .D(n1996), .CP(clk), .RN(n6572), 
        .Q(\registers[18][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][17]  ( .D(n1995), .CP(clk), .RN(n6572), 
        .Q(\registers[18][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][16]  ( .D(n1994), .CP(clk), .RN(n6574), 
        .Q(\registers[18][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][15]  ( .D(n1993), .CP(clk), .RN(n6548), 
        .Q(\registers[18][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][14]  ( .D(n1992), .CP(clk), .RN(n6550), 
        .Q(\registers[18][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][13]  ( .D(n1991), .CP(clk), .RN(n6540), 
        .Q(\registers[18][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][12]  ( .D(n1990), .CP(clk), .RN(n6540), 
        .Q(\registers[18][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][11]  ( .D(n1989), .CP(clk), .RN(n6540), 
        .Q(\registers[18][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][10]  ( .D(n1988), .CP(clk), .RN(n6542), 
        .Q(\registers[18][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][9]  ( .D(n1987), .CP(clk), .RN(n6542), 
        .Q(\registers[18][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][8]  ( .D(n1986), .CP(clk), .RN(n6542), 
        .Q(\registers[18][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][7]  ( .D(n1985), .CP(clk), .RN(n6542), 
        .Q(\registers[18][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][6]  ( .D(n1984), .CP(clk), .RN(n6542), 
        .Q(\registers[18][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][5]  ( .D(n1983), .CP(clk), .RN(n6542), 
        .Q(\registers[18][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][4]  ( .D(n1982), .CP(clk), .RN(n6542), 
        .Q(\registers[18][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][3]  ( .D(n1981), .CP(clk), .RN(n6542), 
        .Q(\registers[18][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][2]  ( .D(n1980), .CP(clk), .RN(n6552), 
        .Q(\registers[18][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][1]  ( .D(n1979), .CP(clk), .RN(n6552), 
        .Q(\registers[18][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][0]  ( .D(n1978), .CP(clk), .RN(n6552), 
        .Q(\registers[18][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][31]  ( .D(n1977), .CP(clk), .RN(n6555), 
        .Q(\registers[17][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][30]  ( .D(n1976), .CP(clk), .RN(n6555), 
        .Q(\registers[17][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][29]  ( .D(n1975), .CP(clk), .RN(n6555), 
        .Q(\registers[17][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][28]  ( .D(n1974), .CP(clk), .RN(n6555), 
        .Q(\registers[17][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][27]  ( .D(n1973), .CP(clk), .RN(n6557), 
        .Q(\registers[17][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][26]  ( .D(n1972), .CP(clk), .RN(n6557), 
        .Q(\registers[17][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][25]  ( .D(n1971), .CP(clk), .RN(n6557), 
        .Q(\registers[17][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][24]  ( .D(n1970), .CP(clk), .RN(n6552), 
        .Q(\registers[17][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][23]  ( .D(n1969), .CP(clk), .RN(n6552), 
        .Q(\registers[17][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][22]  ( .D(n1968), .CP(clk), .RN(n6556), 
        .Q(\registers[17][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][21]  ( .D(n1967), .CP(clk), .RN(n6556), 
        .Q(\registers[17][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][20]  ( .D(n1966), .CP(clk), .RN(n6556), 
        .Q(\registers[17][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][19]  ( .D(n1965), .CP(clk), .RN(n6556), 
        .Q(\registers[17][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][18]  ( .D(n1964), .CP(clk), .RN(n6556), 
        .Q(\registers[17][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][17]  ( .D(n1963), .CP(clk), .RN(n6556), 
        .Q(\registers[17][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][16]  ( .D(n1962), .CP(clk), .RN(n6556), 
        .Q(\registers[17][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][15]  ( .D(n1961), .CP(clk), .RN(n6556), 
        .Q(\registers[17][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][14]  ( .D(n1960), .CP(clk), .RN(n6556), 
        .Q(\registers[17][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][13]  ( .D(n1959), .CP(clk), .RN(n6556), 
        .Q(\registers[17][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][12]  ( .D(n1958), .CP(clk), .RN(n6556), 
        .Q(\registers[17][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][11]  ( .D(n1957), .CP(clk), .RN(n6556), 
        .Q(\registers[17][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][10]  ( .D(n1956), .CP(clk), .RN(n6552), 
        .Q(\registers[17][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][9]  ( .D(n1955), .CP(clk), .RN(n6552), 
        .Q(\registers[17][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][8]  ( .D(n1954), .CP(clk), .RN(n6552), 
        .Q(\registers[17][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][7]  ( .D(n1953), .CP(clk), .RN(n6555), 
        .Q(\registers[17][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][6]  ( .D(n1952), .CP(clk), .RN(n6555), 
        .Q(\registers[17][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][5]  ( .D(n1951), .CP(clk), .RN(n6555), 
        .Q(\registers[17][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][4]  ( .D(n1950), .CP(clk), .RN(n6555), 
        .Q(\registers[17][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][3]  ( .D(n1949), .CP(clk), .RN(n6555), 
        .Q(\registers[17][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][2]  ( .D(n1948), .CP(clk), .RN(n6555), 
        .Q(\registers[17][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][1]  ( .D(n1947), .CP(clk), .RN(n6555), 
        .Q(\registers[17][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][0]  ( .D(n1946), .CP(clk), .RN(n6555), 
        .Q(\registers[17][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][31]  ( .D(n1945), .CP(clk), .RN(n6557), 
        .Q(\registers[16][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][30]  ( .D(n1944), .CP(clk), .RN(n6558), 
        .Q(\registers[16][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][29]  ( .D(n1943), .CP(clk), .RN(n6558), 
        .Q(\registers[16][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][28]  ( .D(n1942), .CP(clk), .RN(n6558), 
        .Q(\registers[16][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][27]  ( .D(n1941), .CP(clk), .RN(n6558), 
        .Q(\registers[16][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][26]  ( .D(n1940), .CP(clk), .RN(n6553), 
        .Q(\registers[16][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][25]  ( .D(n1939), .CP(clk), .RN(n6553), 
        .Q(\registers[16][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][24]  ( .D(n1938), .CP(clk), .RN(n6550), 
        .Q(\registers[16][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][23]  ( .D(n1937), .CP(clk), .RN(n6550), 
        .Q(\registers[16][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][22]  ( .D(n1936), .CP(clk), .RN(n6550), 
        .Q(\registers[16][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][21]  ( .D(n1935), .CP(clk), .RN(n6550), 
        .Q(\registers[16][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][20]  ( .D(n1934), .CP(clk), .RN(n6550), 
        .Q(\registers[16][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][19]  ( .D(n1933), .CP(clk), .RN(n6557), 
        .Q(\registers[16][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][18]  ( .D(n1932), .CP(clk), .RN(n6557), 
        .Q(\registers[16][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][17]  ( .D(n1931), .CP(clk), .RN(n6557), 
        .Q(\registers[16][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][16]  ( .D(n1930), .CP(clk), .RN(n6557), 
        .Q(\registers[16][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][15]  ( .D(n1929), .CP(clk), .RN(n6553), 
        .Q(\registers[16][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][14]  ( .D(n1928), .CP(clk), .RN(n6553), 
        .Q(\registers[16][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][13]  ( .D(n1927), .CP(clk), .RN(n6553), 
        .Q(\registers[16][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][12]  ( .D(n1926), .CP(clk), .RN(n6553), 
        .Q(\registers[16][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][11]  ( .D(n1925), .CP(clk), .RN(n6553), 
        .Q(\registers[16][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][10]  ( .D(n1924), .CP(clk), .RN(n6553), 
        .Q(\registers[16][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][9]  ( .D(n1923), .CP(clk), .RN(n6553), 
        .Q(\registers[16][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][8]  ( .D(n1922), .CP(clk), .RN(n6553), 
        .Q(\registers[16][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][7]  ( .D(n1921), .CP(clk), .RN(n6554), 
        .Q(\registers[16][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][6]  ( .D(n1920), .CP(clk), .RN(n6554), 
        .Q(\registers[16][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][5]  ( .D(n1919), .CP(clk), .RN(n6554), 
        .Q(\registers[16][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][4]  ( .D(n1918), .CP(clk), .RN(n6554), 
        .Q(\registers[16][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][3]  ( .D(n1917), .CP(clk), .RN(n6554), 
        .Q(\registers[16][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][2]  ( .D(n1916), .CP(clk), .RN(n6554), 
        .Q(\registers[16][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][1]  ( .D(n1915), .CP(clk), .RN(n6554), 
        .Q(\registers[16][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][0]  ( .D(n1914), .CP(clk), .RN(n6554), 
        .Q(\registers[16][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][31]  ( .D(n1849), .CP(clk), .RN(n6559), 
        .Q(\registers[13][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][30]  ( .D(n1848), .CP(clk), .RN(n6559), 
        .Q(\registers[13][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][29]  ( .D(n1847), .CP(clk), .RN(n6559), 
        .Q(\registers[13][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][28]  ( .D(n1846), .CP(clk), .RN(n6559), 
        .Q(\registers[13][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][27]  ( .D(n1845), .CP(clk), .RN(n6561), 
        .Q(\registers[13][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][26]  ( .D(n1844), .CP(clk), .RN(n6561), 
        .Q(\registers[13][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][25]  ( .D(n1843), .CP(clk), .RN(n6561), 
        .Q(\registers[13][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][24]  ( .D(n1842), .CP(clk), .RN(n6561), 
        .Q(\registers[13][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][23]  ( .D(n1841), .CP(clk), .RN(n6560), 
        .Q(\registers[13][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][22]  ( .D(n1840), .CP(clk), .RN(n6560), 
        .Q(\registers[13][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][21]  ( .D(n1839), .CP(clk), .RN(n6560), 
        .Q(\registers[13][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][20]  ( .D(n1838), .CP(clk), .RN(n6560), 
        .Q(\registers[13][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][19]  ( .D(n1837), .CP(clk), .RN(n6557), 
        .Q(\registers[13][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][18]  ( .D(n1836), .CP(clk), .RN(n6557), 
        .Q(\registers[13][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][17]  ( .D(n1835), .CP(clk), .RN(n6557), 
        .Q(\registers[13][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][16]  ( .D(n1834), .CP(clk), .RN(n6557), 
        .Q(\registers[13][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][15]  ( .D(n1833), .CP(clk), .RN(n6562), 
        .Q(\registers[13][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][14]  ( .D(n1832), .CP(clk), .RN(n6558), 
        .Q(\registers[13][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][13]  ( .D(n1831), .CP(clk), .RN(n6558), 
        .Q(\registers[13][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][12]  ( .D(n1830), .CP(clk), .RN(n6558), 
        .Q(\registers[13][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][11]  ( .D(n1829), .CP(clk), .RN(n6561), 
        .Q(\registers[13][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][10]  ( .D(n1828), .CP(clk), .RN(n6561), 
        .Q(\registers[13][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][9]  ( .D(n1827), .CP(clk), .RN(n6561), 
        .Q(\registers[13][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][8]  ( .D(n1826), .CP(clk), .RN(n6561), 
        .Q(\registers[13][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][7]  ( .D(n1825), .CP(clk), .RN(n6561), 
        .Q(\registers[13][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][6]  ( .D(n1824), .CP(clk), .RN(n6561), 
        .Q(\registers[13][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][5]  ( .D(n1823), .CP(clk), .RN(n6561), 
        .Q(\registers[13][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][4]  ( .D(n1822), .CP(clk), .RN(n6561), 
        .Q(\registers[13][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][3]  ( .D(n1821), .CP(clk), .RN(n6541), 
        .Q(\registers[13][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][2]  ( .D(n1820), .CP(clk), .RN(n6539), 
        .Q(\registers[13][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][1]  ( .D(n1819), .CP(clk), .RN(n6539), 
        .Q(\registers[13][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][0]  ( .D(n1818), .CP(clk), .RN(n6539), 
        .Q(\registers[13][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][31]  ( .D(n1817), .CP(clk), .RN(n6539), 
        .Q(\registers[12][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][30]  ( .D(n1816), .CP(clk), .RN(n6539), 
        .Q(\registers[12][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][29]  ( .D(n1815), .CP(clk), .RN(n6539), 
        .Q(\registers[12][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][28]  ( .D(n1814), .CP(clk), .RN(n6542), 
        .Q(\registers[12][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][27]  ( .D(n1813), .CP(clk), .RN(n6542), 
        .Q(\registers[12][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][26]  ( .D(n1812), .CP(clk), .RN(n6541), 
        .Q(\registers[12][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][25]  ( .D(n1811), .CP(clk), .RN(n6540), 
        .Q(\registers[12][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][24]  ( .D(n1810), .CP(clk), .RN(n6540), 
        .Q(\registers[12][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][23]  ( .D(n1809), .CP(clk), .RN(n6539), 
        .Q(\registers[12][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][22]  ( .D(n1808), .CP(clk), .RN(n6539), 
        .Q(\registers[12][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][21]  ( .D(n1807), .CP(clk), .RN(n6539), 
        .Q(\registers[12][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][20]  ( .D(n1806), .CP(clk), .RN(n6538), 
        .Q(\registers[12][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][19]  ( .D(n1805), .CP(clk), .RN(n6544), 
        .Q(\registers[12][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][18]  ( .D(n1804), .CP(clk), .RN(n6544), 
        .Q(\registers[12][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][17]  ( .D(n1803), .CP(clk), .RN(n6544), 
        .Q(\registers[12][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][16]  ( .D(n1802), .CP(clk), .RN(n6544), 
        .Q(\registers[12][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][15]  ( .D(n1801), .CP(clk), .RN(n6544), 
        .Q(\registers[12][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][14]  ( .D(n1800), .CP(clk), .RN(n6544), 
        .Q(\registers[12][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][13]  ( .D(n1799), .CP(clk), .RN(n6544), 
        .Q(\registers[12][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][12]  ( .D(n1798), .CP(clk), .RN(n6544), 
        .Q(\registers[12][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][11]  ( .D(n1797), .CP(clk), .RN(n6545), 
        .Q(\registers[12][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][10]  ( .D(n1796), .CP(clk), .RN(n6545), 
        .Q(\registers[12][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][9]  ( .D(n1795), .CP(clk), .RN(n6545), 
        .Q(\registers[12][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][8]  ( .D(n1794), .CP(clk), .RN(n6545), 
        .Q(\registers[12][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][7]  ( .D(n1793), .CP(clk), .RN(n6546), 
        .Q(\registers[12][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][6]  ( .D(n1792), .CP(clk), .RN(n6546), 
        .Q(\registers[12][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][5]  ( .D(n1791), .CP(clk), .RN(n6546), 
        .Q(\registers[12][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][4]  ( .D(n1790), .CP(clk), .RN(n6546), 
        .Q(\registers[12][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][3]  ( .D(n1789), .CP(clk), .RN(n6546), 
        .Q(\registers[12][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][2]  ( .D(n1788), .CP(clk), .RN(n6546), 
        .Q(\registers[12][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][1]  ( .D(n1787), .CP(clk), .RN(n6546), 
        .Q(\registers[12][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][0]  ( .D(n1786), .CP(clk), .RN(n6546), 
        .Q(\registers[12][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][31]  ( .D(n1785), .CP(clk), .RN(n6550), 
        .Q(\registers[11][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][30]  ( .D(n1784), .CP(clk), .RN(n6550), 
        .Q(\registers[11][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][29]  ( .D(n1783), .CP(clk), .RN(n6550), 
        .Q(\registers[11][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][28]  ( .D(n1782), .CP(clk), .RN(n6550), 
        .Q(\registers[11][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][27]  ( .D(n1781), .CP(clk), .RN(n6549), 
        .Q(\registers[11][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][26]  ( .D(n1780), .CP(clk), .RN(n6549), 
        .Q(\registers[11][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][25]  ( .D(n1779), .CP(clk), .RN(n6549), 
        .Q(\registers[11][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][24]  ( .D(n1778), .CP(clk), .RN(n6549), 
        .Q(\registers[11][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][23]  ( .D(n1777), .CP(clk), .RN(n6545), 
        .Q(\registers[11][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][22]  ( .D(n1776), .CP(clk), .RN(n6545), 
        .Q(\registers[11][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][21]  ( .D(n1775), .CP(clk), .RN(n6545), 
        .Q(\registers[11][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][20]  ( .D(n1774), .CP(clk), .RN(n6545), 
        .Q(\registers[11][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][19]  ( .D(n1773), .CP(clk), .RN(n6552), 
        .Q(\registers[11][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][18]  ( .D(n1772), .CP(clk), .RN(n6548), 
        .Q(\registers[11][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][17]  ( .D(n1771), .CP(clk), .RN(n6548), 
        .Q(\registers[11][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][16]  ( .D(n1770), .CP(clk), .RN(n6548), 
        .Q(\registers[11][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][15]  ( .D(n1769), .CP(clk), .RN(n6541), 
        .Q(\registers[11][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][14]  ( .D(n1768), .CP(clk), .RN(n6541), 
        .Q(\registers[11][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][13]  ( .D(n1767), .CP(clk), .RN(n6541), 
        .Q(\registers[11][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][12]  ( .D(n1766), .CP(clk), .RN(n6541), 
        .Q(\registers[11][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][11]  ( .D(n1765), .CP(clk), .RN(n6541), 
        .Q(\registers[11][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][10]  ( .D(n1764), .CP(clk), .RN(n6541), 
        .Q(\registers[11][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][9]  ( .D(n1763), .CP(clk), .RN(n6541), 
        .Q(\registers[11][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][8]  ( .D(n1762), .CP(clk), .RN(n6550), 
        .Q(\registers[11][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][7]  ( .D(n1761), .CP(clk), .RN(n6551), 
        .Q(\registers[11][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][6]  ( .D(n1760), .CP(clk), .RN(n6551), 
        .Q(\registers[11][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][5]  ( .D(n1759), .CP(clk), .RN(n6551), 
        .Q(\registers[11][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][4]  ( .D(n1758), .CP(clk), .RN(n6551), 
        .Q(\registers[11][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][3]  ( .D(n1757), .CP(clk), .RN(n6551), 
        .Q(\registers[11][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][2]  ( .D(n1756), .CP(clk), .RN(n6551), 
        .Q(\registers[11][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][1]  ( .D(n1755), .CP(clk), .RN(n6551), 
        .Q(\registers[11][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][0]  ( .D(n1754), .CP(clk), .RN(n6551), 
        .Q(\registers[11][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][31]  ( .D(n1753), .CP(clk), .RN(n6551), 
        .Q(\registers[10][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][30]  ( .D(n1752), .CP(clk), .RN(n6551), 
        .Q(\registers[10][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][29]  ( .D(n1751), .CP(clk), .RN(n6551), 
        .Q(\registers[10][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][28]  ( .D(n1750), .CP(clk), .RN(n6563), 
        .Q(\registers[10][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][27]  ( .D(n1749), .CP(clk), .RN(n6563), 
        .Q(\registers[10][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][26]  ( .D(n1748), .CP(clk), .RN(n6563), 
        .Q(\registers[10][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][25]  ( .D(n1747), .CP(clk), .RN(n6563), 
        .Q(\registers[10][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][24]  ( .D(n1746), .CP(clk), .RN(n6549), 
        .Q(\registers[10][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][23]  ( .D(n1745), .CP(clk), .RN(n6549), 
        .Q(\registers[10][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][22]  ( .D(n1744), .CP(clk), .RN(n6549), 
        .Q(\registers[10][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][21]  ( .D(n1743), .CP(clk), .RN(n6549), 
        .Q(\registers[10][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][20]  ( .D(n1742), .CP(clk), .RN(n6549), 
        .Q(\registers[10][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][19]  ( .D(n1741), .CP(clk), .RN(n6549), 
        .Q(\registers[10][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][18]  ( .D(n1740), .CP(clk), .RN(n6549), 
        .Q(\registers[10][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][17]  ( .D(n1739), .CP(clk), .RN(n6549), 
        .Q(\registers[10][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][16]  ( .D(n1738), .CP(clk), .RN(n6564), 
        .Q(\registers[10][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][15]  ( .D(n1737), .CP(clk), .RN(n6564), 
        .Q(\registers[10][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][14]  ( .D(n1736), .CP(clk), .RN(n6564), 
        .Q(\registers[10][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][13]  ( .D(n1735), .CP(clk), .RN(n6564), 
        .Q(\registers[10][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][12]  ( .D(n1734), .CP(clk), .RN(n6559), 
        .Q(\registers[10][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][11]  ( .D(n1733), .CP(clk), .RN(n6559), 
        .Q(\registers[10][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][10]  ( .D(n1732), .CP(clk), .RN(n6559), 
        .Q(\registers[10][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][9]  ( .D(n1731), .CP(clk), .RN(n6559), 
        .Q(\registers[10][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][8]  ( .D(n1730), .CP(clk), .RN(n6559), 
        .Q(\registers[10][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][7]  ( .D(n1729), .CP(clk), .RN(n6559), 
        .Q(\registers[10][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][6]  ( .D(n1728), .CP(clk), .RN(n6559), 
        .Q(\registers[10][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][5]  ( .D(n1727), .CP(clk), .RN(n6559), 
        .Q(\registers[10][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][4]  ( .D(n1726), .CP(clk), .RN(n6540), 
        .Q(\registers[10][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][3]  ( .D(n1725), .CP(clk), .RN(n6540), 
        .Q(\registers[10][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][2]  ( .D(n1724), .CP(clk), .RN(n6540), 
        .Q(\registers[10][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][1]  ( .D(n1723), .CP(clk), .RN(n6540), 
        .Q(\registers[10][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][0]  ( .D(n1722), .CP(clk), .RN(n6540), 
        .Q(\registers[10][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][31]  ( .D(n1657), .CP(clk), .RN(n6545), 
        .Q(\registers[7][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][30]  ( .D(n1656), .CP(clk), .RN(n6545), 
        .Q(\registers[7][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][29]  ( .D(n1655), .CP(clk), .RN(n6545), 
        .Q(\registers[7][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][28]  ( .D(n1654), .CP(clk), .RN(n6545), 
        .Q(\registers[7][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][27]  ( .D(n1653), .CP(clk), .RN(n6546), 
        .Q(\registers[7][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][26]  ( .D(n1652), .CP(clk), .RN(n6546), 
        .Q(\registers[7][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][25]  ( .D(n1651), .CP(clk), .RN(n6546), 
        .Q(\registers[7][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][24]  ( .D(n1650), .CP(clk), .RN(n6546), 
        .Q(\registers[7][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][23]  ( .D(n1649), .CP(clk), .RN(n6537), 
        .Q(\registers[7][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][22]  ( .D(n1648), .CP(clk), .RN(n6565), 
        .Q(\registers[7][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][21]  ( .D(n1647), .CP(clk), .RN(n6565), 
        .Q(\registers[7][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][20]  ( .D(n1646), .CP(clk), .RN(n6565), 
        .Q(\registers[7][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][19]  ( .D(n1645), .CP(clk), .RN(n6565), 
        .Q(\registers[7][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][18]  ( .D(n1644), .CP(clk), .RN(n6562), 
        .Q(\registers[7][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][17]  ( .D(n1643), .CP(clk), .RN(n6562), 
        .Q(\registers[7][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][16]  ( .D(n1642), .CP(clk), .RN(n6562), 
        .Q(\registers[7][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][15]  ( .D(n1641), .CP(clk), .RN(n6558), 
        .Q(\registers[7][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][14]  ( .D(n1640), .CP(clk), .RN(n6558), 
        .Q(\registers[7][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][13]  ( .D(n1639), .CP(clk), .RN(n6558), 
        .Q(\registers[7][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][12]  ( .D(n1638), .CP(clk), .RN(n6558), 
        .Q(\registers[7][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][11]  ( .D(n1637), .CP(clk), .RN(n6564), 
        .Q(\registers[7][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][10]  ( .D(n1636), .CP(clk), .RN(n6564), 
        .Q(\registers[7][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][9]  ( .D(n1635), .CP(clk), .RN(n6564), .Q(
        \registers[7][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][8]  ( .D(n1634), .CP(clk), .RN(n6564), .Q(
        \registers[7][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][7]  ( .D(n1633), .CP(clk), .RN(n6562), .Q(
        \registers[7][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][6]  ( .D(n1632), .CP(clk), .RN(n6562), .Q(
        \registers[7][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][5]  ( .D(n1631), .CP(clk), .RN(n6562), .Q(
        \registers[7][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][4]  ( .D(n1630), .CP(clk), .RN(n6562), .Q(
        \registers[7][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][3]  ( .D(n1629), .CP(clk), .RN(n6562), .Q(
        \registers[7][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][2]  ( .D(n1628), .CP(clk), .RN(n6562), .Q(
        \registers[7][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][1]  ( .D(n1627), .CP(clk), .RN(n6562), .Q(
        \registers[7][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][0]  ( .D(n1626), .CP(clk), .RN(n6562), .Q(
        \registers[7][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][31]  ( .D(n1625), .CP(clk), .RN(n6567), 
        .Q(\registers[6][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][30]  ( .D(n1624), .CP(clk), .RN(n6567), 
        .Q(\registers[6][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][29]  ( .D(n1623), .CP(clk), .RN(n6567), 
        .Q(\registers[6][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][28]  ( .D(n1622), .CP(clk), .RN(n6567), 
        .Q(\registers[6][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][27]  ( .D(n1621), .CP(clk), .RN(n6568), 
        .Q(\registers[6][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][26]  ( .D(n1620), .CP(clk), .RN(n6568), 
        .Q(\registers[6][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][25]  ( .D(n1619), .CP(clk), .RN(n6568), 
        .Q(\registers[6][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][24]  ( .D(n1618), .CP(clk), .RN(n6566), 
        .Q(\registers[6][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][23]  ( .D(n1617), .CP(clk), .RN(n6566), 
        .Q(\registers[6][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][22]  ( .D(n1616), .CP(clk), .RN(n6566), 
        .Q(\registers[6][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][21]  ( .D(n1615), .CP(clk), .RN(n6566), 
        .Q(\registers[6][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][20]  ( .D(n1614), .CP(clk), .RN(n6566), 
        .Q(\registers[6][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][19]  ( .D(n1613), .CP(clk), .RN(n6598), 
        .Q(\registers[6][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][18]  ( .D(n1612), .CP(clk), .RN(n6597), 
        .Q(\registers[6][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][17]  ( .D(n1611), .CP(clk), .RN(n6597), 
        .Q(\registers[6][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][16]  ( .D(n1610), .CP(clk), .RN(n6597), 
        .Q(\registers[6][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][15]  ( .D(n1609), .CP(clk), .RN(n6596), 
        .Q(\registers[6][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][14]  ( .D(n1608), .CP(clk), .RN(n6596), 
        .Q(\registers[6][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][13]  ( .D(n1607), .CP(clk), .RN(n6596), 
        .Q(\registers[6][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][12]  ( .D(n1606), .CP(clk), .RN(n6596), 
        .Q(\registers[6][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][11]  ( .D(n1605), .CP(clk), .RN(n6596), 
        .Q(\registers[6][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][10]  ( .D(n1604), .CP(clk), .RN(n6596), 
        .Q(\registers[6][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][9]  ( .D(n1603), .CP(clk), .RN(n6596), .Q(
        \registers[6][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][8]  ( .D(n1602), .CP(clk), .RN(n6596), .Q(
        \registers[6][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][7]  ( .D(n1601), .CP(clk), .RN(n6595), .Q(
        \registers[6][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][6]  ( .D(n1600), .CP(clk), .RN(n6595), .Q(
        \registers[6][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][5]  ( .D(n1599), .CP(clk), .RN(n6595), .Q(
        \registers[6][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][4]  ( .D(n1598), .CP(clk), .RN(n6595), .Q(
        \registers[6][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][3]  ( .D(n1597), .CP(clk), .RN(n6595), .Q(
        \registers[6][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][2]  ( .D(n1596), .CP(clk), .RN(n6595), .Q(
        \registers[6][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][1]  ( .D(n1595), .CP(clk), .RN(n6595), .Q(
        \registers[6][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][0]  ( .D(n1594), .CP(clk), .RN(n6595), .Q(
        \registers[6][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][31]  ( .D(n1593), .CP(clk), .RN(n6537), 
        .Q(\registers[5][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][30]  ( .D(n1592), .CP(clk), .RN(n6537), 
        .Q(\registers[5][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][29]  ( .D(n1591), .CP(clk), .RN(n6537), 
        .Q(\registers[5][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][28]  ( .D(n1590), .CP(clk), .RN(n6544), 
        .Q(\registers[5][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][27]  ( .D(n1589), .CP(clk), .RN(n6544), 
        .Q(\registers[5][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][26]  ( .D(n1588), .CP(clk), .RN(n6544), 
        .Q(\registers[5][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][25]  ( .D(n1587), .CP(clk), .RN(n6544), 
        .Q(\registers[5][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][24]  ( .D(n1586), .CP(clk), .RN(n6538), 
        .Q(\registers[5][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][23]  ( .D(n1585), .CP(clk), .RN(n6538), 
        .Q(\registers[5][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][22]  ( .D(n1584), .CP(clk), .RN(n6538), 
        .Q(\registers[5][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][21]  ( .D(n1583), .CP(clk), .RN(n6538), 
        .Q(\registers[5][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][20]  ( .D(n1582), .CP(clk), .RN(n6598), 
        .Q(\registers[5][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][19]  ( .D(n1581), .CP(clk), .RN(n6598), 
        .Q(\registers[5][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][18]  ( .D(n1580), .CP(clk), .RN(n6597), 
        .Q(\registers[5][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][17]  ( .D(n1579), .CP(clk), .RN(n6597), 
        .Q(\registers[5][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][16]  ( .D(n1578), .CP(clk), .RN(n6543), 
        .Q(\registers[5][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][15]  ( .D(n1577), .CP(clk), .RN(n6543), 
        .Q(\registers[5][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][14]  ( .D(n1576), .CP(clk), .RN(n6543), 
        .Q(\registers[5][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][13]  ( .D(n1575), .CP(clk), .RN(n6543), 
        .Q(\registers[5][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][12]  ( .D(n1574), .CP(clk), .RN(n6537), 
        .Q(\registers[5][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][11]  ( .D(n1573), .CP(clk), .RN(n6537), 
        .Q(\registers[5][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][10]  ( .D(n1572), .CP(clk), .RN(n6537), 
        .Q(\registers[5][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][9]  ( .D(n1571), .CP(clk), .RN(n6537), .Q(
        \registers[5][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][8]  ( .D(n1570), .CP(clk), .RN(n6537), .Q(
        \registers[5][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][7]  ( .D(n1569), .CP(clk), .RN(n6537), .Q(
        \registers[5][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][6]  ( .D(n1568), .CP(clk), .RN(n6537), .Q(
        \registers[5][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][5]  ( .D(n1567), .CP(clk), .RN(n6537), .Q(
        \registers[5][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][4]  ( .D(n1566), .CP(clk), .RN(n6543), .Q(
        \registers[5][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][3]  ( .D(n1565), .CP(clk), .RN(n6543), .Q(
        \registers[5][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][2]  ( .D(n1564), .CP(clk), .RN(n6543), .Q(
        \registers[5][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][1]  ( .D(n1563), .CP(clk), .RN(n6543), .Q(
        \registers[5][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][0]  ( .D(n1562), .CP(clk), .RN(n6543), .Q(
        \registers[5][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][31]  ( .D(n1561), .CP(clk), .RN(n6547), 
        .Q(\registers[4][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][30]  ( .D(n1560), .CP(clk), .RN(n6547), 
        .Q(\registers[4][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][29]  ( .D(n1559), .CP(clk), .RN(n6547), 
        .Q(\registers[4][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][28]  ( .D(n1558), .CP(clk), .RN(n6598), 
        .Q(\registers[4][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][27]  ( .D(n1557), .CP(clk), .RN(n6547), 
        .Q(\registers[4][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][26]  ( .D(n1556), .CP(clk), .RN(n6543), 
        .Q(\registers[4][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][25]  ( .D(n1555), .CP(clk), .RN(n6543), 
        .Q(\registers[4][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][24]  ( .D(n1554), .CP(clk), .RN(n6548), 
        .Q(\registers[4][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][23]  ( .D(n1553), .CP(clk), .RN(n6548), 
        .Q(\registers[4][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][22]  ( .D(n1552), .CP(clk), .RN(n6548), 
        .Q(\registers[4][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][21]  ( .D(n1551), .CP(clk), .RN(n6548), 
        .Q(\registers[4][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][20]  ( .D(n1550), .CP(clk), .RN(n6547), 
        .Q(\registers[4][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][19]  ( .D(n1549), .CP(clk), .RN(n6547), 
        .Q(\registers[4][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][18]  ( .D(n1548), .CP(clk), .RN(n6547), 
        .Q(\registers[4][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][17]  ( .D(n1547), .CP(clk), .RN(n6547), 
        .Q(\registers[4][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][16]  ( .D(n1546), .CP(clk), .RN(n6547), 
        .Q(\registers[4][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][15]  ( .D(n1545), .CP(clk), .RN(n6547), 
        .Q(\registers[4][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][14]  ( .D(n1544), .CP(clk), .RN(n6547), 
        .Q(\registers[4][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][13]  ( .D(n1543), .CP(clk), .RN(n6547), 
        .Q(\registers[4][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][12]  ( .D(n1542), .CP(clk), .RN(n6566), 
        .Q(\registers[4][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][11]  ( .D(n1541), .CP(clk), .RN(n6548), 
        .Q(\registers[4][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][10]  ( .D(n1540), .CP(clk), .RN(n6548), 
        .Q(\registers[4][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][9]  ( .D(n1539), .CP(clk), .RN(n6548), .Q(
        \registers[4][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][8]  ( .D(n1538), .CP(clk), .RN(n6563), .Q(
        \registers[4][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][7]  ( .D(n1537), .CP(clk), .RN(n6563), .Q(
        \registers[4][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][6]  ( .D(n1536), .CP(clk), .RN(n6563), .Q(
        \registers[4][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][5]  ( .D(n1535), .CP(clk), .RN(n6563), .Q(
        \registers[4][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][4]  ( .D(n1534), .CP(clk), .RN(n6563), .Q(
        \registers[4][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][3]  ( .D(n1533), .CP(clk), .RN(n6563), .Q(
        \registers[4][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][2]  ( .D(n1532), .CP(clk), .RN(n6563), .Q(
        \registers[4][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][1]  ( .D(n1531), .CP(clk), .RN(n6563), .Q(
        \registers[4][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][0]  ( .D(n1530), .CP(clk), .RN(n6548), .Q(
        \registers[4][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][31]  ( .D(n1529), .CP(clk), .RN(n6554), 
        .Q(\registers[3][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][30]  ( .D(n1528), .CP(clk), .RN(n6554), 
        .Q(\registers[3][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][29]  ( .D(n1527), .CP(clk), .RN(n6554), 
        .Q(\registers[3][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][28]  ( .D(n1526), .CP(clk), .RN(n6554), 
        .Q(\registers[3][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][27]  ( .D(n1525), .CP(clk), .RN(n6553), 
        .Q(\registers[3][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][26]  ( .D(n1524), .CP(clk), .RN(n6553), 
        .Q(\registers[3][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][25]  ( .D(n1523), .CP(clk), .RN(n6551), 
        .Q(\registers[3][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][24]  ( .D(n1522), .CP(clk), .RN(n6550), 
        .Q(\registers[3][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][23]  ( .D(n1521), .CP(clk), .RN(n6552), 
        .Q(\registers[3][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][22]  ( .D(n1520), .CP(clk), .RN(n6552), 
        .Q(\registers[3][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][21]  ( .D(n1519), .CP(clk), .RN(n6552), 
        .Q(\registers[3][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][20]  ( .D(n1518), .CP(clk), .RN(n6576), 
        .Q(\registers[3][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][19]  ( .D(n1517), .CP(clk), .RN(n6576), 
        .Q(\registers[3][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][18]  ( .D(n1516), .CP(clk), .RN(n6576), 
        .Q(\registers[3][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][17]  ( .D(n1515), .CP(clk), .RN(n6567), 
        .Q(\registers[3][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][16]  ( .D(n1514), .CP(clk), .RN(n6578), 
        .Q(\registers[3][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][15]  ( .D(n1513), .CP(clk), .RN(n6575), 
        .Q(\registers[3][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][14]  ( .D(n1512), .CP(clk), .RN(n6575), 
        .Q(\registers[3][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][13]  ( .D(n1511), .CP(clk), .RN(n6575), 
        .Q(\registers[3][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][12]  ( .D(n1510), .CP(clk), .RN(n6575), 
        .Q(\registers[3][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][11]  ( .D(n1509), .CP(clk), .RN(n6575), 
        .Q(\registers[3][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][10]  ( .D(n1508), .CP(clk), .RN(n6575), 
        .Q(\registers[3][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][9]  ( .D(n1507), .CP(clk), .RN(n6575), .Q(
        \registers[3][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][8]  ( .D(n1506), .CP(clk), .RN(n6567), .Q(
        \registers[3][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][7]  ( .D(n1505), .CP(clk), .RN(n6565), .Q(
        \registers[3][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][6]  ( .D(n1504), .CP(clk), .RN(n6565), .Q(
        \registers[3][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][5]  ( .D(n1503), .CP(clk), .RN(n6565), .Q(
        \registers[3][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][4]  ( .D(n1502), .CP(clk), .RN(n6565), .Q(
        \registers[3][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][3]  ( .D(n1501), .CP(clk), .RN(n6565), .Q(
        \registers[3][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][2]  ( .D(n1500), .CP(clk), .RN(n6565), .Q(
        \registers[3][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][1]  ( .D(n1499), .CP(clk), .RN(n6565), .Q(
        \registers[3][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][0]  ( .D(n1498), .CP(clk), .RN(n6565), .Q(
        \registers[3][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][31]  ( .D(n1497), .CP(clk), .RN(n6575), 
        .Q(\registers[2][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][30]  ( .D(n1496), .CP(clk), .RN(n6575), 
        .Q(\registers[2][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][29]  ( .D(n1495), .CP(clk), .RN(n6575), 
        .Q(\registers[2][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][28]  ( .D(n1494), .CP(clk), .RN(n6580), 
        .Q(\registers[2][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][27]  ( .D(n1493), .CP(clk), .RN(n6580), 
        .Q(\registers[2][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][26]  ( .D(n1492), .CP(clk), .RN(n6580), 
        .Q(\registers[2][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][25]  ( .D(n1491), .CP(clk), .RN(n6580), 
        .Q(\registers[2][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][24]  ( .D(n1490), .CP(clk), .RN(n6568), 
        .Q(\registers[2][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][23]  ( .D(n1489), .CP(clk), .RN(n6566), 
        .Q(\registers[2][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][22]  ( .D(n1488), .CP(clk), .RN(n6566), 
        .Q(\registers[2][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][21]  ( .D(n1487), .CP(clk), .RN(n6566), 
        .Q(\registers[2][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][20]  ( .D(n1486), .CP(clk), .RN(n6566), 
        .Q(\registers[2][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][19]  ( .D(n1485), .CP(clk), .RN(n6566), 
        .Q(\registers[2][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][18]  ( .D(n1484), .CP(clk), .RN(n6566), 
        .Q(\registers[2][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][17]  ( .D(n1483), .CP(clk), .RN(n6579), 
        .Q(\registers[2][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][16]  ( .D(n1482), .CP(clk), .RN(n6579), 
        .Q(\registers[2][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][15]  ( .D(n1481), .CP(clk), .RN(n6578), 
        .Q(\registers[2][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][14]  ( .D(n1480), .CP(clk), .RN(n6575), 
        .Q(\registers[2][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][13]  ( .D(n1479), .CP(clk), .RN(n6579), 
        .Q(\registers[2][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][12]  ( .D(n1478), .CP(clk), .RN(n6579), 
        .Q(\registers[2][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][11]  ( .D(n1477), .CP(clk), .RN(n6579), 
        .Q(\registers[2][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][10]  ( .D(n1476), .CP(clk), .RN(n6579), 
        .Q(\registers[2][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][9]  ( .D(n1475), .CP(clk), .RN(n6579), .Q(
        \registers[2][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][8]  ( .D(n1474), .CP(clk), .RN(n6579), .Q(
        \registers[2][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][7]  ( .D(n1473), .CP(clk), .RN(n6579), .Q(
        \registers[2][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][6]  ( .D(n1472), .CP(clk), .RN(n6579), .Q(
        \registers[2][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][5]  ( .D(n1471), .CP(clk), .RN(n6567), .Q(
        \registers[2][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][4]  ( .D(n1470), .CP(clk), .RN(n6567), .Q(
        \registers[2][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][3]  ( .D(n1469), .CP(clk), .RN(n6567), .Q(
        \registers[2][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][2]  ( .D(n1468), .CP(clk), .RN(n6567), .Q(
        \registers[2][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][1]  ( .D(n1467), .CP(clk), .RN(n6567), .Q(
        \registers[2][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][0]  ( .D(n1466), .CP(clk), .RN(n6567), .Q(
        \registers[2][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][31]  ( .D(n1465), .CP(clk), .RN(n6582), 
        .Q(\registers[1][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][30]  ( .D(n1464), .CP(clk), .RN(n6582), 
        .Q(\registers[1][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][29]  ( .D(n1463), .CP(clk), .RN(n6582), 
        .Q(\registers[1][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][28]  ( .D(n1462), .CP(clk), .RN(n6582), 
        .Q(\registers[1][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][27]  ( .D(n1461), .CP(clk), .RN(n6575), 
        .Q(\registers[1][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][26]  ( .D(n1460), .CP(clk), .RN(n6576), 
        .Q(\registers[1][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][25]  ( .D(n1459), .CP(clk), .RN(n6581), 
        .Q(\registers[1][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][24]  ( .D(n1458), .CP(clk), .RN(n6581), 
        .Q(\registers[1][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][23]  ( .D(n1457), .CP(clk), .RN(n6581), 
        .Q(\registers[1][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][22]  ( .D(n1456), .CP(clk), .RN(n6581), 
        .Q(\registers[1][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][21]  ( .D(n1455), .CP(clk), .RN(n6581), 
        .Q(\registers[1][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][20]  ( .D(n1454), .CP(clk), .RN(n6581), 
        .Q(\registers[1][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][19]  ( .D(n1453), .CP(clk), .RN(n6581), 
        .Q(\registers[1][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][18]  ( .D(n1452), .CP(clk), .RN(n6581), 
        .Q(\registers[1][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][17]  ( .D(n1451), .CP(clk), .RN(n6581), 
        .Q(\registers[1][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][16]  ( .D(n1450), .CP(clk), .RN(n6581), 
        .Q(\registers[1][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][15]  ( .D(n1449), .CP(clk), .RN(n6581), 
        .Q(\registers[1][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][14]  ( .D(n1448), .CP(clk), .RN(n6581), 
        .Q(\registers[1][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][13]  ( .D(n1447), .CP(clk), .RN(n6564), 
        .Q(\registers[1][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][12]  ( .D(n1446), .CP(clk), .RN(n6564), 
        .Q(\registers[1][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][11]  ( .D(n1445), .CP(clk), .RN(n6564), 
        .Q(\registers[1][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][10]  ( .D(n1444), .CP(clk), .RN(n6564), 
        .Q(\registers[1][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][9]  ( .D(n1443), .CP(clk), .RN(n6560), .Q(
        \registers[1][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][8]  ( .D(n1442), .CP(clk), .RN(n6560), .Q(
        \registers[1][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][7]  ( .D(n1441), .CP(clk), .RN(n6560), .Q(
        \registers[1][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][6]  ( .D(n1440), .CP(clk), .RN(n6560), .Q(
        \registers[1][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][5]  ( .D(n1439), .CP(clk), .RN(n6560), .Q(
        \registers[1][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][4]  ( .D(n1438), .CP(clk), .RN(n6560), .Q(
        \registers[1][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][3]  ( .D(n1437), .CP(clk), .RN(n6560), .Q(
        \registers[1][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][2]  ( .D(n1436), .CP(clk), .RN(n6560), .Q(
        \registers[1][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][1]  ( .D(n1435), .CP(clk), .RN(n6558), .Q(
        \registers[1][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][0]  ( .D(n1434), .CP(clk), .RN(n6543), .Q(
        \registers[1][0] ) );
  HS65_LH_DFPRQNX9 \registers_reg[27][31]  ( .D(n2297), .CP(clk), .RN(n6616), 
        .QN(n65) );
  HS65_LH_DFPRQNX9 \registers_reg[27][30]  ( .D(n2296), .CP(clk), .RN(n6616), 
        .QN(n66) );
  HS65_LH_DFPRQNX9 \registers_reg[27][29]  ( .D(n2295), .CP(clk), .RN(n6616), 
        .QN(n67) );
  HS65_LH_DFPRQNX9 \registers_reg[27][28]  ( .D(n2294), .CP(clk), .RN(n6616), 
        .QN(n68) );
  HS65_LH_DFPRQNX9 \registers_reg[27][27]  ( .D(n2293), .CP(clk), .RN(n6616), 
        .QN(n69) );
  HS65_LH_DFPRQNX9 \registers_reg[27][26]  ( .D(n2292), .CP(clk), .RN(n6616), 
        .QN(n70) );
  HS65_LH_DFPRQNX9 \registers_reg[27][25]  ( .D(n2291), .CP(clk), .RN(n6616), 
        .QN(n71) );
  HS65_LH_DFPRQNX9 \registers_reg[27][24]  ( .D(n2290), .CP(clk), .RN(n6616), 
        .QN(n72) );
  HS65_LH_DFPRQNX9 \registers_reg[27][23]  ( .D(n2289), .CP(clk), .RN(n6615), 
        .QN(n73) );
  HS65_LH_DFPRQNX9 \registers_reg[27][22]  ( .D(n2288), .CP(clk), .RN(n6615), 
        .QN(n74) );
  HS65_LH_DFPRQNX9 \registers_reg[27][21]  ( .D(n2287), .CP(clk), .RN(n6615), 
        .QN(n75) );
  HS65_LH_DFPRQNX9 \registers_reg[27][20]  ( .D(n2286), .CP(clk), .RN(n6615), 
        .QN(n76) );
  HS65_LH_DFPRQNX9 \registers_reg[27][19]  ( .D(n2285), .CP(clk), .RN(n6615), 
        .QN(n77) );
  HS65_LH_DFPRQNX9 \registers_reg[27][18]  ( .D(n2284), .CP(clk), .RN(n6615), 
        .QN(n78) );
  HS65_LH_DFPRQNX9 \registers_reg[27][17]  ( .D(n2283), .CP(clk), .RN(n6615), 
        .QN(n79) );
  HS65_LH_DFPRQNX9 \registers_reg[27][16]  ( .D(n2282), .CP(clk), .RN(n6615), 
        .QN(n80) );
  HS65_LH_DFPRQNX9 \registers_reg[27][15]  ( .D(n2281), .CP(clk), .RN(n6615), 
        .QN(n81) );
  HS65_LH_DFPRQNX9 \registers_reg[27][14]  ( .D(n2280), .CP(clk), .RN(n6615), 
        .QN(n82) );
  HS65_LH_DFPRQNX9 \registers_reg[27][13]  ( .D(n2279), .CP(clk), .RN(n6615), 
        .QN(n83) );
  HS65_LH_DFPRQNX9 \registers_reg[27][12]  ( .D(n2278), .CP(clk), .RN(n6615), 
        .QN(n84) );
  HS65_LH_DFPRQNX9 \registers_reg[27][11]  ( .D(n2277), .CP(clk), .RN(n6615), 
        .QN(n85) );
  HS65_LH_DFPRQNX9 \registers_reg[27][10]  ( .D(n2276), .CP(clk), .RN(n6615), 
        .QN(n86) );
  HS65_LH_DFPRQNX9 \registers_reg[27][9]  ( .D(n2275), .CP(clk), .RN(n6614), 
        .QN(n87) );
  HS65_LH_DFPRQNX9 \registers_reg[27][8]  ( .D(n2274), .CP(clk), .RN(n6614), 
        .QN(n88) );
  HS65_LH_DFPRQNX9 \registers_reg[27][7]  ( .D(n2273), .CP(clk), .RN(n6614), 
        .QN(n89) );
  HS65_LH_DFPRQNX9 \registers_reg[27][6]  ( .D(n2272), .CP(clk), .RN(n6614), 
        .QN(n90) );
  HS65_LH_DFPRQNX9 \registers_reg[27][5]  ( .D(n2271), .CP(clk), .RN(n6614), 
        .QN(n91) );
  HS65_LH_DFPRQNX9 \registers_reg[27][4]  ( .D(n2270), .CP(clk), .RN(n6614), 
        .QN(n92) );
  HS65_LH_DFPRQNX9 \registers_reg[27][3]  ( .D(n2269), .CP(clk), .RN(n6614), 
        .QN(n93) );
  HS65_LH_DFPRQNX9 \registers_reg[27][2]  ( .D(n2268), .CP(clk), .RN(n6614), 
        .QN(n94) );
  HS65_LH_DFPRQNX9 \registers_reg[27][1]  ( .D(n2267), .CP(clk), .RN(n6614), 
        .QN(n95) );
  HS65_LH_DFPRQNX9 \registers_reg[27][0]  ( .D(n2266), .CP(clk), .RN(n6614), 
        .QN(n96) );
  HS65_LH_DFPRQNX9 \registers_reg[28][31]  ( .D(n2329), .CP(clk), .RN(n6611), 
        .QN(n33) );
  HS65_LH_DFPRQNX9 \registers_reg[28][30]  ( .D(n2328), .CP(clk), .RN(n6611), 
        .QN(n34) );
  HS65_LH_DFPRQNX9 \registers_reg[28][29]  ( .D(n2327), .CP(clk), .RN(n6611), 
        .QN(n35) );
  HS65_LH_DFPRQNX9 \registers_reg[28][28]  ( .D(n2326), .CP(clk), .RN(n6611), 
        .QN(n36) );
  HS65_LH_DFPRQNX9 \registers_reg[28][27]  ( .D(n2325), .CP(clk), .RN(n6611), 
        .QN(n37) );
  HS65_LH_DFPRQNX9 \registers_reg[28][26]  ( .D(n2324), .CP(clk), .RN(n6611), 
        .QN(n38) );
  HS65_LH_DFPRQNX9 \registers_reg[28][25]  ( .D(n2323), .CP(clk), .RN(n6611), 
        .QN(n39) );
  HS65_LH_DFPRQNX9 \registers_reg[28][24]  ( .D(n2322), .CP(clk), .RN(n6611), 
        .QN(n40) );
  HS65_LH_DFPRQNX9 \registers_reg[28][23]  ( .D(n2321), .CP(clk), .RN(n6611), 
        .QN(n41) );
  HS65_LH_DFPRQNX9 \registers_reg[28][22]  ( .D(n2320), .CP(clk), .RN(n6611), 
        .QN(n42) );
  HS65_LH_DFPRQNX9 \registers_reg[28][21]  ( .D(n2319), .CP(clk), .RN(n6611), 
        .QN(n43) );
  HS65_LH_DFPRQNX9 \registers_reg[28][20]  ( .D(n2318), .CP(clk), .RN(n6611), 
        .QN(n44) );
  HS65_LH_DFPRQNX9 \registers_reg[28][19]  ( .D(n2317), .CP(clk), .RN(n6611), 
        .QN(n45) );
  HS65_LH_DFPRQNX9 \registers_reg[28][18]  ( .D(n2316), .CP(clk), .RN(n6611), 
        .QN(n46) );
  HS65_LH_DFPRQNX9 \registers_reg[28][17]  ( .D(n2315), .CP(clk), .RN(n6610), 
        .QN(n47) );
  HS65_LH_DFPRQNX9 \registers_reg[28][16]  ( .D(n2314), .CP(clk), .RN(n6610), 
        .QN(n48) );
  HS65_LH_DFPRQNX9 \registers_reg[28][15]  ( .D(n2313), .CP(clk), .RN(n6610), 
        .QN(n49) );
  HS65_LH_DFPRQNX9 \registers_reg[28][14]  ( .D(n2312), .CP(clk), .RN(n6610), 
        .QN(n50) );
  HS65_LH_DFPRQNX9 \registers_reg[28][13]  ( .D(n2311), .CP(clk), .RN(n6610), 
        .QN(n51) );
  HS65_LH_DFPRQNX9 \registers_reg[28][12]  ( .D(n2310), .CP(clk), .RN(n6610), 
        .QN(n52) );
  HS65_LH_DFPRQNX9 \registers_reg[28][11]  ( .D(n2309), .CP(clk), .RN(n6610), 
        .QN(n53) );
  HS65_LH_DFPRQNX9 \registers_reg[28][10]  ( .D(n2308), .CP(clk), .RN(n6610), 
        .QN(n54) );
  HS65_LH_DFPRQNX9 \registers_reg[28][9]  ( .D(n2307), .CP(clk), .RN(n6610), 
        .QN(n55) );
  HS65_LH_DFPRQNX9 \registers_reg[28][8]  ( .D(n2306), .CP(clk), .RN(n6610), 
        .QN(n56) );
  HS65_LH_DFPRQNX9 \registers_reg[28][7]  ( .D(n2305), .CP(clk), .RN(n6610), 
        .QN(n57) );
  HS65_LH_DFPRQNX9 \registers_reg[28][6]  ( .D(n2304), .CP(clk), .RN(n6610), 
        .QN(n58) );
  HS65_LH_DFPRQNX9 \registers_reg[28][5]  ( .D(n2303), .CP(clk), .RN(n6610), 
        .QN(n59) );
  HS65_LH_DFPRQNX9 \registers_reg[28][4]  ( .D(n2302), .CP(clk), .RN(n6610), 
        .QN(n60) );
  HS65_LH_DFPRQNX9 \registers_reg[28][3]  ( .D(n2301), .CP(clk), .RN(n6609), 
        .QN(n61) );
  HS65_LH_DFPRQNX9 \registers_reg[28][2]  ( .D(n2300), .CP(clk), .RN(n6609), 
        .QN(n62) );
  HS65_LH_DFPRQNX9 \registers_reg[28][1]  ( .D(n2299), .CP(clk), .RN(n6609), 
        .QN(n63) );
  HS65_LH_DFPRQNX9 \registers_reg[28][0]  ( .D(n2298), .CP(clk), .RN(n6609), 
        .QN(n64) );
  HS65_LH_DFPRQNX9 \registers_reg[14][31]  ( .D(n1881), .CP(clk), .RN(n6609), 
        .QN(n161) );
  HS65_LH_DFPRQNX9 \registers_reg[14][30]  ( .D(n1880), .CP(clk), .RN(n6609), 
        .QN(n162) );
  HS65_LH_DFPRQNX9 \registers_reg[14][29]  ( .D(n1879), .CP(clk), .RN(n6609), 
        .QN(n163) );
  HS65_LH_DFPRQNX9 \registers_reg[14][28]  ( .D(n1878), .CP(clk), .RN(n6609), 
        .QN(n164) );
  HS65_LH_DFPRQNX9 \registers_reg[14][27]  ( .D(n1877), .CP(clk), .RN(n6609), 
        .QN(n165) );
  HS65_LH_DFPRQNX9 \registers_reg[14][26]  ( .D(n1876), .CP(clk), .RN(n6609), 
        .QN(n166) );
  HS65_LH_DFPRQNX9 \registers_reg[14][25]  ( .D(n1875), .CP(clk), .RN(n6609), 
        .QN(n167) );
  HS65_LH_DFPRQNX9 \registers_reg[14][24]  ( .D(n1874), .CP(clk), .RN(n6609), 
        .QN(n168) );
  HS65_LH_DFPRQNX9 \registers_reg[14][23]  ( .D(n1873), .CP(clk), .RN(n6609), 
        .QN(n169) );
  HS65_LH_DFPRQNX9 \registers_reg[14][22]  ( .D(n1872), .CP(clk), .RN(n6609), 
        .QN(n170) );
  HS65_LH_DFPRQNX9 \registers_reg[14][21]  ( .D(n1871), .CP(clk), .RN(n6608), 
        .QN(n171) );
  HS65_LH_DFPRQNX9 \registers_reg[14][20]  ( .D(n1870), .CP(clk), .RN(n6608), 
        .QN(n172) );
  HS65_LH_DFPRQNX9 \registers_reg[14][19]  ( .D(n1869), .CP(clk), .RN(n6608), 
        .QN(n173) );
  HS65_LH_DFPRQNX9 \registers_reg[14][18]  ( .D(n1868), .CP(clk), .RN(n6608), 
        .QN(n174) );
  HS65_LH_DFPRQNX9 \registers_reg[14][17]  ( .D(n1867), .CP(clk), .RN(n6608), 
        .QN(n175) );
  HS65_LH_DFPRQNX9 \registers_reg[14][16]  ( .D(n1866), .CP(clk), .RN(n6608), 
        .QN(n176) );
  HS65_LH_DFPRQNX9 \registers_reg[14][15]  ( .D(n1865), .CP(clk), .RN(n6608), 
        .QN(n177) );
  HS65_LH_DFPRQNX9 \registers_reg[14][14]  ( .D(n1864), .CP(clk), .RN(n6608), 
        .QN(n178) );
  HS65_LH_DFPRQNX9 \registers_reg[14][13]  ( .D(n1863), .CP(clk), .RN(n6608), 
        .QN(n179) );
  HS65_LH_DFPRQNX9 \registers_reg[14][12]  ( .D(n1862), .CP(clk), .RN(n6608), 
        .QN(n180) );
  HS65_LH_DFPRQNX9 \registers_reg[14][11]  ( .D(n1861), .CP(clk), .RN(n6608), 
        .QN(n181) );
  HS65_LH_DFPRQNX9 \registers_reg[14][10]  ( .D(n1860), .CP(clk), .RN(n6608), 
        .QN(n182) );
  HS65_LH_DFPRQNX9 \registers_reg[14][9]  ( .D(n1859), .CP(clk), .RN(n6608), 
        .QN(n183) );
  HS65_LH_DFPRQNX9 \registers_reg[14][8]  ( .D(n1858), .CP(clk), .RN(n6608), 
        .QN(n184) );
  HS65_LH_DFPRQNX9 \registers_reg[14][7]  ( .D(n1857), .CP(clk), .RN(n6607), 
        .QN(n185) );
  HS65_LH_DFPRQNX9 \registers_reg[14][6]  ( .D(n1856), .CP(clk), .RN(n6607), 
        .QN(n186) );
  HS65_LH_DFPRQNX9 \registers_reg[14][5]  ( .D(n1855), .CP(clk), .RN(n6607), 
        .QN(n187) );
  HS65_LH_DFPRQNX9 \registers_reg[14][4]  ( .D(n1854), .CP(clk), .RN(n6607), 
        .QN(n188) );
  HS65_LH_DFPRQNX9 \registers_reg[14][3]  ( .D(n1853), .CP(clk), .RN(n6607), 
        .QN(n189) );
  HS65_LH_DFPRQNX9 \registers_reg[14][2]  ( .D(n1852), .CP(clk), .RN(n6607), 
        .QN(n190) );
  HS65_LH_DFPRQNX9 \registers_reg[14][1]  ( .D(n1851), .CP(clk), .RN(n6607), 
        .QN(n191) );
  HS65_LH_DFPRQNX9 \registers_reg[14][0]  ( .D(n1850), .CP(clk), .RN(n6607), 
        .QN(n192) );
  HS65_LH_DFPRQNX9 \registers_reg[26][31]  ( .D(n2265), .CP(clk), .RN(n6607), 
        .QN(n97) );
  HS65_LH_DFPRQNX9 \registers_reg[26][30]  ( .D(n2264), .CP(clk), .RN(n6607), 
        .QN(n98) );
  HS65_LH_DFPRQNX9 \registers_reg[26][29]  ( .D(n2263), .CP(clk), .RN(n6607), 
        .QN(n99) );
  HS65_LH_DFPRQNX9 \registers_reg[26][28]  ( .D(n2262), .CP(clk), .RN(n6607), 
        .QN(n100) );
  HS65_LH_DFPRQNX9 \registers_reg[26][27]  ( .D(n2261), .CP(clk), .RN(n6607), 
        .QN(n101) );
  HS65_LH_DFPRQNX9 \registers_reg[26][26]  ( .D(n2260), .CP(clk), .RN(n6607), 
        .QN(n102) );
  HS65_LH_DFPRQNX9 \registers_reg[26][25]  ( .D(n2259), .CP(clk), .RN(n6606), 
        .QN(n103) );
  HS65_LH_DFPRQNX9 \registers_reg[26][24]  ( .D(n2258), .CP(clk), .RN(n6606), 
        .QN(n104) );
  HS65_LH_DFPRQNX9 \registers_reg[26][23]  ( .D(n2257), .CP(clk), .RN(n6606), 
        .QN(n105) );
  HS65_LH_DFPRQNX9 \registers_reg[26][22]  ( .D(n2256), .CP(clk), .RN(n6606), 
        .QN(n106) );
  HS65_LH_DFPRQNX9 \registers_reg[26][21]  ( .D(n2255), .CP(clk), .RN(n6606), 
        .QN(n107) );
  HS65_LH_DFPRQNX9 \registers_reg[26][20]  ( .D(n2254), .CP(clk), .RN(n6606), 
        .QN(n108) );
  HS65_LH_DFPRQNX9 \registers_reg[26][19]  ( .D(n2253), .CP(clk), .RN(n6606), 
        .QN(n109) );
  HS65_LH_DFPRQNX9 \registers_reg[26][18]  ( .D(n2252), .CP(clk), .RN(n6606), 
        .QN(n110) );
  HS65_LH_DFPRQNX9 \registers_reg[26][17]  ( .D(n2251), .CP(clk), .RN(n6606), 
        .QN(n111) );
  HS65_LH_DFPRQNX9 \registers_reg[26][16]  ( .D(n2250), .CP(clk), .RN(n6606), 
        .QN(n112) );
  HS65_LH_DFPRQNX9 \registers_reg[26][15]  ( .D(n2249), .CP(clk), .RN(n6606), 
        .QN(n113) );
  HS65_LH_DFPRQNX9 \registers_reg[26][14]  ( .D(n2248), .CP(clk), .RN(n6606), 
        .QN(n114) );
  HS65_LH_DFPRQNX9 \registers_reg[26][13]  ( .D(n2247), .CP(clk), .RN(n6606), 
        .QN(n115) );
  HS65_LH_DFPRQNX9 \registers_reg[26][12]  ( .D(n2246), .CP(clk), .RN(n6606), 
        .QN(n116) );
  HS65_LH_DFPRQNX9 \registers_reg[26][11]  ( .D(n2245), .CP(clk), .RN(n6605), 
        .QN(n117) );
  HS65_LH_DFPRQNX9 \registers_reg[26][10]  ( .D(n2244), .CP(clk), .RN(n6605), 
        .QN(n118) );
  HS65_LH_DFPRQNX9 \registers_reg[26][9]  ( .D(n2243), .CP(clk), .RN(n6605), 
        .QN(n119) );
  HS65_LH_DFPRQNX9 \registers_reg[26][8]  ( .D(n2242), .CP(clk), .RN(n6605), 
        .QN(n120) );
  HS65_LH_DFPRQNX9 \registers_reg[26][7]  ( .D(n2241), .CP(clk), .RN(n6605), 
        .QN(n121) );
  HS65_LH_DFPRQNX9 \registers_reg[26][6]  ( .D(n2240), .CP(clk), .RN(n6605), 
        .QN(n122) );
  HS65_LH_DFPRQNX9 \registers_reg[26][5]  ( .D(n2239), .CP(clk), .RN(n6605), 
        .QN(n123) );
  HS65_LH_DFPRQNX9 \registers_reg[26][4]  ( .D(n2238), .CP(clk), .RN(n6605), 
        .QN(n124) );
  HS65_LH_DFPRQNX9 \registers_reg[26][3]  ( .D(n2237), .CP(clk), .RN(n6605), 
        .QN(n125) );
  HS65_LH_DFPRQNX9 \registers_reg[26][2]  ( .D(n2236), .CP(clk), .RN(n6605), 
        .QN(n126) );
  HS65_LH_DFPRQNX9 \registers_reg[26][1]  ( .D(n2235), .CP(clk), .RN(n6605), 
        .QN(n127) );
  HS65_LH_DFPRQNX9 \registers_reg[26][0]  ( .D(n2234), .CP(clk), .RN(n6605), 
        .QN(n128) );
  HS65_LH_DFPRQNX9 \registers_reg[29][31]  ( .D(n2361), .CP(clk), .RN(n6605), 
        .QN(n1) );
  HS65_LH_DFPRQNX9 \registers_reg[29][30]  ( .D(n2360), .CP(clk), .RN(n6605), 
        .QN(n2) );
  HS65_LH_DFPRQNX9 \registers_reg[29][29]  ( .D(n2359), .CP(clk), .RN(n6604), 
        .QN(n3) );
  HS65_LH_DFPRQNX9 \registers_reg[29][28]  ( .D(n2358), .CP(clk), .RN(n6604), 
        .QN(n4) );
  HS65_LH_DFPRQNX9 \registers_reg[29][27]  ( .D(n2357), .CP(clk), .RN(n6604), 
        .QN(n5) );
  HS65_LH_DFPRQNX9 \registers_reg[29][26]  ( .D(n2356), .CP(clk), .RN(n6604), 
        .QN(n6) );
  HS65_LH_DFPRQNX9 \registers_reg[29][25]  ( .D(n2355), .CP(clk), .RN(n6604), 
        .QN(n7) );
  HS65_LH_DFPRQNX9 \registers_reg[29][24]  ( .D(n2354), .CP(clk), .RN(n6604), 
        .QN(n8) );
  HS65_LH_DFPRQNX9 \registers_reg[29][23]  ( .D(n2353), .CP(clk), .RN(n6604), 
        .QN(n9) );
  HS65_LH_DFPRQNX9 \registers_reg[29][22]  ( .D(n2352), .CP(clk), .RN(n6604), 
        .QN(n10) );
  HS65_LH_DFPRQNX9 \registers_reg[29][21]  ( .D(n2351), .CP(clk), .RN(n6604), 
        .QN(n11) );
  HS65_LH_DFPRQNX9 \registers_reg[29][20]  ( .D(n2350), .CP(clk), .RN(n6604), 
        .QN(n12) );
  HS65_LH_DFPRQNX9 \registers_reg[29][19]  ( .D(n2349), .CP(clk), .RN(n6604), 
        .QN(n13) );
  HS65_LH_DFPRQNX9 \registers_reg[29][18]  ( .D(n2348), .CP(clk), .RN(n6604), 
        .QN(n14) );
  HS65_LH_DFPRQNX9 \registers_reg[29][17]  ( .D(n2347), .CP(clk), .RN(n6604), 
        .QN(n15) );
  HS65_LH_DFPRQNX9 \registers_reg[29][16]  ( .D(n2346), .CP(clk), .RN(n6604), 
        .QN(n16) );
  HS65_LH_DFPRQNX9 \registers_reg[29][15]  ( .D(n2345), .CP(clk), .RN(n6603), 
        .QN(n17) );
  HS65_LH_DFPRQNX9 \registers_reg[29][14]  ( .D(n2344), .CP(clk), .RN(n6603), 
        .QN(n18) );
  HS65_LH_DFPRQNX9 \registers_reg[29][13]  ( .D(n2343), .CP(clk), .RN(n6603), 
        .QN(n19) );
  HS65_LH_DFPRQNX9 \registers_reg[29][12]  ( .D(n2342), .CP(clk), .RN(n6603), 
        .QN(n20) );
  HS65_LH_DFPRQNX9 \registers_reg[29][11]  ( .D(n2341), .CP(clk), .RN(n6603), 
        .QN(n21) );
  HS65_LH_DFPRQNX9 \registers_reg[29][10]  ( .D(n2340), .CP(clk), .RN(n6603), 
        .QN(n22) );
  HS65_LH_DFPRQNX9 \registers_reg[29][9]  ( .D(n2339), .CP(clk), .RN(n6603), 
        .QN(n23) );
  HS65_LH_DFPRQNX9 \registers_reg[29][8]  ( .D(n2338), .CP(clk), .RN(n6603), 
        .QN(n24) );
  HS65_LH_DFPRQNX9 \registers_reg[29][7]  ( .D(n2337), .CP(clk), .RN(n6603), 
        .QN(n25) );
  HS65_LH_DFPRQNX9 \registers_reg[29][6]  ( .D(n2336), .CP(clk), .RN(n6603), 
        .QN(n26) );
  HS65_LH_DFPRQNX9 \registers_reg[29][5]  ( .D(n2335), .CP(clk), .RN(n6603), 
        .QN(n27) );
  HS65_LH_DFPRQNX9 \registers_reg[29][4]  ( .D(n2334), .CP(clk), .RN(n6603), 
        .QN(n28) );
  HS65_LH_DFPRQNX9 \registers_reg[29][3]  ( .D(n2333), .CP(clk), .RN(n6603), 
        .QN(n29) );
  HS65_LH_DFPRQNX9 \registers_reg[29][2]  ( .D(n2332), .CP(clk), .RN(n6603), 
        .QN(n30) );
  HS65_LH_DFPRQNX9 \registers_reg[29][1]  ( .D(n2331), .CP(clk), .RN(n6602), 
        .QN(n31) );
  HS65_LH_DFPRQNX9 \registers_reg[29][0]  ( .D(n2330), .CP(clk), .RN(n6602), 
        .QN(n32) );
  HS65_LH_DFPRQNX9 \registers_reg[8][31]  ( .D(n1689), .CP(clk), .RN(n6600), 
        .QN(n225) );
  HS65_LH_DFPRQNX9 \registers_reg[8][30]  ( .D(n1688), .CP(clk), .RN(n6600), 
        .QN(n226) );
  HS65_LH_DFPRQNX9 \registers_reg[8][29]  ( .D(n1687), .CP(clk), .RN(n6600), 
        .QN(n227) );
  HS65_LH_DFPRQNX9 \registers_reg[8][28]  ( .D(n1686), .CP(clk), .RN(n6600), 
        .QN(n228) );
  HS65_LH_DFPRQNX9 \registers_reg[8][27]  ( .D(n1685), .CP(clk), .RN(n6600), 
        .QN(n229) );
  HS65_LH_DFPRQNX9 \registers_reg[8][26]  ( .D(n1684), .CP(clk), .RN(n6600), 
        .QN(n230) );
  HS65_LH_DFPRQNX9 \registers_reg[8][25]  ( .D(n1683), .CP(clk), .RN(n6600), 
        .QN(n231) );
  HS65_LH_DFPRQNX9 \registers_reg[8][24]  ( .D(n1682), .CP(clk), .RN(n6600), 
        .QN(n232) );
  HS65_LH_DFPRQNX9 \registers_reg[8][23]  ( .D(n1681), .CP(clk), .RN(n6599), 
        .QN(n233) );
  HS65_LH_DFPRQNX9 \registers_reg[8][22]  ( .D(n1680), .CP(clk), .RN(n6599), 
        .QN(n234) );
  HS65_LH_DFPRQNX9 \registers_reg[8][21]  ( .D(n1679), .CP(clk), .RN(n6599), 
        .QN(n235) );
  HS65_LH_DFPRQNX9 \registers_reg[8][20]  ( .D(n1678), .CP(clk), .RN(n6599), 
        .QN(n236) );
  HS65_LH_DFPRQNX9 \registers_reg[8][19]  ( .D(n1677), .CP(clk), .RN(n6599), 
        .QN(n237) );
  HS65_LH_DFPRQNX9 \registers_reg[8][18]  ( .D(n1676), .CP(clk), .RN(n6599), 
        .QN(n238) );
  HS65_LH_DFPRQNX9 \registers_reg[8][17]  ( .D(n1675), .CP(clk), .RN(n6599), 
        .QN(n239) );
  HS65_LH_DFPRQNX9 \registers_reg[8][16]  ( .D(n1674), .CP(clk), .RN(n6599), 
        .QN(n240) );
  HS65_LH_DFPRQNX9 \registers_reg[8][15]  ( .D(n1673), .CP(clk), .RN(n6599), 
        .QN(n241) );
  HS65_LH_DFPRQNX9 \registers_reg[8][14]  ( .D(n1672), .CP(clk), .RN(n6599), 
        .QN(n242) );
  HS65_LH_DFPRQNX9 \registers_reg[8][13]  ( .D(n1671), .CP(clk), .RN(n6599), 
        .QN(n243) );
  HS65_LH_DFPRQNX9 \registers_reg[8][12]  ( .D(n1670), .CP(clk), .RN(n6599), 
        .QN(n244) );
  HS65_LH_DFPRQNX9 \registers_reg[8][11]  ( .D(n1669), .CP(clk), .RN(n6599), 
        .QN(n245) );
  HS65_LH_DFPRQNX9 \registers_reg[8][10]  ( .D(n1668), .CP(clk), .RN(n6599), 
        .QN(n246) );
  HS65_LH_DFPRQNX9 \registers_reg[8][9]  ( .D(n1667), .CP(clk), .RN(n6598), 
        .QN(n247) );
  HS65_LH_DFPRQNX9 \registers_reg[8][8]  ( .D(n1666), .CP(clk), .RN(n6598), 
        .QN(n248) );
  HS65_LH_DFPRQNX9 \registers_reg[8][7]  ( .D(n1665), .CP(clk), .RN(n6598), 
        .QN(n249) );
  HS65_LH_DFPRQNX9 \registers_reg[8][6]  ( .D(n1664), .CP(clk), .RN(n6598), 
        .QN(n250) );
  HS65_LH_DFPRQNX9 \registers_reg[8][5]  ( .D(n1663), .CP(clk), .RN(n6598), 
        .QN(n251) );
  HS65_LH_DFPRQNX9 \registers_reg[8][4]  ( .D(n1662), .CP(clk), .RN(n6598), 
        .QN(n252) );
  HS65_LH_DFPRQNX9 \registers_reg[8][3]  ( .D(n1661), .CP(clk), .RN(n6598), 
        .QN(n253) );
  HS65_LH_DFPRQNX9 \registers_reg[8][2]  ( .D(n1660), .CP(clk), .RN(n6598), 
        .QN(n254) );
  HS65_LH_DFPRQNX9 \registers_reg[8][1]  ( .D(n1659), .CP(clk), .RN(n6598), 
        .QN(n255) );
  HS65_LH_DFPRQNX9 \registers_reg[8][0]  ( .D(n1658), .CP(clk), .RN(n6598), 
        .QN(n256) );
  HS65_LH_DFPRQNX9 \registers_reg[15][31]  ( .D(n1913), .CP(clk), .RN(n6614), 
        .QN(n129) );
  HS65_LH_DFPRQNX9 \registers_reg[15][30]  ( .D(n1912), .CP(clk), .RN(n6614), 
        .QN(n130) );
  HS65_LH_DFPRQNX9 \registers_reg[15][29]  ( .D(n1911), .CP(clk), .RN(n6614), 
        .QN(n131) );
  HS65_LH_DFPRQNX9 \registers_reg[15][28]  ( .D(n1910), .CP(clk), .RN(n6614), 
        .QN(n132) );
  HS65_LH_DFPRQNX9 \registers_reg[15][27]  ( .D(n1909), .CP(clk), .RN(n6613), 
        .QN(n133) );
  HS65_LH_DFPRQNX9 \registers_reg[15][26]  ( .D(n1908), .CP(clk), .RN(n6613), 
        .QN(n134) );
  HS65_LH_DFPRQNX9 \registers_reg[15][25]  ( .D(n1907), .CP(clk), .RN(n6613), 
        .QN(n135) );
  HS65_LH_DFPRQNX9 \registers_reg[15][24]  ( .D(n1906), .CP(clk), .RN(n6613), 
        .QN(n136) );
  HS65_LH_DFPRQNX9 \registers_reg[15][23]  ( .D(n1905), .CP(clk), .RN(n6613), 
        .QN(n137) );
  HS65_LH_DFPRQNX9 \registers_reg[15][22]  ( .D(n1904), .CP(clk), .RN(n6613), 
        .QN(n138) );
  HS65_LH_DFPRQNX9 \registers_reg[15][21]  ( .D(n1903), .CP(clk), .RN(n6613), 
        .QN(n139) );
  HS65_LH_DFPRQNX9 \registers_reg[15][20]  ( .D(n1902), .CP(clk), .RN(n6613), 
        .QN(n140) );
  HS65_LH_DFPRQNX9 \registers_reg[15][19]  ( .D(n1901), .CP(clk), .RN(n6613), 
        .QN(n141) );
  HS65_LH_DFPRQNX9 \registers_reg[15][18]  ( .D(n1900), .CP(clk), .RN(n6613), 
        .QN(n142) );
  HS65_LH_DFPRQNX9 \registers_reg[15][17]  ( .D(n1899), .CP(clk), .RN(n6613), 
        .QN(n143) );
  HS65_LH_DFPRQNX9 \registers_reg[15][16]  ( .D(n1898), .CP(clk), .RN(n6613), 
        .QN(n144) );
  HS65_LH_DFPRQNX9 \registers_reg[15][15]  ( .D(n1897), .CP(clk), .RN(n6613), 
        .QN(n145) );
  HS65_LH_DFPRQNX9 \registers_reg[15][14]  ( .D(n1896), .CP(clk), .RN(n6613), 
        .QN(n146) );
  HS65_LH_DFPRQNX9 \registers_reg[15][13]  ( .D(n1895), .CP(clk), .RN(n6612), 
        .QN(n147) );
  HS65_LH_DFPRQNX9 \registers_reg[15][12]  ( .D(n1894), .CP(clk), .RN(n6612), 
        .QN(n148) );
  HS65_LH_DFPRQNX9 \registers_reg[15][11]  ( .D(n1893), .CP(clk), .RN(n6612), 
        .QN(n149) );
  HS65_LH_DFPRQNX9 \registers_reg[15][10]  ( .D(n1892), .CP(clk), .RN(n6612), 
        .QN(n150) );
  HS65_LH_DFPRQNX9 \registers_reg[15][9]  ( .D(n1891), .CP(clk), .RN(n6612), 
        .QN(n151) );
  HS65_LH_DFPRQNX9 \registers_reg[15][8]  ( .D(n1890), .CP(clk), .RN(n6612), 
        .QN(n152) );
  HS65_LH_DFPRQNX9 \registers_reg[15][7]  ( .D(n1889), .CP(clk), .RN(n6612), 
        .QN(n153) );
  HS65_LH_DFPRQNX9 \registers_reg[15][6]  ( .D(n1888), .CP(clk), .RN(n6612), 
        .QN(n154) );
  HS65_LH_DFPRQNX9 \registers_reg[15][5]  ( .D(n1887), .CP(clk), .RN(n6612), 
        .QN(n155) );
  HS65_LH_DFPRQNX9 \registers_reg[15][4]  ( .D(n1886), .CP(clk), .RN(n6612), 
        .QN(n156) );
  HS65_LH_DFPRQNX9 \registers_reg[15][3]  ( .D(n1885), .CP(clk), .RN(n6612), 
        .QN(n157) );
  HS65_LH_DFPRQNX9 \registers_reg[15][2]  ( .D(n1884), .CP(clk), .RN(n6612), 
        .QN(n158) );
  HS65_LH_DFPRQNX9 \registers_reg[15][1]  ( .D(n1883), .CP(clk), .RN(n6612), 
        .QN(n159) );
  HS65_LH_DFPRQNX9 \registers_reg[15][0]  ( .D(n1882), .CP(clk), .RN(n6612), 
        .QN(n160) );
  HS65_LH_DFPRQNX9 \registers_reg[9][31]  ( .D(n1721), .CP(clk), .RN(n6602), 
        .QN(n193) );
  HS65_LH_DFPRQNX9 \registers_reg[9][30]  ( .D(n1720), .CP(clk), .RN(n6602), 
        .QN(n194) );
  HS65_LH_DFPRQNX9 \registers_reg[9][29]  ( .D(n1719), .CP(clk), .RN(n6602), 
        .QN(n195) );
  HS65_LH_DFPRQNX9 \registers_reg[9][28]  ( .D(n1718), .CP(clk), .RN(n6602), 
        .QN(n196) );
  HS65_LH_DFPRQNX9 \registers_reg[9][27]  ( .D(n1717), .CP(clk), .RN(n6602), 
        .QN(n197) );
  HS65_LH_DFPRQNX9 \registers_reg[9][26]  ( .D(n1716), .CP(clk), .RN(n6602), 
        .QN(n198) );
  HS65_LH_DFPRQNX9 \registers_reg[9][25]  ( .D(n1715), .CP(clk), .RN(n6602), 
        .QN(n199) );
  HS65_LH_DFPRQNX9 \registers_reg[9][24]  ( .D(n1714), .CP(clk), .RN(n6602), 
        .QN(n200) );
  HS65_LH_DFPRQNX9 \registers_reg[9][23]  ( .D(n1713), .CP(clk), .RN(n6602), 
        .QN(n201) );
  HS65_LH_DFPRQNX9 \registers_reg[9][22]  ( .D(n1712), .CP(clk), .RN(n6602), 
        .QN(n202) );
  HS65_LH_DFPRQNX9 \registers_reg[9][21]  ( .D(n1711), .CP(clk), .RN(n6602), 
        .QN(n203) );
  HS65_LH_DFPRQNX9 \registers_reg[9][20]  ( .D(n1710), .CP(clk), .RN(n6602), 
        .QN(n204) );
  HS65_LH_DFPRQNX9 \registers_reg[9][19]  ( .D(n1709), .CP(clk), .RN(n6601), 
        .QN(n205) );
  HS65_LH_DFPRQNX9 \registers_reg[9][18]  ( .D(n1708), .CP(clk), .RN(n6601), 
        .QN(n206) );
  HS65_LH_DFPRQNX9 \registers_reg[9][17]  ( .D(n1707), .CP(clk), .RN(n6601), 
        .QN(n207) );
  HS65_LH_DFPRQNX9 \registers_reg[9][16]  ( .D(n1706), .CP(clk), .RN(n6601), 
        .QN(n208) );
  HS65_LH_DFPRQNX9 \registers_reg[9][15]  ( .D(n1705), .CP(clk), .RN(n6601), 
        .QN(n209) );
  HS65_LH_DFPRQNX9 \registers_reg[9][14]  ( .D(n1704), .CP(clk), .RN(n6601), 
        .QN(n210) );
  HS65_LH_DFPRQNX9 \registers_reg[9][13]  ( .D(n1703), .CP(clk), .RN(n6601), 
        .QN(n211) );
  HS65_LH_DFPRQNX9 \registers_reg[9][12]  ( .D(n1702), .CP(clk), .RN(n6601), 
        .QN(n212) );
  HS65_LH_DFPRQNX9 \registers_reg[9][11]  ( .D(n1701), .CP(clk), .RN(n6601), 
        .QN(n213) );
  HS65_LH_DFPRQNX9 \registers_reg[9][10]  ( .D(n1700), .CP(clk), .RN(n6601), 
        .QN(n214) );
  HS65_LH_DFPRQNX9 \registers_reg[9][9]  ( .D(n1699), .CP(clk), .RN(n6601), 
        .QN(n215) );
  HS65_LH_DFPRQNX9 \registers_reg[9][8]  ( .D(n1698), .CP(clk), .RN(n6601), 
        .QN(n216) );
  HS65_LH_DFPRQNX9 \registers_reg[9][7]  ( .D(n1697), .CP(clk), .RN(n6601), 
        .QN(n217) );
  HS65_LH_DFPRQNX9 \registers_reg[9][6]  ( .D(n1696), .CP(clk), .RN(n6601), 
        .QN(n218) );
  HS65_LH_DFPRQNX9 \registers_reg[9][5]  ( .D(n1695), .CP(clk), .RN(n6600), 
        .QN(n219) );
  HS65_LH_DFPRQNX9 \registers_reg[9][4]  ( .D(n1694), .CP(clk), .RN(n6600), 
        .QN(n220) );
  HS65_LH_DFPRQNX9 \registers_reg[9][3]  ( .D(n1693), .CP(clk), .RN(n6600), 
        .QN(n221) );
  HS65_LH_DFPRQNX9 \registers_reg[9][2]  ( .D(n1692), .CP(clk), .RN(n6600), 
        .QN(n222) );
  HS65_LH_DFPRQNX9 \registers_reg[9][1]  ( .D(n1691), .CP(clk), .RN(n6600), 
        .QN(n223) );
  HS65_LH_DFPRQNX9 \registers_reg[9][0]  ( .D(n1690), .CP(clk), .RN(n6600), 
        .QN(n224) );
  HS65_LH_AND2X4 U3 ( .A(n2824), .B(n2825), .Z(n6167) );
  HS65_LH_AND2X4 U4 ( .A(n2827), .B(n2825), .Z(n6168) );
  HS65_LH_AND2X4 U5 ( .A(n2850), .B(n2829), .Z(n6169) );
  HS65_LH_AND2X4 U6 ( .A(n2850), .B(n2833), .Z(n6170) );
  HS65_LH_AND2X4 U7 ( .A(n2841), .B(n2833), .Z(n6171) );
  HS65_LH_AND2X4 U8 ( .A(n2841), .B(n2831), .Z(n6172) );
  HS65_LH_AND2X4 U9 ( .A(n2841), .B(n2829), .Z(n6173) );
  HS65_LH_AND2X4 U10 ( .A(n2841), .B(n2824), .Z(n6174) );
  HS65_LH_AND2X4 U11 ( .A(n2841), .B(n2827), .Z(n6175) );
  HS65_LH_AND2X4 U12 ( .A(n2859), .B(n2831), .Z(n6176) );
  HS65_LH_AND2X4 U13 ( .A(n2859), .B(n2833), .Z(n6177) );
  HS65_LH_AND2X4 U14 ( .A(n2859), .B(n2835), .Z(n6178) );
  HS65_LH_AND2X4 U15 ( .A(n2859), .B(n2829), .Z(n6179) );
  HS65_LH_AND2X4 U16 ( .A(n2859), .B(n2837), .Z(n6180) );
  HS65_LH_AND2X4 U17 ( .A(n2859), .B(n2824), .Z(n6181) );
  HS65_LH_AND2X4 U18 ( .A(n1323), .B(n1330), .Z(n882) );
  HS65_LH_AND2X4 U19 ( .A(n2806), .B(n2819), .Z(n1373) );
  HS65_LH_AND2X4 U20 ( .A(n1322), .B(n1327), .Z(n862) );
  HS65_LH_AND2X4 U21 ( .A(n1326), .B(n1327), .Z(n857) );
  HS65_LH_AND2X4 U22 ( .A(n1329), .B(n1327), .Z(n868) );
  HS65_LH_AND2X4 U23 ( .A(n1329), .B(n1323), .Z(n870) );
  HS65_LH_AND2X4 U24 ( .A(n1326), .B(n1323), .Z(n866) );
  HS65_LH_AND2X4 U25 ( .A(n1324), .B(n1323), .Z(n865) );
  HS65_LH_AND2X4 U26 ( .A(n2822), .B(n2806), .Z(n1381) );
  HS65_LH_AND2X4 U27 ( .A(n2810), .B(n2806), .Z(n1354) );
  HS65_LH_AND2X4 U28 ( .A(n2813), .B(n2806), .Z(n1359) );
  HS65_LH_AND2X4 U29 ( .A(n2811), .B(n2806), .Z(n1355) );
  HS65_LH_AND2X4 U30 ( .A(n2811), .B(n2808), .Z(n1353) );
  HS65_LH_AND2X4 U31 ( .A(n2805), .B(n2808), .Z(n1348) );
  HS65_LH_AND2X4 U32 ( .A(n2813), .B(n2808), .Z(n1357) );
  HS65_LH_AND2X4 U33 ( .A(n2810), .B(n2808), .Z(n1356) );
  HS65_LH_AND2X4 U34 ( .A(n1330), .B(n1325), .Z(n881) );
  HS65_LH_AND2X4 U35 ( .A(n1338), .B(n1325), .Z(n888) );
  HS65_LH_AND2X4 U36 ( .A(n1331), .B(n1325), .Z(n892) );
  HS65_LH_AND2X4 U37 ( .A(n1329), .B(n1325), .Z(n871) );
  HS65_LH_AND2X4 U38 ( .A(n1326), .B(n1325), .Z(n869) );
  HS65_LH_AND2X4 U39 ( .A(n1322), .B(n1325), .Z(n864) );
  HS65_LH_AND2X4 U40 ( .A(n2805), .B(n2812), .Z(n1352) );
  HS65_LH_AND2X4 U41 ( .A(n2813), .B(n2812), .Z(n1361) );
  HS65_LH_AND2X4 U42 ( .A(n2810), .B(n2812), .Z(n1360) );
  HS65_LH_AND2X4 U43 ( .A(n2812), .B(n2822), .Z(n1380) );
  HS65_LH_AND2X4 U44 ( .A(n2820), .B(n2807), .Z(n1367) );
  HS65_LH_AND2X4 U45 ( .A(n2813), .B(n2807), .Z(n1362) );
  HS65_LH_AND2X4 U46 ( .A(n2811), .B(n2807), .Z(n1358) );
  HS65_LH_AND2X4 U47 ( .A(n1324), .B(n1328), .Z(n886) );
  HS65_LH_AND2X4 U48 ( .A(n1329), .B(n1328), .Z(n863) );
  HS65_LH_AND2X4 U49 ( .A(n1326), .B(n1328), .Z(n856) );
  HS65_LH_AND2X4 U50 ( .A(n1327), .B(n1331), .Z(n891) );
  HS65_LH_AND2X4 U51 ( .A(n1327), .B(n1330), .Z(n861) );
  HS65_LH_AND2X4 U52 ( .A(n1323), .B(n1331), .Z(n867) );
  HS65_LH_AND2X4 U53 ( .A(n2808), .B(n2819), .Z(n1372) );
  HS65_LH_AND2X4 U54 ( .A(n2812), .B(n2809), .Z(n1379) );
  HS65_LH_AND2X4 U55 ( .A(n2812), .B(n2819), .Z(n1377) );
  HS65_LH_AND2X4 U56 ( .A(n2806), .B(n2809), .Z(n1378) );
  HS65_LH_AND2X4 U57 ( .A(n2808), .B(n2809), .Z(n1347) );
  HS65_LH_AND2X4 U58 ( .A(n1325), .B(n1337), .Z(n876) );
  HS65_LH_AND2X4 U59 ( .A(n1327), .B(n1337), .Z(n889) );
  HS65_LH_AND2X4 U60 ( .A(n1323), .B(n1337), .Z(n890) );
  HS65_LH_AND2X4 U61 ( .A(n2812), .B(n2811), .Z(n1384) );
  HS65_LH_AND2X4 U62 ( .A(n1328), .B(n1338), .Z(n877) );
  HS65_LH_AND2X4 U63 ( .A(n1323), .B(n1338), .Z(n887) );
  HS65_LH_AND2X4 U64 ( .A(n1327), .B(n1338), .Z(n893) );
  HS65_LH_AND2X4 U65 ( .A(n2808), .B(n2820), .Z(n1368) );
  HS65_LH_AND2X4 U66 ( .A(n2806), .B(n2820), .Z(n1383) );
  HS65_LH_AND2X4 U67 ( .A(n2812), .B(n2820), .Z(n1382) );
  HS65_LH_NOR3AX2 U68 ( .A(\regfile_i[WR_EN] ), .B(n795), .C(
        \regfile_i[ADRWRITE][3] ), .Z(n2841) );
  HS65_LH_NOR3AX2 U69 ( .A(\regfile_i[WR_EN] ), .B(n811), .C(
        \regfile_i[ADRWRITE][4] ), .Z(n2850) );
  HS65_LH_NOR3AX2 U70 ( .A(\regfile_i[WR_EN] ), .B(n795), .C(n811), .Z(n2825)
         );
  HS65_LH_NOR3AX2 U71 ( .A(\regfile_i[WR_EN] ), .B(\regfile_i[ADRWRITE][3] ), 
        .C(\regfile_i[ADRWRITE][4] ), .Z(n2859) );
  HS65_LH_IVX9 U72 ( .A(\regfile_i[FORWARD_B] ), .Z(n848) );
  HS65_LH_IVX9 U73 ( .A(\regfile_i[FORWARD_A] ), .Z(n847) );
  HS65_LH_BFX9 U74 ( .A(n6626), .Z(n6598) );
  HS65_LH_BFX9 U75 ( .A(n6625), .Z(n6599) );
  HS65_LH_BFX9 U76 ( .A(n6625), .Z(n6600) );
  HS65_LH_BFX9 U77 ( .A(n6624), .Z(n6601) );
  HS65_LH_BFX9 U78 ( .A(n6624), .Z(n6602) );
  HS65_LH_BFX9 U79 ( .A(n6623), .Z(n6603) );
  HS65_LH_BFX9 U80 ( .A(n6623), .Z(n6604) );
  HS65_LH_BFX9 U81 ( .A(n6622), .Z(n6605) );
  HS65_LH_BFX9 U82 ( .A(n6622), .Z(n6606) );
  HS65_LH_BFX9 U83 ( .A(n6621), .Z(n6607) );
  HS65_LH_BFX9 U84 ( .A(n6621), .Z(n6608) );
  HS65_LH_BFX9 U85 ( .A(n6620), .Z(n6609) );
  HS65_LH_BFX9 U86 ( .A(n6620), .Z(n6610) );
  HS65_LH_BFX9 U87 ( .A(n6619), .Z(n6611) );
  HS65_LH_BFX9 U88 ( .A(n6619), .Z(n6612) );
  HS65_LH_BFX9 U89 ( .A(n6618), .Z(n6613) );
  HS65_LH_BFX9 U90 ( .A(n6618), .Z(n6614) );
  HS65_LH_BFX9 U91 ( .A(n6617), .Z(n6615) );
  HS65_LH_BFX9 U92 ( .A(n6634), .Z(n6581) );
  HS65_LH_BFX9 U93 ( .A(n6637), .Z(n6575) );
  HS65_LH_BFX9 U94 ( .A(n6651), .Z(n6547) );
  HS65_LH_BFX9 U95 ( .A(n6653), .Z(n6543) );
  HS65_LH_BFX9 U96 ( .A(n6642), .Z(n6566) );
  HS65_LH_BFX9 U97 ( .A(n6641), .Z(n6567) );
  HS65_LH_BFX9 U98 ( .A(n6642), .Z(n6565) );
  HS65_LH_BFX9 U99 ( .A(n6656), .Z(n6537) );
  HS65_LH_BFX9 U100 ( .A(n6643), .Z(n6564) );
  HS65_LH_BFX9 U101 ( .A(n6643), .Z(n6563) );
  HS65_LH_BFX9 U102 ( .A(n6649), .Z(n6551) );
  HS65_LH_BFX9 U103 ( .A(n6650), .Z(n6549) );
  HS65_LH_BFX9 U104 ( .A(n6652), .Z(n6546) );
  HS65_LH_BFX9 U105 ( .A(n6652), .Z(n6545) );
  HS65_LH_BFX9 U106 ( .A(n6653), .Z(n6544) );
  HS65_LH_BFX9 U107 ( .A(n6644), .Z(n6562) );
  HS65_LH_BFX9 U108 ( .A(n6645), .Z(n6560) );
  HS65_LH_BFX9 U109 ( .A(n6644), .Z(n6561) );
  HS65_LH_BFX9 U110 ( .A(n6645), .Z(n6559) );
  HS65_LH_BFX9 U111 ( .A(n6648), .Z(n6554) );
  HS65_LH_BFX9 U112 ( .A(n6648), .Z(n6553) );
  HS65_LH_BFX9 U113 ( .A(n6646), .Z(n6558) );
  HS65_LH_BFX9 U114 ( .A(n6647), .Z(n6556) );
  HS65_LH_BFX9 U115 ( .A(n6646), .Z(n6557) );
  HS65_LH_BFX9 U116 ( .A(n6647), .Z(n6555) );
  HS65_LH_BFX9 U117 ( .A(n6649), .Z(n6552) );
  HS65_LH_BFX9 U118 ( .A(n6650), .Z(n6550) );
  HS65_LH_BFX9 U119 ( .A(n6651), .Z(n6548) );
  HS65_LH_BFX9 U120 ( .A(n6631), .Z(n6587) );
  HS65_LH_BFX9 U121 ( .A(n6636), .Z(n6577) );
  HS65_LH_BFX9 U122 ( .A(n6637), .Z(n6576) );
  HS65_LH_BFX9 U123 ( .A(n6638), .Z(n6574) );
  HS65_LH_BFX9 U124 ( .A(n6638), .Z(n6573) );
  HS65_LH_BFX9 U125 ( .A(n6655), .Z(n6540) );
  HS65_LH_BFX9 U126 ( .A(n6654), .Z(n6542) );
  HS65_LH_BFX9 U127 ( .A(n6654), .Z(n6541) );
  HS65_LH_BFX9 U128 ( .A(n6656), .Z(n6538) );
  HS65_LH_BFX9 U129 ( .A(n6626), .Z(n6597) );
  HS65_LH_BFX9 U130 ( .A(n6627), .Z(n6596) );
  HS65_LH_BFX9 U131 ( .A(n6627), .Z(n6595) );
  HS65_LH_BFX9 U132 ( .A(n6628), .Z(n6594) );
  HS65_LH_BFX9 U133 ( .A(n6628), .Z(n6593) );
  HS65_LH_BFX9 U134 ( .A(n6629), .Z(n6592) );
  HS65_LH_BFX9 U135 ( .A(n6630), .Z(n6590) );
  HS65_LH_BFX9 U136 ( .A(n6629), .Z(n6591) );
  HS65_LH_BFX9 U137 ( .A(n6631), .Z(n6588) );
  HS65_LH_BFX9 U138 ( .A(n6630), .Z(n6589) );
  HS65_LH_BFX9 U139 ( .A(n6632), .Z(n6586) );
  HS65_LH_BFX9 U140 ( .A(n6634), .Z(n6582) );
  HS65_LH_BFX9 U141 ( .A(n6632), .Z(n6585) );
  HS65_LH_BFX9 U142 ( .A(n6635), .Z(n6579) );
  HS65_LH_BFX9 U143 ( .A(n6633), .Z(n6584) );
  HS65_LH_BFX9 U144 ( .A(n6633), .Z(n6583) );
  HS65_LH_BFX9 U145 ( .A(n6635), .Z(n6580) );
  HS65_LH_BFX9 U146 ( .A(n6636), .Z(n6578) );
  HS65_LH_BFX9 U147 ( .A(n6641), .Z(n6568) );
  HS65_LH_BFX9 U148 ( .A(n6639), .Z(n6572) );
  HS65_LH_BFX9 U149 ( .A(n6640), .Z(n6570) );
  HS65_LH_BFX9 U150 ( .A(n6639), .Z(n6571) );
  HS65_LH_BFX9 U151 ( .A(n6640), .Z(n6569) );
  HS65_LH_BFX9 U152 ( .A(n6655), .Z(n6539) );
  HS65_LH_BFX9 U153 ( .A(n6617), .Z(n6616) );
  HS65_LH_IVX9 U154 ( .A(n6239), .Z(n6238) );
  HS65_LH_IVX9 U155 ( .A(n6239), .Z(n6237) );
  HS65_LH_IVX9 U156 ( .A(n6259), .Z(n6258) );
  HS65_LH_IVX9 U157 ( .A(n6259), .Z(n6257) );
  HS65_LH_IVX9 U158 ( .A(n6264), .Z(n6263) );
  HS65_LH_IVX9 U159 ( .A(n6264), .Z(n6262) );
  HS65_LH_IVX9 U160 ( .A(n6209), .Z(n6208) );
  HS65_LH_IVX9 U161 ( .A(n6209), .Z(n6207) );
  HS65_LH_IVX9 U162 ( .A(n6299), .Z(n6298) );
  HS65_LH_IVX9 U163 ( .A(n6299), .Z(n6297) );
  HS65_LH_IVX9 U164 ( .A(n6304), .Z(n6303) );
  HS65_LH_IVX9 U165 ( .A(n6304), .Z(n6302) );
  HS65_LH_IVX9 U166 ( .A(n6229), .Z(n6228) );
  HS65_LH_IVX9 U167 ( .A(n6229), .Z(n6227) );
  HS65_LH_IVX9 U168 ( .A(n6269), .Z(n6268) );
  HS65_LH_IVX9 U169 ( .A(n6269), .Z(n6267) );
  HS65_LH_BFX9 U170 ( .A(n1373), .Z(n6367) );
  HS65_LH_BFX9 U171 ( .A(n1373), .Z(n6368) );
  HS65_LH_BFX9 U172 ( .A(n882), .Z(n6460) );
  HS65_LH_BFX9 U173 ( .A(n882), .Z(n6461) );
  HS65_LH_IVX9 U174 ( .A(n6324), .Z(n6323) );
  HS65_LH_IVX9 U175 ( .A(n6324), .Z(n6322) );
  HS65_LH_IVX9 U176 ( .A(n6309), .Z(n6308) );
  HS65_LH_IVX9 U177 ( .A(n6309), .Z(n6307) );
  HS65_LH_IVX9 U178 ( .A(n6319), .Z(n6318) );
  HS65_LH_IVX9 U179 ( .A(n6319), .Z(n6317) );
  HS65_LH_IVX9 U180 ( .A(n6314), .Z(n6313) );
  HS65_LH_IVX9 U181 ( .A(n6314), .Z(n6312) );
  HS65_LH_IVX9 U182 ( .A(n6219), .Z(n6218) );
  HS65_LH_IVX9 U183 ( .A(n6219), .Z(n6217) );
  HS65_LH_IVX9 U184 ( .A(n6224), .Z(n6223) );
  HS65_LH_IVX9 U185 ( .A(n6224), .Z(n6222) );
  HS65_LH_IVX9 U186 ( .A(n6249), .Z(n6248) );
  HS65_LH_IVX9 U187 ( .A(n6249), .Z(n6247) );
  HS65_LH_IVX9 U188 ( .A(n6254), .Z(n6253) );
  HS65_LH_IVX9 U189 ( .A(n6254), .Z(n6252) );
  HS65_LH_BFX9 U190 ( .A(n6168), .Z(n6330) );
  HS65_LH_BFX9 U191 ( .A(n6167), .Z(n6335) );
  HS65_LH_BFX9 U192 ( .A(n6171), .Z(n6275) );
  HS65_LH_BFX9 U193 ( .A(n6172), .Z(n6280) );
  HS65_LH_BFX9 U194 ( .A(n6173), .Z(n6285) );
  HS65_LH_BFX9 U195 ( .A(n6175), .Z(n6290) );
  HS65_LH_BFX9 U196 ( .A(n6174), .Z(n6295) );
  HS65_LH_BFX9 U197 ( .A(n6180), .Z(n6185) );
  HS65_LH_BFX9 U198 ( .A(n6181), .Z(n6215) );
  HS65_LH_BFX9 U199 ( .A(n6170), .Z(n6235) );
  HS65_LH_BFX9 U200 ( .A(n6169), .Z(n6245) );
  HS65_LH_BFX9 U201 ( .A(n6178), .Z(n6190) );
  HS65_LH_BFX9 U202 ( .A(n6177), .Z(n6195) );
  HS65_LH_BFX9 U203 ( .A(n6176), .Z(n6200) );
  HS65_LH_BFX9 U204 ( .A(n6179), .Z(n6205) );
  HS65_LH_BFX9 U205 ( .A(n1373), .Z(n6369) );
  HS65_LH_BFX9 U206 ( .A(n882), .Z(n6462) );
  HS65_LH_IVX9 U207 ( .A(n6234), .Z(n6232) );
  HS65_LH_IVX9 U208 ( .A(n6234), .Z(n6233) );
  HS65_LH_IVX9 U209 ( .A(n6244), .Z(n6242) );
  HS65_LH_IVX9 U210 ( .A(n6244), .Z(n6243) );
  HS65_LH_IVX9 U211 ( .A(n6189), .Z(n6187) );
  HS65_LH_IVX9 U212 ( .A(n6189), .Z(n6188) );
  HS65_LH_IVX9 U213 ( .A(n6194), .Z(n6192) );
  HS65_LH_IVX9 U214 ( .A(n6194), .Z(n6193) );
  HS65_LH_IVX9 U215 ( .A(n6199), .Z(n6197) );
  HS65_LH_IVX9 U216 ( .A(n6199), .Z(n6198) );
  HS65_LH_IVX9 U217 ( .A(n6204), .Z(n6202) );
  HS65_LH_IVX9 U218 ( .A(n6204), .Z(n6203) );
  HS65_LH_IVX9 U219 ( .A(n6274), .Z(n6272) );
  HS65_LH_IVX9 U220 ( .A(n6274), .Z(n6273) );
  HS65_LH_IVX9 U221 ( .A(n6279), .Z(n6277) );
  HS65_LH_IVX9 U222 ( .A(n6279), .Z(n6278) );
  HS65_LH_IVX9 U223 ( .A(n6284), .Z(n6282) );
  HS65_LH_IVX9 U224 ( .A(n6284), .Z(n6283) );
  HS65_LH_IVX9 U225 ( .A(n6289), .Z(n6287) );
  HS65_LH_IVX9 U226 ( .A(n6289), .Z(n6288) );
  HS65_LH_IVX9 U227 ( .A(n6294), .Z(n6292) );
  HS65_LH_IVX9 U228 ( .A(n6294), .Z(n6293) );
  HS65_LH_IVX9 U229 ( .A(n6184), .Z(n6182) );
  HS65_LH_IVX9 U230 ( .A(n6184), .Z(n6183) );
  HS65_LH_IVX9 U231 ( .A(n6214), .Z(n6212) );
  HS65_LH_IVX9 U232 ( .A(n6214), .Z(n6213) );
  HS65_LH_IVX9 U233 ( .A(n6329), .Z(n6327) );
  HS65_LH_IVX9 U234 ( .A(n6329), .Z(n6328) );
  HS65_LH_IVX9 U235 ( .A(n6334), .Z(n6332) );
  HS65_LH_IVX9 U236 ( .A(n6334), .Z(n6333) );
  HS65_LH_BFX9 U237 ( .A(n6168), .Z(n6331) );
  HS65_LH_BFX9 U238 ( .A(n6167), .Z(n6336) );
  HS65_LH_BFX9 U239 ( .A(n6171), .Z(n6276) );
  HS65_LH_BFX9 U240 ( .A(n6172), .Z(n6281) );
  HS65_LH_BFX9 U241 ( .A(n6173), .Z(n6286) );
  HS65_LH_BFX9 U242 ( .A(n6175), .Z(n6291) );
  HS65_LH_BFX9 U243 ( .A(n6174), .Z(n6296) );
  HS65_LH_BFX9 U244 ( .A(n6180), .Z(n6186) );
  HS65_LH_BFX9 U245 ( .A(n6181), .Z(n6216) );
  HS65_LH_BFX9 U246 ( .A(n6170), .Z(n6236) );
  HS65_LH_BFX9 U247 ( .A(n6169), .Z(n6246) );
  HS65_LH_BFX9 U248 ( .A(n6178), .Z(n6191) );
  HS65_LH_BFX9 U249 ( .A(n6177), .Z(n6196) );
  HS65_LH_BFX9 U250 ( .A(n6176), .Z(n6201) );
  HS65_LH_BFX9 U251 ( .A(n6179), .Z(n6206) );
  HS65_LH_BFX9 U252 ( .A(n6659), .Z(n6642) );
  HS65_LH_BFX9 U253 ( .A(n6659), .Z(n6643) );
  HS65_LH_BFX9 U254 ( .A(n6657), .Z(n6652) );
  HS65_LH_BFX9 U255 ( .A(n6657), .Z(n6653) );
  HS65_LH_BFX9 U256 ( .A(n6659), .Z(n6644) );
  HS65_LH_BFX9 U257 ( .A(n6659), .Z(n6645) );
  HS65_LH_BFX9 U258 ( .A(n6658), .Z(n6648) );
  HS65_LH_BFX9 U259 ( .A(n6659), .Z(n6646) );
  HS65_LH_BFX9 U260 ( .A(n6658), .Z(n6647) );
  HS65_LH_BFX9 U261 ( .A(n6658), .Z(n6649) );
  HS65_LH_BFX9 U262 ( .A(n6658), .Z(n6650) );
  HS65_LH_BFX9 U263 ( .A(n6658), .Z(n6651) );
  HS65_LH_BFX9 U264 ( .A(n6660), .Z(n6637) );
  HS65_LH_BFX9 U265 ( .A(n6660), .Z(n6638) );
  HS65_LH_BFX9 U266 ( .A(n6657), .Z(n6654) );
  HS65_LH_BFX9 U267 ( .A(n6657), .Z(n6656) );
  HS65_LH_BFX9 U268 ( .A(n6662), .Z(n6627) );
  HS65_LH_BFX9 U269 ( .A(n6662), .Z(n6628) );
  HS65_LH_BFX9 U270 ( .A(n6662), .Z(n6629) );
  HS65_LH_BFX9 U271 ( .A(n6662), .Z(n6631) );
  HS65_LH_BFX9 U272 ( .A(n6662), .Z(n6630) );
  HS65_LH_BFX9 U273 ( .A(n6661), .Z(n6634) );
  HS65_LH_BFX9 U274 ( .A(n6661), .Z(n6632) );
  HS65_LH_BFX9 U275 ( .A(n6661), .Z(n6633) );
  HS65_LH_BFX9 U276 ( .A(n6661), .Z(n6635) );
  HS65_LH_BFX9 U277 ( .A(n6661), .Z(n6636) );
  HS65_LH_BFX9 U278 ( .A(n6660), .Z(n6641) );
  HS65_LH_BFX9 U279 ( .A(n6660), .Z(n6639) );
  HS65_LH_BFX9 U280 ( .A(n6660), .Z(n6640) );
  HS65_LH_BFX9 U281 ( .A(n6657), .Z(n6655) );
  HS65_LH_BFX9 U282 ( .A(n6663), .Z(n6625) );
  HS65_LH_BFX9 U283 ( .A(n6663), .Z(n6624) );
  HS65_LH_BFX9 U284 ( .A(n6663), .Z(n6623) );
  HS65_LH_BFX9 U285 ( .A(n6663), .Z(n6622) );
  HS65_LH_BFX9 U286 ( .A(n6664), .Z(n6621) );
  HS65_LH_BFX9 U287 ( .A(n6664), .Z(n6620) );
  HS65_LH_BFX9 U288 ( .A(n6664), .Z(n6619) );
  HS65_LH_BFX9 U289 ( .A(n6664), .Z(n6618) );
  HS65_LH_BFX9 U290 ( .A(n6664), .Z(n6617) );
  HS65_LH_BFX9 U291 ( .A(n6663), .Z(n6626) );
  HS65_LH_BFX9 U292 ( .A(n2853), .Z(n6239) );
  HS65_LH_BFX9 U293 ( .A(n2848), .Z(n6259) );
  HS65_LH_BFX9 U294 ( .A(n2847), .Z(n6264) );
  HS65_LH_BFX9 U295 ( .A(n2860), .Z(n6209) );
  HS65_LH_BFX9 U296 ( .A(n2857), .Z(n6219) );
  HS65_LH_BFX9 U297 ( .A(n2856), .Z(n6224) );
  HS65_LH_BFX9 U298 ( .A(n2851), .Z(n6249) );
  HS65_LH_BFX9 U299 ( .A(n2849), .Z(n6254) );
  HS65_LH_BFX9 U300 ( .A(n2855), .Z(n6229) );
  HS65_LH_BFX9 U301 ( .A(n2846), .Z(n6269) );
  HS65_LH_BFX9 U302 ( .A(n2828), .Z(n6324) );
  HS65_LH_BFX9 U303 ( .A(n2834), .Z(n6309) );
  HS65_LH_BFX9 U304 ( .A(n2830), .Z(n6319) );
  HS65_LH_BFX9 U305 ( .A(n2832), .Z(n6314) );
  HS65_LH_BFX9 U306 ( .A(n2838), .Z(n6299) );
  HS65_LH_BFX9 U307 ( .A(n2836), .Z(n6304) );
  HS65_LH_BFX9 U308 ( .A(n2857), .Z(n6220) );
  HS65_LH_BFX9 U309 ( .A(n2856), .Z(n6225) );
  HS65_LH_BFX9 U310 ( .A(n2851), .Z(n6250) );
  HS65_LH_BFX9 U311 ( .A(n2849), .Z(n6255) );
  HS65_LH_BFX9 U312 ( .A(n2855), .Z(n6230) );
  HS65_LH_BFX9 U313 ( .A(n2846), .Z(n6270) );
  HS65_LH_BFX9 U314 ( .A(n2828), .Z(n6325) );
  HS65_LH_BFX9 U315 ( .A(n2834), .Z(n6310) );
  HS65_LH_BFX9 U316 ( .A(n2830), .Z(n6320) );
  HS65_LH_BFX9 U317 ( .A(n2832), .Z(n6315) );
  HS65_LH_BFX9 U318 ( .A(n2838), .Z(n6300) );
  HS65_LH_BFX9 U319 ( .A(n2836), .Z(n6305) );
  HS65_LH_BFX9 U320 ( .A(n2853), .Z(n6240) );
  HS65_LH_BFX9 U321 ( .A(n2848), .Z(n6260) );
  HS65_LH_BFX9 U322 ( .A(n2847), .Z(n6265) );
  HS65_LH_BFX9 U323 ( .A(n2860), .Z(n6210) );
  HS65_LH_BFX9 U324 ( .A(n1352), .Z(n6415) );
  HS65_LH_BFX9 U325 ( .A(n1352), .Z(n6416) );
  HS65_LH_BFX9 U326 ( .A(n861), .Z(n6508) );
  HS65_LH_BFX9 U327 ( .A(n861), .Z(n6509) );
  HS65_LH_BFX9 U328 ( .A(n6168), .Z(n6329) );
  HS65_LH_BFX9 U329 ( .A(n6167), .Z(n6334) );
  HS65_LH_BFX9 U330 ( .A(n6171), .Z(n6274) );
  HS65_LH_BFX9 U331 ( .A(n6172), .Z(n6279) );
  HS65_LH_BFX9 U332 ( .A(n6173), .Z(n6284) );
  HS65_LH_BFX9 U333 ( .A(n6175), .Z(n6289) );
  HS65_LH_BFX9 U334 ( .A(n6174), .Z(n6294) );
  HS65_LH_BFX9 U335 ( .A(n6180), .Z(n6184) );
  HS65_LH_BFX9 U336 ( .A(n6181), .Z(n6214) );
  HS65_LH_BFX9 U337 ( .A(n6170), .Z(n6234) );
  HS65_LH_BFX9 U338 ( .A(n6169), .Z(n6244) );
  HS65_LH_BFX9 U339 ( .A(n6178), .Z(n6189) );
  HS65_LH_BFX9 U340 ( .A(n6177), .Z(n6194) );
  HS65_LH_BFX9 U341 ( .A(n6176), .Z(n6199) );
  HS65_LH_BFX9 U342 ( .A(n6179), .Z(n6204) );
  HS65_LH_BFX9 U343 ( .A(n1353), .Z(n6412) );
  HS65_LH_BFX9 U344 ( .A(n1353), .Z(n6413) );
  HS65_LH_BFX9 U345 ( .A(n1354), .Z(n6409) );
  HS65_LH_BFX9 U346 ( .A(n1354), .Z(n6410) );
  HS65_LH_BFX9 U347 ( .A(n862), .Z(n6505) );
  HS65_LH_BFX9 U348 ( .A(n862), .Z(n6506) );
  HS65_LH_BFX9 U349 ( .A(n863), .Z(n6502) );
  HS65_LH_BFX9 U350 ( .A(n863), .Z(n6503) );
  HS65_LH_BFX9 U351 ( .A(n881), .Z(n6463) );
  HS65_LH_BFX9 U352 ( .A(n856), .Z(n6520) );
  HS65_LH_BFX9 U353 ( .A(n881), .Z(n6464) );
  HS65_LH_BFX9 U354 ( .A(n856), .Z(n6521) );
  HS65_LH_BFX9 U355 ( .A(n1372), .Z(n6370) );
  HS65_LH_BFX9 U356 ( .A(n1367), .Z(n6382) );
  HS65_LH_BFX9 U357 ( .A(n1347), .Z(n6427) );
  HS65_LH_BFX9 U358 ( .A(n1372), .Z(n6371) );
  HS65_LH_BFX9 U359 ( .A(n1367), .Z(n6383) );
  HS65_LH_BFX9 U360 ( .A(n1347), .Z(n6428) );
  HS65_LH_BFX9 U361 ( .A(n885), .Z(n6454) );
  HS65_LH_BFX9 U362 ( .A(n885), .Z(n6455) );
  HS65_LH_BFX9 U363 ( .A(n860), .Z(n6511) );
  HS65_LH_BFX9 U364 ( .A(n860), .Z(n6512) );
  HS65_LH_BFX9 U365 ( .A(n880), .Z(n6466) );
  HS65_LH_BFX9 U366 ( .A(n880), .Z(n6467) );
  HS65_LH_BFX9 U367 ( .A(n1348), .Z(n6424) );
  HS65_LH_BFX9 U368 ( .A(n1348), .Z(n6425) );
  HS65_LH_BFX9 U369 ( .A(n1368), .Z(n6379) );
  HS65_LH_BFX9 U370 ( .A(n1368), .Z(n6380) );
  HS65_LH_BFX9 U371 ( .A(n876), .Z(n6475) );
  HS65_LH_BFX9 U372 ( .A(n876), .Z(n6476) );
  HS65_LH_BFX9 U373 ( .A(n879), .Z(n6469) );
  HS65_LH_BFX9 U374 ( .A(n879), .Z(n6470) );
  HS65_LH_BFX9 U375 ( .A(n1371), .Z(n6373) );
  HS65_LH_BFX9 U376 ( .A(n1371), .Z(n6374) );
  HS65_LH_BFX9 U377 ( .A(n877), .Z(n6472) );
  HS65_LH_BFX9 U378 ( .A(n857), .Z(n6517) );
  HS65_LH_BFX9 U379 ( .A(n877), .Z(n6473) );
  HS65_LH_BFX9 U380 ( .A(n857), .Z(n6518) );
  HS65_LH_BFX9 U381 ( .A(n1376), .Z(n6361) );
  HS65_LH_BFX9 U382 ( .A(n1351), .Z(n6418) );
  HS65_LH_BFX9 U383 ( .A(n1376), .Z(n6362) );
  HS65_LH_BFX9 U384 ( .A(n1351), .Z(n6419) );
  HS65_LH_BFX9 U385 ( .A(n859), .Z(n6514) );
  HS65_LH_BFX9 U386 ( .A(n859), .Z(n6515) );
  HS65_LH_BFX9 U387 ( .A(n884), .Z(n6457) );
  HS65_LH_BFX9 U388 ( .A(n884), .Z(n6458) );
  HS65_LH_BFX9 U389 ( .A(n2853), .Z(n6241) );
  HS65_LH_BFX9 U390 ( .A(n2848), .Z(n6261) );
  HS65_LH_BFX9 U391 ( .A(n2847), .Z(n6266) );
  HS65_LH_BFX9 U392 ( .A(n1352), .Z(n6417) );
  HS65_LH_BFX9 U393 ( .A(n861), .Z(n6510) );
  HS65_LH_BFX9 U394 ( .A(n2860), .Z(n6211) );
  HS65_LH_BFX9 U395 ( .A(n1375), .Z(n6364) );
  HS65_LH_BFX9 U396 ( .A(n1370), .Z(n6376) );
  HS65_LH_BFX9 U397 ( .A(n1350), .Z(n6421) );
  HS65_LH_BFX9 U398 ( .A(n1375), .Z(n6365) );
  HS65_LH_BFX9 U399 ( .A(n1370), .Z(n6377) );
  HS65_LH_BFX9 U400 ( .A(n1350), .Z(n6422) );
  HS65_LH_BFX9 U401 ( .A(n1353), .Z(n6414) );
  HS65_LH_BFX9 U402 ( .A(n862), .Z(n6507) );
  HS65_LH_BFX9 U403 ( .A(n2857), .Z(n6221) );
  HS65_LH_BFX9 U404 ( .A(n2856), .Z(n6226) );
  HS65_LH_BFX9 U405 ( .A(n2851), .Z(n6251) );
  HS65_LH_BFX9 U406 ( .A(n2849), .Z(n6256) );
  HS65_LH_BFX9 U407 ( .A(n2855), .Z(n6231) );
  HS65_LH_BFX9 U408 ( .A(n2846), .Z(n6271) );
  HS65_LH_BFX9 U409 ( .A(n2828), .Z(n6326) );
  HS65_LH_BFX9 U410 ( .A(n2834), .Z(n6311) );
  HS65_LH_BFX9 U411 ( .A(n2830), .Z(n6321) );
  HS65_LH_BFX9 U412 ( .A(n2832), .Z(n6316) );
  HS65_LH_BFX9 U413 ( .A(n2838), .Z(n6301) );
  HS65_LH_BFX9 U414 ( .A(n2836), .Z(n6306) );
  HS65_LH_BFX9 U415 ( .A(n863), .Z(n6504) );
  HS65_LH_BFX9 U416 ( .A(n888), .Z(n6445) );
  HS65_LH_BFX9 U417 ( .A(n866), .Z(n6493) );
  HS65_LH_BFX9 U418 ( .A(n888), .Z(n6446) );
  HS65_LH_BFX9 U419 ( .A(n866), .Z(n6494) );
  HS65_LH_BFX9 U420 ( .A(n1379), .Z(n6352) );
  HS65_LH_BFX9 U421 ( .A(n1383), .Z(n6340) );
  HS65_LH_BFX9 U422 ( .A(n1361), .Z(n6388) );
  HS65_LH_BFX9 U423 ( .A(n1357), .Z(n6400) );
  HS65_LH_BFX9 U424 ( .A(n1379), .Z(n6353) );
  HS65_LH_BFX9 U425 ( .A(n1383), .Z(n6341) );
  HS65_LH_BFX9 U426 ( .A(n1361), .Z(n6389) );
  HS65_LH_BFX9 U427 ( .A(n1357), .Z(n6401) );
  HS65_LH_BFX9 U428 ( .A(n886), .Z(n6451) );
  HS65_LH_BFX9 U429 ( .A(n886), .Z(n6452) );
  HS65_LH_BFX9 U430 ( .A(n1381), .Z(n6346) );
  HS65_LH_BFX9 U431 ( .A(n1381), .Z(n6347) );
  HS65_LH_BFX9 U432 ( .A(n1377), .Z(n6358) );
  HS65_LH_BFX9 U433 ( .A(n1359), .Z(n6394) );
  HS65_LH_BFX9 U434 ( .A(n1355), .Z(n6406) );
  HS65_LH_BFX9 U435 ( .A(n1377), .Z(n6359) );
  HS65_LH_BFX9 U436 ( .A(n1359), .Z(n6395) );
  HS65_LH_BFX9 U437 ( .A(n1355), .Z(n6407) );
  HS65_LH_BFX9 U438 ( .A(n865), .Z(n6496) );
  HS65_LH_BFX9 U439 ( .A(n865), .Z(n6497) );
  HS65_LH_BFX9 U440 ( .A(n1378), .Z(n6355) );
  HS65_LH_BFX9 U441 ( .A(n1382), .Z(n6343) );
  HS65_LH_BFX9 U442 ( .A(n1360), .Z(n6391) );
  HS65_LH_BFX9 U443 ( .A(n1356), .Z(n6403) );
  HS65_LH_BFX9 U444 ( .A(n1378), .Z(n6356) );
  HS65_LH_BFX9 U445 ( .A(n1382), .Z(n6344) );
  HS65_LH_BFX9 U446 ( .A(n1360), .Z(n6392) );
  HS65_LH_BFX9 U447 ( .A(n1356), .Z(n6404) );
  HS65_LH_BFX9 U448 ( .A(n893), .Z(n6430) );
  HS65_LH_BFX9 U449 ( .A(n893), .Z(n6431) );
  HS65_LH_BFX9 U450 ( .A(n1380), .Z(n6349) );
  HS65_LH_BFX9 U451 ( .A(n1384), .Z(n6337) );
  HS65_LH_BFX9 U452 ( .A(n1362), .Z(n6385) );
  HS65_LH_BFX9 U453 ( .A(n1358), .Z(n6397) );
  HS65_LH_BFX9 U454 ( .A(n1380), .Z(n6350) );
  HS65_LH_BFX9 U455 ( .A(n1384), .Z(n6338) );
  HS65_LH_BFX9 U456 ( .A(n1362), .Z(n6386) );
  HS65_LH_BFX9 U457 ( .A(n1358), .Z(n6398) );
  HS65_LH_BFX9 U458 ( .A(n876), .Z(n6477) );
  HS65_LH_BFX9 U459 ( .A(n889), .Z(n6442) );
  HS65_LH_BFX9 U460 ( .A(n871), .Z(n6478) );
  HS65_LH_BFX9 U461 ( .A(n867), .Z(n6490) );
  HS65_LH_BFX9 U462 ( .A(n889), .Z(n6443) );
  HS65_LH_BFX9 U463 ( .A(n871), .Z(n6479) );
  HS65_LH_BFX9 U464 ( .A(n867), .Z(n6491) );
  HS65_LH_BFX9 U465 ( .A(n887), .Z(n6448) );
  HS65_LH_BFX9 U466 ( .A(n891), .Z(n6436) );
  HS65_LH_BFX9 U467 ( .A(n869), .Z(n6484) );
  HS65_LH_BFX9 U468 ( .A(n887), .Z(n6449) );
  HS65_LH_BFX9 U469 ( .A(n891), .Z(n6437) );
  HS65_LH_BFX9 U470 ( .A(n869), .Z(n6485) );
  HS65_LH_BFX9 U471 ( .A(n879), .Z(n6471) );
  HS65_LH_BFX9 U472 ( .A(n884), .Z(n6459) );
  HS65_LH_BFX9 U473 ( .A(n859), .Z(n6516) );
  HS65_LH_BFX9 U474 ( .A(n890), .Z(n6439) );
  HS65_LH_BFX9 U475 ( .A(n868), .Z(n6487) );
  HS65_LH_BFX9 U476 ( .A(n864), .Z(n6499) );
  HS65_LH_BFX9 U477 ( .A(n890), .Z(n6440) );
  HS65_LH_BFX9 U478 ( .A(n868), .Z(n6488) );
  HS65_LH_BFX9 U479 ( .A(n864), .Z(n6500) );
  HS65_LH_BFX9 U480 ( .A(n1354), .Z(n6411) );
  HS65_LH_BFX9 U481 ( .A(n892), .Z(n6433) );
  HS65_LH_BFX9 U482 ( .A(n870), .Z(n6481) );
  HS65_LH_BFX9 U483 ( .A(n892), .Z(n6434) );
  HS65_LH_BFX9 U484 ( .A(n870), .Z(n6482) );
  HS65_LH_BFX9 U485 ( .A(n1375), .Z(n6366) );
  HS65_LH_BFX9 U486 ( .A(n1370), .Z(n6378) );
  HS65_LH_BFX9 U487 ( .A(n1350), .Z(n6423) );
  HS65_LH_BFX9 U488 ( .A(n881), .Z(n6465) );
  HS65_LH_BFX9 U489 ( .A(n856), .Z(n6522) );
  HS65_LH_BFX9 U490 ( .A(n1372), .Z(n6372) );
  HS65_LH_BFX9 U491 ( .A(n1367), .Z(n6384) );
  HS65_LH_BFX9 U492 ( .A(n1347), .Z(n6429) );
  HS65_LH_BFX9 U493 ( .A(n885), .Z(n6456) );
  HS65_LH_BFX9 U494 ( .A(n860), .Z(n6513) );
  HS65_LH_BFX9 U495 ( .A(n880), .Z(n6468) );
  HS65_LH_BFX9 U496 ( .A(n1371), .Z(n6375) );
  HS65_LH_BFX9 U497 ( .A(n1351), .Z(n6420) );
  HS65_LH_BFX9 U498 ( .A(n1376), .Z(n6363) );
  HS65_LH_BFX9 U499 ( .A(n1348), .Z(n6426) );
  HS65_LH_BFX9 U500 ( .A(n1368), .Z(n6381) );
  HS65_LH_BFX9 U501 ( .A(n877), .Z(n6474) );
  HS65_LH_BFX9 U502 ( .A(n857), .Z(n6519) );
  HS65_LH_BFX9 U503 ( .A(n865), .Z(n6498) );
  HS65_LH_BFX9 U504 ( .A(n1378), .Z(n6357) );
  HS65_LH_BFX9 U505 ( .A(n1382), .Z(n6345) );
  HS65_LH_BFX9 U506 ( .A(n1360), .Z(n6393) );
  HS65_LH_BFX9 U507 ( .A(n1356), .Z(n6405) );
  HS65_LH_BFX9 U508 ( .A(n893), .Z(n6432) );
  HS65_LH_BFX9 U509 ( .A(n1380), .Z(n6351) );
  HS65_LH_BFX9 U510 ( .A(n1384), .Z(n6339) );
  HS65_LH_BFX9 U511 ( .A(n1362), .Z(n6387) );
  HS65_LH_BFX9 U512 ( .A(n1358), .Z(n6399) );
  HS65_LH_BFX9 U513 ( .A(n889), .Z(n6444) );
  HS65_LH_BFX9 U514 ( .A(n871), .Z(n6480) );
  HS65_LH_BFX9 U515 ( .A(n867), .Z(n6492) );
  HS65_LH_BFX9 U516 ( .A(n887), .Z(n6450) );
  HS65_LH_BFX9 U517 ( .A(n891), .Z(n6438) );
  HS65_LH_BFX9 U518 ( .A(n869), .Z(n6486) );
  HS65_LH_BFX9 U519 ( .A(n890), .Z(n6441) );
  HS65_LH_BFX9 U520 ( .A(n868), .Z(n6489) );
  HS65_LH_BFX9 U521 ( .A(n864), .Z(n6501) );
  HS65_LH_BFX9 U522 ( .A(n892), .Z(n6435) );
  HS65_LH_BFX9 U523 ( .A(n870), .Z(n6483) );
  HS65_LH_BFX9 U524 ( .A(n888), .Z(n6447) );
  HS65_LH_BFX9 U525 ( .A(n866), .Z(n6495) );
  HS65_LH_BFX9 U526 ( .A(n1379), .Z(n6354) );
  HS65_LH_BFX9 U527 ( .A(n1383), .Z(n6342) );
  HS65_LH_BFX9 U528 ( .A(n1361), .Z(n6390) );
  HS65_LH_BFX9 U529 ( .A(n1357), .Z(n6402) );
  HS65_LH_BFX9 U530 ( .A(n886), .Z(n6453) );
  HS65_LH_BFX9 U531 ( .A(n1381), .Z(n6348) );
  HS65_LH_BFX9 U532 ( .A(n1377), .Z(n6360) );
  HS65_LH_BFX9 U533 ( .A(n1359), .Z(n6396) );
  HS65_LH_BFX9 U534 ( .A(n1355), .Z(n6408) );
  HS65_LH_BFX9 U535 ( .A(n6533), .Z(n6659) );
  HS65_LH_BFX9 U536 ( .A(n6533), .Z(n6658) );
  HS65_LH_BFX9 U537 ( .A(n6534), .Z(n6662) );
  HS65_LH_BFX9 U538 ( .A(n6534), .Z(n6661) );
  HS65_LH_BFX9 U539 ( .A(n6534), .Z(n6660) );
  HS65_LH_BFX9 U540 ( .A(n6533), .Z(n6657) );
  HS65_LH_BFX9 U541 ( .A(n6535), .Z(n6664) );
  HS65_LH_BFX9 U542 ( .A(n6535), .Z(n6663) );
  HS65_LH_OAI22X6 U543 ( .A(n6303), .B(n288), .C(n846), .D(n6304), .Z(n2202)
         );
  HS65_LH_OAI22X6 U544 ( .A(n6302), .B(n287), .C(n845), .D(n6305), .Z(n2203)
         );
  HS65_LH_OAI22X6 U545 ( .A(n6303), .B(n286), .C(n844), .D(n6305), .Z(n2204)
         );
  HS65_LH_OAI22X6 U546 ( .A(n6302), .B(n285), .C(n843), .D(n6305), .Z(n2205)
         );
  HS65_LH_OAI22X6 U547 ( .A(n6303), .B(n284), .C(n842), .D(n6305), .Z(n2206)
         );
  HS65_LH_OAI22X6 U548 ( .A(n6302), .B(n283), .C(n841), .D(n6305), .Z(n2207)
         );
  HS65_LH_OAI22X6 U549 ( .A(n6303), .B(n282), .C(n840), .D(n6305), .Z(n2208)
         );
  HS65_LH_OAI22X6 U550 ( .A(n6302), .B(n281), .C(n839), .D(n6305), .Z(n2209)
         );
  HS65_LH_OAI22X6 U551 ( .A(n6303), .B(n280), .C(n838), .D(n6305), .Z(n2210)
         );
  HS65_LH_OAI22X6 U552 ( .A(n6303), .B(n279), .C(n837), .D(n6305), .Z(n2211)
         );
  HS65_LH_OAI22X6 U553 ( .A(n6303), .B(n278), .C(n836), .D(n6305), .Z(n2212)
         );
  HS65_LH_OAI22X6 U554 ( .A(n6303), .B(n277), .C(n835), .D(n6305), .Z(n2213)
         );
  HS65_LH_OAI22X6 U555 ( .A(n6303), .B(n276), .C(n834), .D(n6305), .Z(n2214)
         );
  HS65_LH_OAI22X6 U556 ( .A(n6303), .B(n275), .C(n833), .D(n6305), .Z(n2215)
         );
  HS65_LH_OAI22X6 U557 ( .A(n6303), .B(n274), .C(n832), .D(n6305), .Z(n2216)
         );
  HS65_LH_OAI22X6 U558 ( .A(n6303), .B(n273), .C(n831), .D(n6305), .Z(n2217)
         );
  HS65_LH_OAI22X6 U559 ( .A(n6303), .B(n272), .C(n830), .D(n6305), .Z(n2218)
         );
  HS65_LH_OAI22X6 U560 ( .A(n6303), .B(n271), .C(n829), .D(n6305), .Z(n2219)
         );
  HS65_LH_OAI22X6 U561 ( .A(n6303), .B(n270), .C(n828), .D(n6305), .Z(n2220)
         );
  HS65_LH_OAI22X6 U562 ( .A(n6303), .B(n269), .C(n827), .D(n6305), .Z(n2221)
         );
  HS65_LH_OAI22X6 U563 ( .A(n6302), .B(n268), .C(n826), .D(n6306), .Z(n2222)
         );
  HS65_LH_OAI22X6 U564 ( .A(n6302), .B(n267), .C(n825), .D(n6306), .Z(n2223)
         );
  HS65_LH_OAI22X6 U565 ( .A(n6302), .B(n266), .C(n824), .D(n6306), .Z(n2224)
         );
  HS65_LH_OAI22X6 U566 ( .A(n6302), .B(n265), .C(n823), .D(n6306), .Z(n2225)
         );
  HS65_LH_OAI22X6 U567 ( .A(n6302), .B(n264), .C(n822), .D(n6306), .Z(n2226)
         );
  HS65_LH_OAI22X6 U568 ( .A(n6302), .B(n263), .C(n821), .D(n6306), .Z(n2227)
         );
  HS65_LH_OAI22X6 U569 ( .A(n6302), .B(n262), .C(n820), .D(n6306), .Z(n2228)
         );
  HS65_LH_OAI22X6 U570 ( .A(n6302), .B(n261), .C(n819), .D(n6306), .Z(n2229)
         );
  HS65_LH_OAI22X6 U571 ( .A(n6302), .B(n260), .C(n818), .D(n6306), .Z(n2230)
         );
  HS65_LH_OAI22X6 U572 ( .A(n6302), .B(n259), .C(n817), .D(n6306), .Z(n2231)
         );
  HS65_LH_OAI22X6 U573 ( .A(n6302), .B(n258), .C(n816), .D(n6306), .Z(n2232)
         );
  HS65_LH_OAI22X6 U574 ( .A(n6302), .B(n257), .C(n815), .D(n6306), .Z(n2233)
         );
  HS65_LH_OAI22X6 U575 ( .A(n6228), .B(n480), .C(n846), .D(n6229), .Z(n1722)
         );
  HS65_LH_OAI22X6 U576 ( .A(n6227), .B(n479), .C(n845), .D(n6230), .Z(n1723)
         );
  HS65_LH_OAI22X6 U577 ( .A(n6228), .B(n478), .C(n844), .D(n6230), .Z(n1724)
         );
  HS65_LH_OAI22X6 U578 ( .A(n6227), .B(n477), .C(n843), .D(n6230), .Z(n1725)
         );
  HS65_LH_OAI22X6 U579 ( .A(n6228), .B(n476), .C(n842), .D(n6230), .Z(n1726)
         );
  HS65_LH_OAI22X6 U580 ( .A(n6227), .B(n475), .C(n841), .D(n6230), .Z(n1727)
         );
  HS65_LH_OAI22X6 U581 ( .A(n6228), .B(n474), .C(n840), .D(n6230), .Z(n1728)
         );
  HS65_LH_OAI22X6 U582 ( .A(n6227), .B(n473), .C(n839), .D(n6230), .Z(n1729)
         );
  HS65_LH_OAI22X6 U583 ( .A(n6228), .B(n472), .C(n838), .D(n6230), .Z(n1730)
         );
  HS65_LH_OAI22X6 U584 ( .A(n6228), .B(n471), .C(n837), .D(n6230), .Z(n1731)
         );
  HS65_LH_OAI22X6 U585 ( .A(n6228), .B(n470), .C(n836), .D(n6230), .Z(n1732)
         );
  HS65_LH_OAI22X6 U586 ( .A(n6228), .B(n469), .C(n835), .D(n6230), .Z(n1733)
         );
  HS65_LH_OAI22X6 U587 ( .A(n6228), .B(n468), .C(n834), .D(n6230), .Z(n1734)
         );
  HS65_LH_OAI22X6 U588 ( .A(n6228), .B(n467), .C(n833), .D(n6230), .Z(n1735)
         );
  HS65_LH_OAI22X6 U589 ( .A(n6228), .B(n466), .C(n832), .D(n6230), .Z(n1736)
         );
  HS65_LH_OAI22X6 U590 ( .A(n6228), .B(n465), .C(n831), .D(n6230), .Z(n1737)
         );
  HS65_LH_OAI22X6 U591 ( .A(n6228), .B(n464), .C(n830), .D(n6230), .Z(n1738)
         );
  HS65_LH_OAI22X6 U592 ( .A(n6228), .B(n463), .C(n829), .D(n6230), .Z(n1739)
         );
  HS65_LH_OAI22X6 U593 ( .A(n6228), .B(n462), .C(n828), .D(n6230), .Z(n1740)
         );
  HS65_LH_OAI22X6 U594 ( .A(n6228), .B(n461), .C(n827), .D(n6230), .Z(n1741)
         );
  HS65_LH_OAI22X6 U595 ( .A(n6227), .B(n460), .C(n826), .D(n6231), .Z(n1742)
         );
  HS65_LH_OAI22X6 U596 ( .A(n6227), .B(n459), .C(n825), .D(n6231), .Z(n1743)
         );
  HS65_LH_OAI22X6 U597 ( .A(n6227), .B(n458), .C(n824), .D(n6231), .Z(n1744)
         );
  HS65_LH_OAI22X6 U598 ( .A(n6227), .B(n457), .C(n823), .D(n6231), .Z(n1745)
         );
  HS65_LH_OAI22X6 U599 ( .A(n6227), .B(n456), .C(n822), .D(n6231), .Z(n1746)
         );
  HS65_LH_OAI22X6 U600 ( .A(n6227), .B(n455), .C(n821), .D(n6231), .Z(n1747)
         );
  HS65_LH_OAI22X6 U601 ( .A(n6227), .B(n454), .C(n820), .D(n6231), .Z(n1748)
         );
  HS65_LH_OAI22X6 U602 ( .A(n6227), .B(n453), .C(n819), .D(n6231), .Z(n1749)
         );
  HS65_LH_OAI22X6 U603 ( .A(n6227), .B(n452), .C(n818), .D(n6231), .Z(n1750)
         );
  HS65_LH_OAI22X6 U604 ( .A(n6227), .B(n451), .C(n817), .D(n6231), .Z(n1751)
         );
  HS65_LH_OAI22X6 U605 ( .A(n6227), .B(n450), .C(n816), .D(n6231), .Z(n1752)
         );
  HS65_LH_OAI22X6 U606 ( .A(n6227), .B(n449), .C(n815), .D(n6231), .Z(n1753)
         );
  HS65_LH_OAI22X6 U607 ( .A(n6268), .B(n352), .C(n846), .D(n6269), .Z(n1978)
         );
  HS65_LH_OAI22X6 U608 ( .A(n6267), .B(n351), .C(n845), .D(n6270), .Z(n1979)
         );
  HS65_LH_OAI22X6 U609 ( .A(n6268), .B(n350), .C(n844), .D(n6270), .Z(n1980)
         );
  HS65_LH_OAI22X6 U610 ( .A(n6267), .B(n349), .C(n843), .D(n6270), .Z(n1981)
         );
  HS65_LH_OAI22X6 U611 ( .A(n6268), .B(n348), .C(n842), .D(n6270), .Z(n1982)
         );
  HS65_LH_OAI22X6 U612 ( .A(n6267), .B(n347), .C(n841), .D(n6270), .Z(n1983)
         );
  HS65_LH_OAI22X6 U613 ( .A(n6268), .B(n346), .C(n840), .D(n6270), .Z(n1984)
         );
  HS65_LH_OAI22X6 U614 ( .A(n6267), .B(n345), .C(n839), .D(n6270), .Z(n1985)
         );
  HS65_LH_OAI22X6 U615 ( .A(n6268), .B(n344), .C(n838), .D(n6270), .Z(n1986)
         );
  HS65_LH_OAI22X6 U616 ( .A(n6268), .B(n343), .C(n837), .D(n6270), .Z(n1987)
         );
  HS65_LH_OAI22X6 U617 ( .A(n6268), .B(n342), .C(n836), .D(n6270), .Z(n1988)
         );
  HS65_LH_OAI22X6 U618 ( .A(n6268), .B(n341), .C(n835), .D(n6270), .Z(n1989)
         );
  HS65_LH_OAI22X6 U619 ( .A(n6268), .B(n340), .C(n834), .D(n6270), .Z(n1990)
         );
  HS65_LH_OAI22X6 U620 ( .A(n6268), .B(n339), .C(n833), .D(n6270), .Z(n1991)
         );
  HS65_LH_OAI22X6 U621 ( .A(n6268), .B(n338), .C(n832), .D(n6270), .Z(n1992)
         );
  HS65_LH_OAI22X6 U622 ( .A(n6268), .B(n337), .C(n831), .D(n6270), .Z(n1993)
         );
  HS65_LH_OAI22X6 U623 ( .A(n6268), .B(n336), .C(n830), .D(n6270), .Z(n1994)
         );
  HS65_LH_OAI22X6 U624 ( .A(n6268), .B(n335), .C(n829), .D(n6270), .Z(n1995)
         );
  HS65_LH_OAI22X6 U625 ( .A(n6268), .B(n334), .C(n828), .D(n6270), .Z(n1996)
         );
  HS65_LH_OAI22X6 U626 ( .A(n6268), .B(n333), .C(n827), .D(n6270), .Z(n1997)
         );
  HS65_LH_OAI22X6 U627 ( .A(n6267), .B(n332), .C(n826), .D(n6271), .Z(n1998)
         );
  HS65_LH_OAI22X6 U628 ( .A(n6267), .B(n331), .C(n825), .D(n6271), .Z(n1999)
         );
  HS65_LH_OAI22X6 U629 ( .A(n6267), .B(n330), .C(n824), .D(n6271), .Z(n2000)
         );
  HS65_LH_OAI22X6 U630 ( .A(n6267), .B(n329), .C(n823), .D(n6271), .Z(n2001)
         );
  HS65_LH_OAI22X6 U631 ( .A(n6267), .B(n328), .C(n822), .D(n6271), .Z(n2002)
         );
  HS65_LH_OAI22X6 U632 ( .A(n6267), .B(n327), .C(n821), .D(n6271), .Z(n2003)
         );
  HS65_LH_OAI22X6 U633 ( .A(n6267), .B(n326), .C(n820), .D(n6271), .Z(n2004)
         );
  HS65_LH_OAI22X6 U634 ( .A(n6267), .B(n325), .C(n819), .D(n6271), .Z(n2005)
         );
  HS65_LH_OAI22X6 U635 ( .A(n6267), .B(n324), .C(n818), .D(n6271), .Z(n2006)
         );
  HS65_LH_OAI22X6 U636 ( .A(n6267), .B(n323), .C(n817), .D(n6271), .Z(n2007)
         );
  HS65_LH_OAI22X6 U637 ( .A(n6267), .B(n322), .C(n816), .D(n6271), .Z(n2008)
         );
  HS65_LH_OAI22X6 U638 ( .A(n6267), .B(n321), .C(n815), .D(n6271), .Z(n2009)
         );
  HS65_LH_OAI22X6 U639 ( .A(n6298), .B(n320), .C(n846), .D(n6299), .Z(n2170)
         );
  HS65_LH_OAI22X6 U640 ( .A(n6297), .B(n319), .C(n845), .D(n6300), .Z(n2171)
         );
  HS65_LH_OAI22X6 U641 ( .A(n6298), .B(n318), .C(n844), .D(n6300), .Z(n2172)
         );
  HS65_LH_OAI22X6 U642 ( .A(n6297), .B(n317), .C(n843), .D(n6300), .Z(n2173)
         );
  HS65_LH_OAI22X6 U643 ( .A(n6298), .B(n316), .C(n842), .D(n6300), .Z(n2174)
         );
  HS65_LH_OAI22X6 U644 ( .A(n6297), .B(n315), .C(n841), .D(n6300), .Z(n2175)
         );
  HS65_LH_OAI22X6 U645 ( .A(n6298), .B(n314), .C(n840), .D(n6300), .Z(n2176)
         );
  HS65_LH_OAI22X6 U646 ( .A(n6297), .B(n313), .C(n839), .D(n6300), .Z(n2177)
         );
  HS65_LH_OAI22X6 U647 ( .A(n6298), .B(n312), .C(n838), .D(n6300), .Z(n2178)
         );
  HS65_LH_OAI22X6 U648 ( .A(n6298), .B(n311), .C(n837), .D(n6300), .Z(n2179)
         );
  HS65_LH_OAI22X6 U649 ( .A(n6298), .B(n310), .C(n836), .D(n6300), .Z(n2180)
         );
  HS65_LH_OAI22X6 U650 ( .A(n6298), .B(n309), .C(n835), .D(n6300), .Z(n2181)
         );
  HS65_LH_OAI22X6 U651 ( .A(n6298), .B(n308), .C(n834), .D(n6300), .Z(n2182)
         );
  HS65_LH_OAI22X6 U652 ( .A(n6298), .B(n307), .C(n833), .D(n6300), .Z(n2183)
         );
  HS65_LH_OAI22X6 U653 ( .A(n6298), .B(n306), .C(n832), .D(n6300), .Z(n2184)
         );
  HS65_LH_OAI22X6 U654 ( .A(n6298), .B(n305), .C(n831), .D(n6300), .Z(n2185)
         );
  HS65_LH_OAI22X6 U655 ( .A(n6298), .B(n304), .C(n830), .D(n6300), .Z(n2186)
         );
  HS65_LH_OAI22X6 U656 ( .A(n6298), .B(n303), .C(n829), .D(n6300), .Z(n2187)
         );
  HS65_LH_OAI22X6 U657 ( .A(n6298), .B(n302), .C(n828), .D(n6300), .Z(n2188)
         );
  HS65_LH_OAI22X6 U658 ( .A(n6298), .B(n301), .C(n827), .D(n6300), .Z(n2189)
         );
  HS65_LH_OAI22X6 U659 ( .A(n6297), .B(n300), .C(n826), .D(n6301), .Z(n2190)
         );
  HS65_LH_OAI22X6 U660 ( .A(n6297), .B(n299), .C(n825), .D(n6301), .Z(n2191)
         );
  HS65_LH_OAI22X6 U661 ( .A(n6297), .B(n298), .C(n824), .D(n6301), .Z(n2192)
         );
  HS65_LH_OAI22X6 U662 ( .A(n6297), .B(n297), .C(n823), .D(n6301), .Z(n2193)
         );
  HS65_LH_OAI22X6 U663 ( .A(n6297), .B(n296), .C(n822), .D(n6301), .Z(n2194)
         );
  HS65_LH_OAI22X6 U664 ( .A(n6297), .B(n295), .C(n821), .D(n6301), .Z(n2195)
         );
  HS65_LH_OAI22X6 U665 ( .A(n6297), .B(n294), .C(n820), .D(n6301), .Z(n2196)
         );
  HS65_LH_OAI22X6 U666 ( .A(n6297), .B(n293), .C(n819), .D(n6301), .Z(n2197)
         );
  HS65_LH_OAI22X6 U667 ( .A(n6297), .B(n292), .C(n818), .D(n6301), .Z(n2198)
         );
  HS65_LH_OAI22X6 U668 ( .A(n6297), .B(n291), .C(n817), .D(n6301), .Z(n2199)
         );
  HS65_LH_OAI22X6 U669 ( .A(n6297), .B(n290), .C(n816), .D(n6301), .Z(n2200)
         );
  HS65_LH_OAI22X6 U670 ( .A(n6297), .B(n289), .C(n815), .D(n6301), .Z(n2201)
         );
  HS65_LH_OAI22X6 U671 ( .A(n846), .B(n6239), .C(n6238), .D(n448), .Z(n1786)
         );
  HS65_LH_OAI22X6 U672 ( .A(n846), .B(n6259), .C(n6258), .D(n416), .Z(n1914)
         );
  HS65_LH_OAI22X6 U673 ( .A(n846), .B(n6264), .C(n6263), .D(n384), .Z(n1946)
         );
  HS65_LH_OAI22X6 U674 ( .A(n846), .B(n6209), .C(n6208), .D(n512), .Z(n1594)
         );
  HS65_LH_OAI22X6 U675 ( .A(n845), .B(n6240), .C(n6237), .D(n447), .Z(n1787)
         );
  HS65_LH_OAI22X6 U676 ( .A(n844), .B(n6240), .C(n6238), .D(n446), .Z(n1788)
         );
  HS65_LH_OAI22X6 U677 ( .A(n843), .B(n6240), .C(n6237), .D(n445), .Z(n1789)
         );
  HS65_LH_OAI22X6 U678 ( .A(n842), .B(n6240), .C(n6238), .D(n444), .Z(n1790)
         );
  HS65_LH_OAI22X6 U679 ( .A(n841), .B(n6240), .C(n6237), .D(n443), .Z(n1791)
         );
  HS65_LH_OAI22X6 U680 ( .A(n840), .B(n6240), .C(n6238), .D(n442), .Z(n1792)
         );
  HS65_LH_OAI22X6 U681 ( .A(n839), .B(n6240), .C(n6238), .D(n441), .Z(n1793)
         );
  HS65_LH_OAI22X6 U682 ( .A(n838), .B(n6240), .C(n6238), .D(n440), .Z(n1794)
         );
  HS65_LH_OAI22X6 U683 ( .A(n837), .B(n6240), .C(n6238), .D(n439), .Z(n1795)
         );
  HS65_LH_OAI22X6 U684 ( .A(n836), .B(n6240), .C(n6238), .D(n438), .Z(n1796)
         );
  HS65_LH_OAI22X6 U685 ( .A(n835), .B(n6240), .C(n6238), .D(n437), .Z(n1797)
         );
  HS65_LH_OAI22X6 U686 ( .A(n834), .B(n6240), .C(n6238), .D(n436), .Z(n1798)
         );
  HS65_LH_OAI22X6 U687 ( .A(n833), .B(n6240), .C(n6238), .D(n435), .Z(n1799)
         );
  HS65_LH_OAI22X6 U688 ( .A(n832), .B(n6240), .C(n6238), .D(n434), .Z(n1800)
         );
  HS65_LH_OAI22X6 U689 ( .A(n831), .B(n6240), .C(n6238), .D(n433), .Z(n1801)
         );
  HS65_LH_OAI22X6 U690 ( .A(n830), .B(n6240), .C(n6238), .D(n432), .Z(n1802)
         );
  HS65_LH_OAI22X6 U691 ( .A(n829), .B(n6240), .C(n6238), .D(n431), .Z(n1803)
         );
  HS65_LH_OAI22X6 U692 ( .A(n828), .B(n6240), .C(n6238), .D(n430), .Z(n1804)
         );
  HS65_LH_OAI22X6 U693 ( .A(n845), .B(n6260), .C(n6257), .D(n415), .Z(n1915)
         );
  HS65_LH_OAI22X6 U694 ( .A(n844), .B(n6260), .C(n6258), .D(n414), .Z(n1916)
         );
  HS65_LH_OAI22X6 U695 ( .A(n843), .B(n6260), .C(n6257), .D(n413), .Z(n1917)
         );
  HS65_LH_OAI22X6 U696 ( .A(n842), .B(n6260), .C(n6258), .D(n412), .Z(n1918)
         );
  HS65_LH_OAI22X6 U697 ( .A(n841), .B(n6260), .C(n6257), .D(n411), .Z(n1919)
         );
  HS65_LH_OAI22X6 U698 ( .A(n840), .B(n6260), .C(n6258), .D(n410), .Z(n1920)
         );
  HS65_LH_OAI22X6 U699 ( .A(n839), .B(n6260), .C(n6258), .D(n409), .Z(n1921)
         );
  HS65_LH_OAI22X6 U700 ( .A(n838), .B(n6260), .C(n6258), .D(n408), .Z(n1922)
         );
  HS65_LH_OAI22X6 U701 ( .A(n837), .B(n6260), .C(n6258), .D(n407), .Z(n1923)
         );
  HS65_LH_OAI22X6 U702 ( .A(n836), .B(n6260), .C(n6258), .D(n406), .Z(n1924)
         );
  HS65_LH_OAI22X6 U703 ( .A(n835), .B(n6260), .C(n6258), .D(n405), .Z(n1925)
         );
  HS65_LH_OAI22X6 U704 ( .A(n834), .B(n6260), .C(n6258), .D(n404), .Z(n1926)
         );
  HS65_LH_OAI22X6 U705 ( .A(n833), .B(n6260), .C(n6258), .D(n403), .Z(n1927)
         );
  HS65_LH_OAI22X6 U706 ( .A(n832), .B(n6260), .C(n6258), .D(n402), .Z(n1928)
         );
  HS65_LH_OAI22X6 U707 ( .A(n831), .B(n6260), .C(n6258), .D(n401), .Z(n1929)
         );
  HS65_LH_OAI22X6 U708 ( .A(n830), .B(n6260), .C(n6258), .D(n400), .Z(n1930)
         );
  HS65_LH_OAI22X6 U709 ( .A(n829), .B(n6260), .C(n6258), .D(n399), .Z(n1931)
         );
  HS65_LH_OAI22X6 U710 ( .A(n828), .B(n6260), .C(n6258), .D(n398), .Z(n1932)
         );
  HS65_LH_OAI22X6 U711 ( .A(n845), .B(n6265), .C(n6262), .D(n383), .Z(n1947)
         );
  HS65_LH_OAI22X6 U712 ( .A(n844), .B(n6265), .C(n6263), .D(n382), .Z(n1948)
         );
  HS65_LH_OAI22X6 U713 ( .A(n843), .B(n6265), .C(n6262), .D(n381), .Z(n1949)
         );
  HS65_LH_OAI22X6 U714 ( .A(n842), .B(n6265), .C(n6263), .D(n380), .Z(n1950)
         );
  HS65_LH_OAI22X6 U715 ( .A(n841), .B(n6265), .C(n6262), .D(n379), .Z(n1951)
         );
  HS65_LH_OAI22X6 U716 ( .A(n840), .B(n6265), .C(n6263), .D(n378), .Z(n1952)
         );
  HS65_LH_OAI22X6 U717 ( .A(n839), .B(n6265), .C(n6263), .D(n377), .Z(n1953)
         );
  HS65_LH_OAI22X6 U718 ( .A(n838), .B(n6265), .C(n6263), .D(n376), .Z(n1954)
         );
  HS65_LH_OAI22X6 U719 ( .A(n837), .B(n6265), .C(n6263), .D(n375), .Z(n1955)
         );
  HS65_LH_OAI22X6 U720 ( .A(n836), .B(n6265), .C(n6263), .D(n374), .Z(n1956)
         );
  HS65_LH_OAI22X6 U721 ( .A(n835), .B(n6265), .C(n6263), .D(n373), .Z(n1957)
         );
  HS65_LH_OAI22X6 U722 ( .A(n834), .B(n6265), .C(n6263), .D(n372), .Z(n1958)
         );
  HS65_LH_OAI22X6 U723 ( .A(n833), .B(n6265), .C(n6263), .D(n371), .Z(n1959)
         );
  HS65_LH_OAI22X6 U724 ( .A(n832), .B(n6265), .C(n6263), .D(n370), .Z(n1960)
         );
  HS65_LH_OAI22X6 U725 ( .A(n831), .B(n6265), .C(n6263), .D(n369), .Z(n1961)
         );
  HS65_LH_OAI22X6 U726 ( .A(n830), .B(n6265), .C(n6263), .D(n368), .Z(n1962)
         );
  HS65_LH_OAI22X6 U727 ( .A(n829), .B(n6265), .C(n6263), .D(n367), .Z(n1963)
         );
  HS65_LH_OAI22X6 U728 ( .A(n828), .B(n6265), .C(n6263), .D(n366), .Z(n1964)
         );
  HS65_LH_OAI22X6 U729 ( .A(n845), .B(n6210), .C(n6207), .D(n511), .Z(n1595)
         );
  HS65_LH_OAI22X6 U730 ( .A(n844), .B(n6210), .C(n6208), .D(n510), .Z(n1596)
         );
  HS65_LH_OAI22X6 U731 ( .A(n843), .B(n6210), .C(n6207), .D(n509), .Z(n1597)
         );
  HS65_LH_OAI22X6 U732 ( .A(n842), .B(n6210), .C(n6208), .D(n508), .Z(n1598)
         );
  HS65_LH_OAI22X6 U733 ( .A(n841), .B(n6210), .C(n6207), .D(n507), .Z(n1599)
         );
  HS65_LH_OAI22X6 U734 ( .A(n840), .B(n6210), .C(n6208), .D(n506), .Z(n1600)
         );
  HS65_LH_OAI22X6 U735 ( .A(n839), .B(n6210), .C(n6208), .D(n505), .Z(n1601)
         );
  HS65_LH_OAI22X6 U736 ( .A(n838), .B(n6210), .C(n6208), .D(n504), .Z(n1602)
         );
  HS65_LH_OAI22X6 U737 ( .A(n837), .B(n6210), .C(n6208), .D(n503), .Z(n1603)
         );
  HS65_LH_OAI22X6 U738 ( .A(n836), .B(n6210), .C(n6208), .D(n502), .Z(n1604)
         );
  HS65_LH_OAI22X6 U739 ( .A(n835), .B(n6210), .C(n6208), .D(n501), .Z(n1605)
         );
  HS65_LH_OAI22X6 U740 ( .A(n834), .B(n6210), .C(n6208), .D(n500), .Z(n1606)
         );
  HS65_LH_OAI22X6 U741 ( .A(n833), .B(n6210), .C(n6208), .D(n499), .Z(n1607)
         );
  HS65_LH_OAI22X6 U742 ( .A(n832), .B(n6210), .C(n6208), .D(n498), .Z(n1608)
         );
  HS65_LH_OAI22X6 U743 ( .A(n831), .B(n6210), .C(n6208), .D(n497), .Z(n1609)
         );
  HS65_LH_OAI22X6 U744 ( .A(n830), .B(n6210), .C(n6208), .D(n496), .Z(n1610)
         );
  HS65_LH_OAI22X6 U745 ( .A(n829), .B(n6210), .C(n6208), .D(n495), .Z(n1611)
         );
  HS65_LH_OAI22X6 U746 ( .A(n828), .B(n6210), .C(n6208), .D(n494), .Z(n1612)
         );
  HS65_LH_OAI22X6 U747 ( .A(n827), .B(n6241), .C(n6237), .D(n429), .Z(n1805)
         );
  HS65_LH_OAI22X6 U748 ( .A(n826), .B(n6241), .C(n6237), .D(n428), .Z(n1806)
         );
  HS65_LH_OAI22X6 U749 ( .A(n825), .B(n6241), .C(n6237), .D(n427), .Z(n1807)
         );
  HS65_LH_OAI22X6 U750 ( .A(n824), .B(n6241), .C(n6237), .D(n426), .Z(n1808)
         );
  HS65_LH_OAI22X6 U751 ( .A(n823), .B(n6241), .C(n6237), .D(n425), .Z(n1809)
         );
  HS65_LH_OAI22X6 U752 ( .A(n822), .B(n6241), .C(n6237), .D(n424), .Z(n1810)
         );
  HS65_LH_OAI22X6 U753 ( .A(n821), .B(n6241), .C(n6237), .D(n423), .Z(n1811)
         );
  HS65_LH_OAI22X6 U754 ( .A(n820), .B(n6241), .C(n6237), .D(n422), .Z(n1812)
         );
  HS65_LH_OAI22X6 U755 ( .A(n819), .B(n6241), .C(n6237), .D(n421), .Z(n1813)
         );
  HS65_LH_OAI22X6 U756 ( .A(n818), .B(n6241), .C(n6237), .D(n420), .Z(n1814)
         );
  HS65_LH_OAI22X6 U757 ( .A(n817), .B(n6241), .C(n6237), .D(n419), .Z(n1815)
         );
  HS65_LH_OAI22X6 U758 ( .A(n816), .B(n6241), .C(n6237), .D(n418), .Z(n1816)
         );
  HS65_LH_OAI22X6 U759 ( .A(n815), .B(n6241), .C(n6237), .D(n417), .Z(n1817)
         );
  HS65_LH_OAI22X6 U760 ( .A(n827), .B(n6261), .C(n6257), .D(n397), .Z(n1933)
         );
  HS65_LH_OAI22X6 U761 ( .A(n826), .B(n6261), .C(n6257), .D(n396), .Z(n1934)
         );
  HS65_LH_OAI22X6 U762 ( .A(n825), .B(n6261), .C(n6257), .D(n395), .Z(n1935)
         );
  HS65_LH_OAI22X6 U763 ( .A(n824), .B(n6261), .C(n6257), .D(n394), .Z(n1936)
         );
  HS65_LH_OAI22X6 U764 ( .A(n823), .B(n6261), .C(n6257), .D(n393), .Z(n1937)
         );
  HS65_LH_OAI22X6 U765 ( .A(n822), .B(n6261), .C(n6257), .D(n392), .Z(n1938)
         );
  HS65_LH_OAI22X6 U766 ( .A(n821), .B(n6261), .C(n6257), .D(n391), .Z(n1939)
         );
  HS65_LH_OAI22X6 U767 ( .A(n820), .B(n6261), .C(n6257), .D(n390), .Z(n1940)
         );
  HS65_LH_OAI22X6 U768 ( .A(n819), .B(n6261), .C(n6257), .D(n389), .Z(n1941)
         );
  HS65_LH_OAI22X6 U769 ( .A(n818), .B(n6261), .C(n6257), .D(n388), .Z(n1942)
         );
  HS65_LH_OAI22X6 U770 ( .A(n817), .B(n6261), .C(n6257), .D(n387), .Z(n1943)
         );
  HS65_LH_OAI22X6 U771 ( .A(n816), .B(n6261), .C(n6257), .D(n386), .Z(n1944)
         );
  HS65_LH_OAI22X6 U772 ( .A(n815), .B(n6261), .C(n6257), .D(n385), .Z(n1945)
         );
  HS65_LH_OAI22X6 U773 ( .A(n827), .B(n6266), .C(n6262), .D(n365), .Z(n1965)
         );
  HS65_LH_OAI22X6 U774 ( .A(n826), .B(n6266), .C(n6262), .D(n364), .Z(n1966)
         );
  HS65_LH_OAI22X6 U775 ( .A(n825), .B(n6266), .C(n6262), .D(n363), .Z(n1967)
         );
  HS65_LH_OAI22X6 U776 ( .A(n824), .B(n6266), .C(n6262), .D(n362), .Z(n1968)
         );
  HS65_LH_OAI22X6 U777 ( .A(n823), .B(n6266), .C(n6262), .D(n361), .Z(n1969)
         );
  HS65_LH_OAI22X6 U778 ( .A(n822), .B(n6266), .C(n6262), .D(n360), .Z(n1970)
         );
  HS65_LH_OAI22X6 U779 ( .A(n821), .B(n6266), .C(n6262), .D(n359), .Z(n1971)
         );
  HS65_LH_OAI22X6 U780 ( .A(n820), .B(n6266), .C(n6262), .D(n358), .Z(n1972)
         );
  HS65_LH_OAI22X6 U781 ( .A(n819), .B(n6266), .C(n6262), .D(n357), .Z(n1973)
         );
  HS65_LH_OAI22X6 U782 ( .A(n818), .B(n6266), .C(n6262), .D(n356), .Z(n1974)
         );
  HS65_LH_OAI22X6 U783 ( .A(n817), .B(n6266), .C(n6262), .D(n355), .Z(n1975)
         );
  HS65_LH_OAI22X6 U784 ( .A(n816), .B(n6266), .C(n6262), .D(n354), .Z(n1976)
         );
  HS65_LH_OAI22X6 U785 ( .A(n815), .B(n6266), .C(n6262), .D(n353), .Z(n1977)
         );
  HS65_LH_OAI22X6 U786 ( .A(n827), .B(n6211), .C(n6207), .D(n493), .Z(n1613)
         );
  HS65_LH_OAI22X6 U787 ( .A(n826), .B(n6211), .C(n6207), .D(n492), .Z(n1614)
         );
  HS65_LH_OAI22X6 U788 ( .A(n825), .B(n6211), .C(n6207), .D(n491), .Z(n1615)
         );
  HS65_LH_OAI22X6 U789 ( .A(n824), .B(n6211), .C(n6207), .D(n490), .Z(n1616)
         );
  HS65_LH_OAI22X6 U790 ( .A(n823), .B(n6211), .C(n6207), .D(n489), .Z(n1617)
         );
  HS65_LH_OAI22X6 U791 ( .A(n822), .B(n6211), .C(n6207), .D(n488), .Z(n1618)
         );
  HS65_LH_OAI22X6 U792 ( .A(n821), .B(n6211), .C(n6207), .D(n487), .Z(n1619)
         );
  HS65_LH_OAI22X6 U793 ( .A(n820), .B(n6211), .C(n6207), .D(n486), .Z(n1620)
         );
  HS65_LH_OAI22X6 U794 ( .A(n819), .B(n6211), .C(n6207), .D(n485), .Z(n1621)
         );
  HS65_LH_OAI22X6 U795 ( .A(n818), .B(n6211), .C(n6207), .D(n484), .Z(n1622)
         );
  HS65_LH_OAI22X6 U796 ( .A(n817), .B(n6211), .C(n6207), .D(n483), .Z(n1623)
         );
  HS65_LH_OAI22X6 U797 ( .A(n816), .B(n6211), .C(n6207), .D(n482), .Z(n1624)
         );
  HS65_LH_OAI22X6 U798 ( .A(n815), .B(n6211), .C(n6207), .D(n481), .Z(n1625)
         );
  HS65_LH_NAND2X7 U799 ( .A(n1327), .B(n1324), .Z(n885) );
  HS65_LH_NAND2X7 U800 ( .A(n1328), .B(n1337), .Z(n879) );
  HS65_LH_NAND2X7 U801 ( .A(n2822), .B(n2807), .Z(n1375) );
  HS65_LH_NAND2X7 U802 ( .A(n2809), .B(n2807), .Z(n1371) );
  HS65_LH_NAND2X7 U803 ( .A(n2819), .B(n2807), .Z(n1370) );
  HS65_LH_NAND2X7 U804 ( .A(n2805), .B(n2807), .Z(n1350) );
  HS65_LH_NAND2X7 U805 ( .A(n1322), .B(n1323), .Z(n860) );
  HS65_LH_NAND2X7 U806 ( .A(n2805), .B(n2806), .Z(n1351) );
  HS65_LH_NAND2X7 U807 ( .A(n2822), .B(n2808), .Z(n1376) );
  HS65_LH_NAND2X7 U808 ( .A(n1330), .B(n1328), .Z(n884) );
  HS65_LH_NAND2X7 U809 ( .A(n1331), .B(n1328), .Z(n880) );
  HS65_LH_NAND2X7 U810 ( .A(n1324), .B(n1325), .Z(n859) );
  HS65_LH_NAND2X7 U811 ( .A(n2829), .B(n2825), .Z(n2828) );
  HS65_LH_NAND2X7 U812 ( .A(n2835), .B(n2825), .Z(n2834) );
  HS65_LH_NAND2X7 U813 ( .A(n2831), .B(n2825), .Z(n2830) );
  HS65_LH_NAND2X7 U814 ( .A(n2833), .B(n2825), .Z(n2832) );
  HS65_LH_NAND2X7 U815 ( .A(n2839), .B(n2825), .Z(n2838) );
  HS65_LH_NAND2X7 U816 ( .A(n2837), .B(n2825), .Z(n2836) );
  HS65_LH_NAND2X7 U817 ( .A(n2841), .B(n2839), .Z(n2848) );
  HS65_LH_NAND2X7 U818 ( .A(n2841), .B(n2837), .Z(n2847) );
  HS65_LH_NAND2X7 U819 ( .A(n2841), .B(n2835), .Z(n2846) );
  HS65_LH_NAND2X7 U820 ( .A(n2850), .B(n2839), .Z(n2857) );
  HS65_LH_NAND2X7 U821 ( .A(n2850), .B(n2837), .Z(n2856) );
  HS65_LH_NAND2X7 U822 ( .A(n2850), .B(n2827), .Z(n2851) );
  HS65_LH_NAND2X7 U823 ( .A(n2850), .B(n2824), .Z(n2849) );
  HS65_LH_NAND2X7 U824 ( .A(n2850), .B(n2835), .Z(n2855) );
  HS65_LH_NAND2X7 U825 ( .A(n2850), .B(n2831), .Z(n2853) );
  HS65_LH_NOR3X4 U826 ( .A(n813), .B(n814), .C(n812), .Z(n2824) );
  HS65_LH_NAND2X7 U827 ( .A(n2859), .B(n2827), .Z(n2860) );
  HS65_LH_NOR3X4 U828 ( .A(n775), .B(n774), .C(n778), .Z(n1330) );
  HS65_LH_NOR3X4 U829 ( .A(n769), .B(n770), .C(n773), .Z(n2819) );
  HS65_LH_NOR2X6 U830 ( .A(n776), .B(n777), .Z(n1323) );
  HS65_LH_NOR2X6 U831 ( .A(n771), .B(n772), .Z(n2806) );
  HS65_LH_OAI22X6 U832 ( .A(n6469), .B(n406), .C(n6466), .D(n374), .Z(n1312)
         );
  HS65_LH_BFX9 U833 ( .A(n847), .Z(n6531) );
  HS65_LH_BFX9 U834 ( .A(n847), .Z(n6530) );
  HS65_LH_BFX9 U835 ( .A(n848), .Z(n6525) );
  HS65_LH_BFX9 U836 ( .A(n848), .Z(n6527) );
  HS65_LH_BFX9 U837 ( .A(n848), .Z(n6526) );
  HS65_LH_BFX9 U838 ( .A(n847), .Z(n6528) );
  HS65_LH_BFX9 U839 ( .A(n847), .Z(n6529) );
  HS65_LH_BFX9 U840 ( .A(n847), .Z(n6532) );
  HS65_LH_BFX9 U841 ( .A(n848), .Z(n6523) );
  HS65_LH_BFX9 U842 ( .A(n848), .Z(n6524) );
  HS65_LH_OAI21X3 U843 ( .A(n6525), .B(n846), .C(n1314), .Z(
        \regfile_o[READ_DATA1][0] ) );
  HS65_LH_OAI21X3 U844 ( .A(n1315), .B(n1316), .C(n6523), .Z(n1314) );
  HS65_LH_NAND4ABX3 U845 ( .A(n1317), .B(n1318), .C(n1319), .D(n1320), .Z(
        n1316) );
  HS65_LH_NAND4ABX3 U846 ( .A(n1332), .B(n1333), .C(n1334), .D(n1335), .Z(
        n1315) );
  HS65_LH_OAI21X3 U847 ( .A(n6527), .B(n845), .C(n1160), .Z(
        \regfile_o[READ_DATA1][1] ) );
  HS65_LH_OAI21X3 U848 ( .A(n1161), .B(n1162), .C(n6524), .Z(n1160) );
  HS65_LH_NAND4ABX3 U849 ( .A(n1163), .B(n1164), .C(n1165), .D(n1166), .Z(
        n1162) );
  HS65_LH_NAND4ABX3 U850 ( .A(n1168), .B(n1169), .C(n1170), .D(n1171), .Z(
        n1161) );
  HS65_LH_OAI21X3 U851 ( .A(n6526), .B(n844), .C(n1006), .Z(
        \regfile_o[READ_DATA1][2] ) );
  HS65_LH_OAI21X3 U852 ( .A(n1007), .B(n1008), .C(n6525), .Z(n1006) );
  HS65_LH_NAND4ABX3 U853 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .Z(
        n1008) );
  HS65_LH_NAND4ABX3 U854 ( .A(n1014), .B(n1015), .C(n1016), .D(n1017), .Z(
        n1007) );
  HS65_LH_OAI21X3 U855 ( .A(n6525), .B(n843), .C(n964), .Z(
        \regfile_o[READ_DATA1][3] ) );
  HS65_LH_OAI21X3 U856 ( .A(n965), .B(n966), .C(n6524), .Z(n964) );
  HS65_LH_NAND4ABX3 U857 ( .A(n967), .B(n968), .C(n969), .D(n970), .Z(n966) );
  HS65_LH_NAND4ABX3 U858 ( .A(n972), .B(n973), .C(n974), .D(n975), .Z(n965) );
  HS65_LH_OAI21X3 U859 ( .A(n6526), .B(n842), .C(n950), .Z(
        \regfile_o[READ_DATA1][4] ) );
  HS65_LH_OAI21X3 U860 ( .A(n951), .B(n952), .C(n6524), .Z(n950) );
  HS65_LH_NAND4ABX3 U861 ( .A(n953), .B(n954), .C(n955), .D(n956), .Z(n952) );
  HS65_LH_NAND4ABX3 U862 ( .A(n958), .B(n959), .C(n960), .D(n961), .Z(n951) );
  HS65_LH_OAI21X3 U863 ( .A(n6525), .B(n841), .C(n936), .Z(
        \regfile_o[READ_DATA1][5] ) );
  HS65_LH_OAI21X3 U864 ( .A(n937), .B(n938), .C(n6524), .Z(n936) );
  HS65_LH_NAND4ABX3 U865 ( .A(n939), .B(n940), .C(n941), .D(n942), .Z(n938) );
  HS65_LH_NAND4ABX3 U866 ( .A(n944), .B(n945), .C(n946), .D(n947), .Z(n937) );
  HS65_LH_OAI21X3 U867 ( .A(n6525), .B(n840), .C(n922), .Z(
        \regfile_o[READ_DATA1][6] ) );
  HS65_LH_OAI21X3 U868 ( .A(n923), .B(n924), .C(n6523), .Z(n922) );
  HS65_LH_NAND4ABX3 U869 ( .A(n925), .B(n926), .C(n927), .D(n928), .Z(n924) );
  HS65_LH_NAND4ABX3 U870 ( .A(n930), .B(n931), .C(n932), .D(n933), .Z(n923) );
  HS65_LH_OAI21X3 U871 ( .A(n6526), .B(n839), .C(n908), .Z(
        \regfile_o[READ_DATA1][7] ) );
  HS65_LH_OAI21X3 U872 ( .A(n909), .B(n910), .C(n6523), .Z(n908) );
  HS65_LH_NAND4ABX3 U873 ( .A(n911), .B(n912), .C(n913), .D(n914), .Z(n910) );
  HS65_LH_NAND4ABX3 U874 ( .A(n916), .B(n917), .C(n918), .D(n919), .Z(n909) );
  HS65_LH_OAI21X3 U875 ( .A(n6525), .B(n838), .C(n894), .Z(
        \regfile_o[READ_DATA1][8] ) );
  HS65_LH_OAI21X3 U876 ( .A(n895), .B(n896), .C(n6523), .Z(n894) );
  HS65_LH_NAND4ABX3 U877 ( .A(n897), .B(n898), .C(n899), .D(n900), .Z(n896) );
  HS65_LH_NAND4ABX3 U878 ( .A(n902), .B(n903), .C(n904), .D(n905), .Z(n895) );
  HS65_LH_OAI21X3 U879 ( .A(n6526), .B(n837), .C(n849), .Z(
        \regfile_o[READ_DATA1][9] ) );
  HS65_LH_OAI21X3 U880 ( .A(n850), .B(n851), .C(n6523), .Z(n849) );
  HS65_LH_NAND4ABX3 U881 ( .A(n852), .B(n853), .C(n854), .D(n855), .Z(n851) );
  HS65_LH_NAND4ABX3 U882 ( .A(n872), .B(n873), .C(n874), .D(n875), .Z(n850) );
  HS65_LH_OAI21X3 U883 ( .A(n848), .B(n836), .C(n1300), .Z(
        \regfile_o[READ_DATA1][10] ) );
  HS65_LH_OAI21X3 U884 ( .A(n1301), .B(n1302), .C(n6523), .Z(n1300) );
  HS65_LH_NAND4ABX3 U885 ( .A(n1303), .B(n1304), .C(n1305), .D(n1306), .Z(
        n1302) );
  HS65_LH_OAI21X3 U886 ( .A(n6527), .B(n835), .C(n1286), .Z(
        \regfile_o[READ_DATA1][11] ) );
  HS65_LH_OAI21X3 U887 ( .A(n1287), .B(n1288), .C(n6523), .Z(n1286) );
  HS65_LH_NAND4ABX3 U888 ( .A(n1289), .B(n1290), .C(n1291), .D(n1292), .Z(
        n1288) );
  HS65_LH_NAND4ABX3 U889 ( .A(n1294), .B(n1295), .C(n1296), .D(n1297), .Z(
        n1287) );
  HS65_LH_OAI21X3 U890 ( .A(n6527), .B(n834), .C(n1272), .Z(
        \regfile_o[READ_DATA1][12] ) );
  HS65_LH_OAI21X3 U891 ( .A(n1273), .B(n1274), .C(n6523), .Z(n1272) );
  HS65_LH_NAND4ABX3 U892 ( .A(n1275), .B(n1276), .C(n1277), .D(n1278), .Z(
        n1274) );
  HS65_LH_NAND4ABX3 U893 ( .A(n1280), .B(n1281), .C(n1282), .D(n1283), .Z(
        n1273) );
  HS65_LH_OAI21X3 U894 ( .A(n6527), .B(n833), .C(n1258), .Z(
        \regfile_o[READ_DATA1][13] ) );
  HS65_LH_OAI21X3 U895 ( .A(n1259), .B(n1260), .C(n6523), .Z(n1258) );
  HS65_LH_NAND4ABX3 U896 ( .A(n1261), .B(n1262), .C(n1263), .D(n1264), .Z(
        n1260) );
  HS65_LH_NAND4ABX3 U897 ( .A(n1266), .B(n1267), .C(n1268), .D(n1269), .Z(
        n1259) );
  HS65_LH_OAI21X3 U898 ( .A(n6527), .B(n832), .C(n1244), .Z(
        \regfile_o[READ_DATA1][14] ) );
  HS65_LH_OAI21X3 U899 ( .A(n1245), .B(n1246), .C(n6523), .Z(n1244) );
  HS65_LH_NAND4ABX3 U900 ( .A(n1247), .B(n1248), .C(n1249), .D(n1250), .Z(
        n1246) );
  HS65_LH_NAND4ABX3 U901 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .Z(
        n1245) );
  HS65_LH_OAI21X3 U902 ( .A(n6527), .B(n831), .C(n1230), .Z(
        \regfile_o[READ_DATA1][15] ) );
  HS65_LH_OAI21X3 U903 ( .A(n1231), .B(n1232), .C(n6523), .Z(n1230) );
  HS65_LH_NAND4ABX3 U904 ( .A(n1233), .B(n1234), .C(n1235), .D(n1236), .Z(
        n1232) );
  HS65_LH_NAND4ABX3 U905 ( .A(n1238), .B(n1239), .C(n1240), .D(n1241), .Z(
        n1231) );
  HS65_LH_OAI21X3 U906 ( .A(n6527), .B(n830), .C(n1216), .Z(
        \regfile_o[READ_DATA1][16] ) );
  HS65_LH_OAI21X3 U907 ( .A(n1217), .B(n1218), .C(n6523), .Z(n1216) );
  HS65_LH_NAND4ABX3 U908 ( .A(n1219), .B(n1220), .C(n1221), .D(n1222), .Z(
        n1218) );
  HS65_LH_NAND4ABX3 U909 ( .A(n1224), .B(n1225), .C(n1226), .D(n1227), .Z(
        n1217) );
  HS65_LH_OAI21X3 U910 ( .A(n6527), .B(n829), .C(n1202), .Z(
        \regfile_o[READ_DATA1][17] ) );
  HS65_LH_OAI21X3 U911 ( .A(n1203), .B(n1204), .C(n6524), .Z(n1202) );
  HS65_LH_NAND4ABX3 U912 ( .A(n1205), .B(n1206), .C(n1207), .D(n1208), .Z(
        n1204) );
  HS65_LH_NAND4ABX3 U913 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .Z(
        n1203) );
  HS65_LH_OAI21X3 U914 ( .A(n6527), .B(n828), .C(n1188), .Z(
        \regfile_o[READ_DATA1][18] ) );
  HS65_LH_OAI21X3 U915 ( .A(n1189), .B(n1190), .C(n6524), .Z(n1188) );
  HS65_LH_NAND4ABX3 U916 ( .A(n1191), .B(n1192), .C(n1193), .D(n1194), .Z(
        n1190) );
  HS65_LH_NAND4ABX3 U917 ( .A(n1196), .B(n1197), .C(n1198), .D(n1199), .Z(
        n1189) );
  HS65_LH_OAI21X3 U918 ( .A(n6527), .B(n827), .C(n1174), .Z(
        \regfile_o[READ_DATA1][19] ) );
  HS65_LH_OAI21X3 U919 ( .A(n1175), .B(n1176), .C(n6524), .Z(n1174) );
  HS65_LH_NAND4ABX3 U920 ( .A(n1177), .B(n1178), .C(n1179), .D(n1180), .Z(
        n1176) );
  HS65_LH_NAND4ABX3 U921 ( .A(n1182), .B(n1183), .C(n1184), .D(n1185), .Z(
        n1175) );
  HS65_LH_OAI21X3 U922 ( .A(n6527), .B(n826), .C(n1146), .Z(
        \regfile_o[READ_DATA1][20] ) );
  HS65_LH_OAI21X3 U923 ( .A(n1147), .B(n1148), .C(n6524), .Z(n1146) );
  HS65_LH_NAND4ABX3 U924 ( .A(n1149), .B(n1150), .C(n1151), .D(n1152), .Z(
        n1148) );
  HS65_LH_NAND4ABX3 U925 ( .A(n1154), .B(n1155), .C(n1156), .D(n1157), .Z(
        n1147) );
  HS65_LH_OAI21X3 U926 ( .A(n6527), .B(n825), .C(n1132), .Z(
        \regfile_o[READ_DATA1][21] ) );
  HS65_LH_OAI21X3 U927 ( .A(n1133), .B(n1134), .C(n6524), .Z(n1132) );
  HS65_LH_NAND4ABX3 U928 ( .A(n1135), .B(n1136), .C(n1137), .D(n1138), .Z(
        n1134) );
  HS65_LH_NAND4ABX3 U929 ( .A(n1140), .B(n1141), .C(n1142), .D(n1143), .Z(
        n1133) );
  HS65_LH_OAI21X3 U930 ( .A(n6527), .B(n824), .C(n1118), .Z(
        \regfile_o[READ_DATA1][22] ) );
  HS65_LH_OAI21X3 U931 ( .A(n1119), .B(n1120), .C(n6524), .Z(n1118) );
  HS65_LH_NAND4ABX3 U932 ( .A(n1121), .B(n1122), .C(n1123), .D(n1124), .Z(
        n1120) );
  HS65_LH_NAND4ABX3 U933 ( .A(n1126), .B(n1127), .C(n1128), .D(n1129), .Z(
        n1119) );
  HS65_LH_OAI21X3 U934 ( .A(n6526), .B(n823), .C(n1104), .Z(
        \regfile_o[READ_DATA1][23] ) );
  HS65_LH_OAI21X3 U935 ( .A(n1105), .B(n1106), .C(n6524), .Z(n1104) );
  HS65_LH_NAND4ABX3 U936 ( .A(n1107), .B(n1108), .C(n1109), .D(n1110), .Z(
        n1106) );
  HS65_LH_NAND4ABX3 U937 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .Z(
        n1105) );
  HS65_LH_OAI21X3 U938 ( .A(n6526), .B(n822), .C(n1090), .Z(
        \regfile_o[READ_DATA1][24] ) );
  HS65_LH_OAI21X3 U939 ( .A(n1091), .B(n1092), .C(n6525), .Z(n1090) );
  HS65_LH_NAND4ABX3 U940 ( .A(n1093), .B(n1094), .C(n1095), .D(n1096), .Z(
        n1092) );
  HS65_LH_NAND4ABX3 U941 ( .A(n1098), .B(n1099), .C(n1100), .D(n1101), .Z(
        n1091) );
  HS65_LH_OAI21X3 U942 ( .A(n6526), .B(n821), .C(n1076), .Z(
        \regfile_o[READ_DATA1][25] ) );
  HS65_LH_OAI21X3 U943 ( .A(n1077), .B(n1078), .C(n6525), .Z(n1076) );
  HS65_LH_NAND4ABX3 U944 ( .A(n1079), .B(n1080), .C(n1081), .D(n1082), .Z(
        n1078) );
  HS65_LH_NAND4ABX3 U945 ( .A(n1084), .B(n1085), .C(n1086), .D(n1087), .Z(
        n1077) );
  HS65_LH_OAI21X3 U946 ( .A(n6526), .B(n820), .C(n1062), .Z(
        \regfile_o[READ_DATA1][26] ) );
  HS65_LH_OAI21X3 U947 ( .A(n1063), .B(n1064), .C(n6524), .Z(n1062) );
  HS65_LH_NAND4ABX3 U948 ( .A(n1065), .B(n1066), .C(n1067), .D(n1068), .Z(
        n1064) );
  HS65_LH_NAND4ABX3 U949 ( .A(n1070), .B(n1071), .C(n1072), .D(n1073), .Z(
        n1063) );
  HS65_LH_OAI21X3 U950 ( .A(n6526), .B(n819), .C(n1048), .Z(
        \regfile_o[READ_DATA1][27] ) );
  HS65_LH_OAI21X3 U951 ( .A(n1049), .B(n1050), .C(n6525), .Z(n1048) );
  HS65_LH_NAND4ABX3 U952 ( .A(n1051), .B(n1052), .C(n1053), .D(n1054), .Z(
        n1050) );
  HS65_LH_NAND4ABX3 U953 ( .A(n1056), .B(n1057), .C(n1058), .D(n1059), .Z(
        n1049) );
  HS65_LH_OAI21X3 U954 ( .A(n6526), .B(n818), .C(n1034), .Z(
        \regfile_o[READ_DATA1][28] ) );
  HS65_LH_OAI21X3 U955 ( .A(n1035), .B(n1036), .C(n6525), .Z(n1034) );
  HS65_LH_NAND4ABX3 U956 ( .A(n1037), .B(n1038), .C(n1039), .D(n1040), .Z(
        n1036) );
  HS65_LH_NAND4ABX3 U957 ( .A(n1042), .B(n1043), .C(n1044), .D(n1045), .Z(
        n1035) );
  HS65_LH_OAI21X3 U958 ( .A(n6526), .B(n817), .C(n1020), .Z(
        \regfile_o[READ_DATA1][29] ) );
  HS65_LH_OAI21X3 U959 ( .A(n1021), .B(n1022), .C(n6525), .Z(n1020) );
  HS65_LH_NAND4ABX3 U960 ( .A(n1023), .B(n1024), .C(n1025), .D(n1026), .Z(
        n1022) );
  HS65_LH_NAND4ABX3 U961 ( .A(n1028), .B(n1029), .C(n1030), .D(n1031), .Z(
        n1021) );
  HS65_LH_OAI21X3 U962 ( .A(n6526), .B(n816), .C(n992), .Z(
        \regfile_o[READ_DATA1][30] ) );
  HS65_LH_OAI21X3 U963 ( .A(n993), .B(n994), .C(n6525), .Z(n992) );
  HS65_LH_NAND4ABX3 U964 ( .A(n995), .B(n996), .C(n997), .D(n998), .Z(n994) );
  HS65_LH_NAND4ABX3 U965 ( .A(n1000), .B(n1001), .C(n1002), .D(n1003), .Z(n993) );
  HS65_LH_OAI21X3 U966 ( .A(n6526), .B(n815), .C(n978), .Z(
        \regfile_o[READ_DATA1][31] ) );
  HS65_LH_OAI21X3 U967 ( .A(n979), .B(n980), .C(n6525), .Z(n978) );
  HS65_LH_NAND4ABX3 U968 ( .A(n981), .B(n982), .C(n983), .D(n984), .Z(n980) );
  HS65_LH_NAND4ABX3 U969 ( .A(n986), .B(n987), .C(n988), .D(n989), .Z(n979) );
  HS65_LH_OAI21X3 U970 ( .A(n844), .B(n6531), .C(n2489), .Z(
        \regfile_o[READ_DATA0][2] ) );
  HS65_LH_OAI21X3 U971 ( .A(n2490), .B(n2491), .C(n6530), .Z(n2489) );
  HS65_LH_NAND4ABX3 U972 ( .A(n2492), .B(n2493), .C(n2494), .D(n2495), .Z(
        n2491) );
  HS65_LH_NAND4ABX3 U973 ( .A(n2497), .B(n2498), .C(n2499), .D(n2500), .Z(
        n2490) );
  HS65_LH_OAI21X3 U974 ( .A(n842), .B(n6531), .C(n2433), .Z(
        \regfile_o[READ_DATA0][4] ) );
  HS65_LH_OAI21X3 U975 ( .A(n2434), .B(n2435), .C(n6529), .Z(n2433) );
  HS65_LH_NAND4ABX3 U976 ( .A(n2436), .B(n2437), .C(n2438), .D(n2439), .Z(
        n2435) );
  HS65_LH_NAND4ABX3 U977 ( .A(n2441), .B(n2442), .C(n2443), .D(n2444), .Z(
        n2434) );
  HS65_LH_OAI21X3 U978 ( .A(n839), .B(n6531), .C(n1399), .Z(
        \regfile_o[READ_DATA0][7] ) );
  HS65_LH_OAI21X3 U979 ( .A(n1400), .B(n1401), .C(n6528), .Z(n1399) );
  HS65_LH_NAND4ABX3 U980 ( .A(n1402), .B(n1403), .C(n1404), .D(n1405), .Z(
        n1401) );
  HS65_LH_NAND4ABX3 U981 ( .A(n1407), .B(n1408), .C(n1409), .D(n1410), .Z(
        n1400) );
  HS65_LH_OAI21X3 U982 ( .A(n837), .B(n6531), .C(n1340), .Z(
        \regfile_o[READ_DATA0][9] ) );
  HS65_LH_OAI21X3 U983 ( .A(n1341), .B(n1342), .C(n6528), .Z(n1340) );
  HS65_LH_NAND4ABX3 U984 ( .A(n1343), .B(n1344), .C(n1345), .D(n1346), .Z(
        n1342) );
  HS65_LH_NAND4ABX3 U985 ( .A(n1363), .B(n1364), .C(n1365), .D(n1366), .Z(
        n1341) );
  HS65_LH_OAI21X3 U986 ( .A(n824), .B(n6531), .C(n2601), .Z(
        \regfile_o[READ_DATA0][22] ) );
  HS65_LH_OAI21X3 U987 ( .A(n2602), .B(n2603), .C(n6529), .Z(n2601) );
  HS65_LH_NAND4ABX3 U988 ( .A(n2604), .B(n2605), .C(n2606), .D(n2607), .Z(
        n2603) );
  HS65_LH_NAND4ABX3 U989 ( .A(n2609), .B(n2610), .C(n2611), .D(n2612), .Z(
        n2602) );
  HS65_LH_OAI21X3 U990 ( .A(n823), .B(n6531), .C(n2587), .Z(
        \regfile_o[READ_DATA0][23] ) );
  HS65_LH_OAI21X3 U991 ( .A(n2588), .B(n2589), .C(n6529), .Z(n2587) );
  HS65_LH_NAND4ABX3 U992 ( .A(n2590), .B(n2591), .C(n2592), .D(n2593), .Z(
        n2589) );
  HS65_LH_NAND4ABX3 U993 ( .A(n2595), .B(n2596), .C(n2597), .D(n2598), .Z(
        n2588) );
  HS65_LH_OAI21X3 U994 ( .A(n822), .B(n6531), .C(n2573), .Z(
        \regfile_o[READ_DATA0][24] ) );
  HS65_LH_OAI21X3 U995 ( .A(n2574), .B(n2575), .C(n6530), .Z(n2573) );
  HS65_LH_NAND4ABX3 U996 ( .A(n2576), .B(n2577), .C(n2578), .D(n2579), .Z(
        n2575) );
  HS65_LH_NAND4ABX3 U997 ( .A(n2581), .B(n2582), .C(n2583), .D(n2584), .Z(
        n2574) );
  HS65_LH_OAI21X3 U998 ( .A(n821), .B(n6531), .C(n2559), .Z(
        \regfile_o[READ_DATA0][25] ) );
  HS65_LH_OAI21X3 U999 ( .A(n2560), .B(n2561), .C(n6530), .Z(n2559) );
  HS65_LH_NAND4ABX3 U1000 ( .A(n2562), .B(n2563), .C(n2564), .D(n2565), .Z(
        n2561) );
  HS65_LH_NAND4ABX3 U1001 ( .A(n2567), .B(n2568), .C(n2569), .D(n2570), .Z(
        n2560) );
  HS65_LH_OAI21X3 U1002 ( .A(n820), .B(n6531), .C(n2545), .Z(
        \regfile_o[READ_DATA0][26] ) );
  HS65_LH_OAI21X3 U1003 ( .A(n2546), .B(n2547), .C(n6529), .Z(n2545) );
  HS65_LH_NAND4ABX3 U1004 ( .A(n2548), .B(n2549), .C(n2550), .D(n2551), .Z(
        n2547) );
  HS65_LH_NAND4ABX3 U1005 ( .A(n2553), .B(n2554), .C(n2555), .D(n2556), .Z(
        n2546) );
  HS65_LH_OAI21X3 U1006 ( .A(n819), .B(n6531), .C(n2531), .Z(
        \regfile_o[READ_DATA0][27] ) );
  HS65_LH_OAI21X3 U1007 ( .A(n2532), .B(n2533), .C(n6530), .Z(n2531) );
  HS65_LH_NAND4ABX3 U1008 ( .A(n2534), .B(n2535), .C(n2536), .D(n2537), .Z(
        n2533) );
  HS65_LH_NAND4ABX3 U1009 ( .A(n2539), .B(n2540), .C(n2541), .D(n2542), .Z(
        n2532) );
  HS65_LH_OAI21X3 U1010 ( .A(n818), .B(n6531), .C(n2517), .Z(
        \regfile_o[READ_DATA0][28] ) );
  HS65_LH_OAI21X3 U1011 ( .A(n2518), .B(n2519), .C(n6530), .Z(n2517) );
  HS65_LH_NAND4ABX3 U1012 ( .A(n2520), .B(n2521), .C(n2522), .D(n2523), .Z(
        n2519) );
  HS65_LH_NAND4ABX3 U1013 ( .A(n2525), .B(n2526), .C(n2527), .D(n2528), .Z(
        n2518) );
  HS65_LH_OAI21X3 U1014 ( .A(n817), .B(n6531), .C(n2503), .Z(
        \regfile_o[READ_DATA0][29] ) );
  HS65_LH_OAI21X3 U1015 ( .A(n2504), .B(n2505), .C(n6530), .Z(n2503) );
  HS65_LH_NAND4ABX3 U1016 ( .A(n2506), .B(n2507), .C(n2508), .D(n2509), .Z(
        n2505) );
  HS65_LH_NAND4ABX3 U1017 ( .A(n2511), .B(n2512), .C(n2513), .D(n2514), .Z(
        n2504) );
  HS65_LH_OAI21X3 U1018 ( .A(n816), .B(n6531), .C(n2475), .Z(
        \regfile_o[READ_DATA0][30] ) );
  HS65_LH_OAI21X3 U1019 ( .A(n2476), .B(n2477), .C(n6530), .Z(n2475) );
  HS65_LH_NAND4ABX3 U1020 ( .A(n2478), .B(n2479), .C(n2480), .D(n2481), .Z(
        n2477) );
  HS65_LH_NAND4ABX3 U1021 ( .A(n2483), .B(n2484), .C(n2485), .D(n2486), .Z(
        n2476) );
  HS65_LH_OAI21X3 U1022 ( .A(n815), .B(n6531), .C(n2461), .Z(
        \regfile_o[READ_DATA0][31] ) );
  HS65_LH_OAI21X3 U1023 ( .A(n2462), .B(n2463), .C(n6530), .Z(n2461) );
  HS65_LH_NAND4ABX3 U1024 ( .A(n2464), .B(n2465), .C(n2466), .D(n2467), .Z(
        n2463) );
  HS65_LH_NAND4ABX3 U1025 ( .A(n2469), .B(n2470), .C(n2471), .D(n2472), .Z(
        n2462) );
  HS65_LH_OAI21X3 U1026 ( .A(n846), .B(n6530), .C(n2797), .Z(
        \regfile_o[READ_DATA0][0] ) );
  HS65_LH_OAI21X3 U1027 ( .A(n2798), .B(n2799), .C(n6528), .Z(n2797) );
  HS65_LH_NAND4ABX3 U1028 ( .A(n2800), .B(n2801), .C(n2802), .D(n2803), .Z(
        n2799) );
  HS65_LH_NAND4ABX3 U1029 ( .A(n2814), .B(n2815), .C(n2816), .D(n2817), .Z(
        n2798) );
  HS65_LH_OAI21X3 U1030 ( .A(n843), .B(n6530), .C(n2447), .Z(
        \regfile_o[READ_DATA0][3] ) );
  HS65_LH_OAI21X3 U1031 ( .A(n2448), .B(n2449), .C(n6529), .Z(n2447) );
  HS65_LH_NAND4ABX3 U1032 ( .A(n2450), .B(n2451), .C(n2452), .D(n2453), .Z(
        n2449) );
  HS65_LH_NAND4ABX3 U1033 ( .A(n2455), .B(n2456), .C(n2457), .D(n2458), .Z(
        n2448) );
  HS65_LH_OAI21X3 U1034 ( .A(n841), .B(n6530), .C(n1427), .Z(
        \regfile_o[READ_DATA0][5] ) );
  HS65_LH_OAI21X3 U1035 ( .A(n1428), .B(n1429), .C(n6529), .Z(n1427) );
  HS65_LH_NAND4ABX3 U1036 ( .A(n1430), .B(n1431), .C(n1432), .D(n1433), .Z(
        n1429) );
  HS65_LH_NAND4ABX3 U1037 ( .A(n2427), .B(n2428), .C(n2429), .D(n2430), .Z(
        n1428) );
  HS65_LH_OAI21X3 U1038 ( .A(n840), .B(n6530), .C(n1413), .Z(
        \regfile_o[READ_DATA0][6] ) );
  HS65_LH_OAI21X3 U1039 ( .A(n1414), .B(n1415), .C(n6528), .Z(n1413) );
  HS65_LH_NAND4ABX3 U1040 ( .A(n1416), .B(n1417), .C(n1418), .D(n1419), .Z(
        n1415) );
  HS65_LH_NAND4ABX3 U1041 ( .A(n1421), .B(n1422), .C(n1423), .D(n1424), .Z(
        n1414) );
  HS65_LH_OAI21X3 U1042 ( .A(n838), .B(n6530), .C(n1385), .Z(
        \regfile_o[READ_DATA0][8] ) );
  HS65_LH_OAI21X3 U1043 ( .A(n1386), .B(n1387), .C(n6528), .Z(n1385) );
  HS65_LH_NAND4ABX3 U1044 ( .A(n1388), .B(n1389), .C(n1390), .D(n1391), .Z(
        n1387) );
  HS65_LH_NAND4ABX3 U1045 ( .A(n1393), .B(n1394), .C(n1395), .D(n1396), .Z(
        n1386) );
  HS65_LH_OAI21X3 U1046 ( .A(n845), .B(n6532), .C(n2643), .Z(
        \regfile_o[READ_DATA0][1] ) );
  HS65_LH_OAI21X3 U1047 ( .A(n2644), .B(n2645), .C(n6529), .Z(n2643) );
  HS65_LH_NAND4ABX3 U1048 ( .A(n2646), .B(n2647), .C(n2648), .D(n2649), .Z(
        n2645) );
  HS65_LH_NAND4ABX3 U1049 ( .A(n2651), .B(n2652), .C(n2653), .D(n2654), .Z(
        n2644) );
  HS65_LH_OAI21X3 U1050 ( .A(n836), .B(n6532), .C(n2783), .Z(
        \regfile_o[READ_DATA0][10] ) );
  HS65_LH_OAI21X3 U1051 ( .A(n2784), .B(n2785), .C(n6528), .Z(n2783) );
  HS65_LH_NAND4ABX3 U1052 ( .A(n2786), .B(n2787), .C(n2788), .D(n2789), .Z(
        n2785) );
  HS65_LH_NAND4ABX3 U1053 ( .A(n2791), .B(n2792), .C(n2793), .D(n2794), .Z(
        n2784) );
  HS65_LH_OAI21X3 U1054 ( .A(n835), .B(n6532), .C(n2769), .Z(
        \regfile_o[READ_DATA0][11] ) );
  HS65_LH_OAI21X3 U1055 ( .A(n2770), .B(n2771), .C(n6528), .Z(n2769) );
  HS65_LH_NAND4ABX3 U1056 ( .A(n2772), .B(n2773), .C(n2774), .D(n2775), .Z(
        n2771) );
  HS65_LH_NAND4ABX3 U1057 ( .A(n2777), .B(n2778), .C(n2779), .D(n2780), .Z(
        n2770) );
  HS65_LH_OAI21X3 U1058 ( .A(n834), .B(n6532), .C(n2755), .Z(
        \regfile_o[READ_DATA0][12] ) );
  HS65_LH_OAI21X3 U1059 ( .A(n2756), .B(n2757), .C(n6528), .Z(n2755) );
  HS65_LH_NAND4ABX3 U1060 ( .A(n2758), .B(n2759), .C(n2760), .D(n2761), .Z(
        n2757) );
  HS65_LH_NAND4ABX3 U1061 ( .A(n2763), .B(n2764), .C(n2765), .D(n2766), .Z(
        n2756) );
  HS65_LH_OAI21X3 U1062 ( .A(n833), .B(n6532), .C(n2741), .Z(
        \regfile_o[READ_DATA0][13] ) );
  HS65_LH_OAI21X3 U1063 ( .A(n2742), .B(n2743), .C(n6528), .Z(n2741) );
  HS65_LH_NAND4ABX3 U1064 ( .A(n2744), .B(n2745), .C(n2746), .D(n2747), .Z(
        n2743) );
  HS65_LH_NAND4ABX3 U1065 ( .A(n2749), .B(n2750), .C(n2751), .D(n2752), .Z(
        n2742) );
  HS65_LH_OAI21X3 U1066 ( .A(n832), .B(n6532), .C(n2727), .Z(
        \regfile_o[READ_DATA0][14] ) );
  HS65_LH_OAI21X3 U1067 ( .A(n2728), .B(n2729), .C(n6528), .Z(n2727) );
  HS65_LH_NAND4ABX3 U1068 ( .A(n2730), .B(n2731), .C(n2732), .D(n2733), .Z(
        n2729) );
  HS65_LH_NAND4ABX3 U1069 ( .A(n2735), .B(n2736), .C(n2737), .D(n2738), .Z(
        n2728) );
  HS65_LH_OAI21X3 U1070 ( .A(n831), .B(n6532), .C(n2713), .Z(
        \regfile_o[READ_DATA0][15] ) );
  HS65_LH_OAI21X3 U1071 ( .A(n2714), .B(n2715), .C(n6528), .Z(n2713) );
  HS65_LH_NAND4ABX3 U1072 ( .A(n2716), .B(n2717), .C(n2718), .D(n2719), .Z(
        n2715) );
  HS65_LH_NAND4ABX3 U1073 ( .A(n2721), .B(n2722), .C(n2723), .D(n2724), .Z(
        n2714) );
  HS65_LH_OAI21X3 U1074 ( .A(n830), .B(n6532), .C(n2699), .Z(
        \regfile_o[READ_DATA0][16] ) );
  HS65_LH_OAI21X3 U1075 ( .A(n2700), .B(n2701), .C(n6528), .Z(n2699) );
  HS65_LH_NAND4ABX3 U1076 ( .A(n2702), .B(n2703), .C(n2704), .D(n2705), .Z(
        n2701) );
  HS65_LH_NAND4ABX3 U1077 ( .A(n2707), .B(n2708), .C(n2709), .D(n2710), .Z(
        n2700) );
  HS65_LH_OAI21X3 U1078 ( .A(n829), .B(n6532), .C(n2685), .Z(
        \regfile_o[READ_DATA0][17] ) );
  HS65_LH_OAI21X3 U1079 ( .A(n2686), .B(n2687), .C(n6529), .Z(n2685) );
  HS65_LH_NAND4ABX3 U1080 ( .A(n2688), .B(n2689), .C(n2690), .D(n2691), .Z(
        n2687) );
  HS65_LH_NAND4ABX3 U1081 ( .A(n2693), .B(n2694), .C(n2695), .D(n2696), .Z(
        n2686) );
  HS65_LH_OAI21X3 U1082 ( .A(n828), .B(n6532), .C(n2671), .Z(
        \regfile_o[READ_DATA0][18] ) );
  HS65_LH_OAI21X3 U1083 ( .A(n2672), .B(n2673), .C(n6529), .Z(n2671) );
  HS65_LH_NAND4ABX3 U1084 ( .A(n2674), .B(n2675), .C(n2676), .D(n2677), .Z(
        n2673) );
  HS65_LH_NAND4ABX3 U1085 ( .A(n2679), .B(n2680), .C(n2681), .D(n2682), .Z(
        n2672) );
  HS65_LH_OAI21X3 U1086 ( .A(n827), .B(n6532), .C(n2657), .Z(
        \regfile_o[READ_DATA0][19] ) );
  HS65_LH_OAI21X3 U1087 ( .A(n2658), .B(n2659), .C(n6529), .Z(n2657) );
  HS65_LH_NAND4ABX3 U1088 ( .A(n2660), .B(n2661), .C(n2662), .D(n2663), .Z(
        n2659) );
  HS65_LH_NAND4ABX3 U1089 ( .A(n2665), .B(n2666), .C(n2667), .D(n2668), .Z(
        n2658) );
  HS65_LH_OAI21X3 U1090 ( .A(n826), .B(n6532), .C(n2629), .Z(
        \regfile_o[READ_DATA0][20] ) );
  HS65_LH_OAI21X3 U1091 ( .A(n2630), .B(n2631), .C(n6529), .Z(n2629) );
  HS65_LH_NAND4ABX3 U1092 ( .A(n2632), .B(n2633), .C(n2634), .D(n2635), .Z(
        n2631) );
  HS65_LH_NAND4ABX3 U1093 ( .A(n2637), .B(n2638), .C(n2639), .D(n2640), .Z(
        n2630) );
  HS65_LH_OAI21X3 U1094 ( .A(n825), .B(n6532), .C(n2615), .Z(
        \regfile_o[READ_DATA0][21] ) );
  HS65_LH_OAI21X3 U1095 ( .A(n2616), .B(n2617), .C(n6529), .Z(n2615) );
  HS65_LH_NAND4ABX3 U1096 ( .A(n2618), .B(n2619), .C(n2620), .D(n2621), .Z(
        n2617) );
  HS65_LH_NAND4ABX3 U1097 ( .A(n2623), .B(n2624), .C(n2625), .D(n2626), .Z(
        n2616) );
  HS65_LH_BFX9 U1098 ( .A(n6536), .Z(n6534) );
  HS65_LH_BFX9 U1099 ( .A(n6536), .Z(n6533) );
  HS65_LH_BFX9 U1100 ( .A(n6536), .Z(n6535) );
  HS65_LH_OAI22X6 U1101 ( .A(n248), .B(n6218), .C(n838), .D(n6220), .Z(n1666)
         );
  HS65_LH_OAI22X6 U1102 ( .A(n247), .B(n6218), .C(n837), .D(n6220), .Z(n1667)
         );
  HS65_LH_OAI22X6 U1103 ( .A(n246), .B(n6218), .C(n836), .D(n6220), .Z(n1668)
         );
  HS65_LH_OAI22X6 U1104 ( .A(n245), .B(n6218), .C(n835), .D(n6220), .Z(n1669)
         );
  HS65_LH_OAI22X6 U1105 ( .A(n244), .B(n6218), .C(n834), .D(n6220), .Z(n1670)
         );
  HS65_LH_OAI22X6 U1106 ( .A(n243), .B(n6218), .C(n833), .D(n6220), .Z(n1671)
         );
  HS65_LH_OAI22X6 U1107 ( .A(n242), .B(n6218), .C(n832), .D(n6220), .Z(n1672)
         );
  HS65_LH_OAI22X6 U1108 ( .A(n241), .B(n6218), .C(n831), .D(n6220), .Z(n1673)
         );
  HS65_LH_OAI22X6 U1109 ( .A(n240), .B(n6218), .C(n830), .D(n6220), .Z(n1674)
         );
  HS65_LH_OAI22X6 U1110 ( .A(n239), .B(n6218), .C(n829), .D(n6220), .Z(n1675)
         );
  HS65_LH_OAI22X6 U1111 ( .A(n238), .B(n6218), .C(n828), .D(n6220), .Z(n1676)
         );
  HS65_LH_OAI22X6 U1112 ( .A(n237), .B(n6218), .C(n827), .D(n6220), .Z(n1677)
         );
  HS65_LH_OAI22X6 U1113 ( .A(n236), .B(n6217), .C(n826), .D(n6221), .Z(n1678)
         );
  HS65_LH_OAI22X6 U1114 ( .A(n235), .B(n6217), .C(n825), .D(n6221), .Z(n1679)
         );
  HS65_LH_OAI22X6 U1115 ( .A(n234), .B(n6217), .C(n824), .D(n6221), .Z(n1680)
         );
  HS65_LH_OAI22X6 U1116 ( .A(n233), .B(n6217), .C(n823), .D(n6221), .Z(n1681)
         );
  HS65_LH_OAI22X6 U1117 ( .A(n232), .B(n6217), .C(n822), .D(n6221), .Z(n1682)
         );
  HS65_LH_OAI22X6 U1118 ( .A(n231), .B(n6217), .C(n821), .D(n6221), .Z(n1683)
         );
  HS65_LH_OAI22X6 U1119 ( .A(n230), .B(n6217), .C(n820), .D(n6221), .Z(n1684)
         );
  HS65_LH_OAI22X6 U1120 ( .A(n229), .B(n6217), .C(n819), .D(n6221), .Z(n1685)
         );
  HS65_LH_OAI22X6 U1121 ( .A(n228), .B(n6217), .C(n818), .D(n6221), .Z(n1686)
         );
  HS65_LH_OAI22X6 U1122 ( .A(n227), .B(n6217), .C(n817), .D(n6221), .Z(n1687)
         );
  HS65_LH_OAI22X6 U1123 ( .A(n226), .B(n6217), .C(n816), .D(n6221), .Z(n1688)
         );
  HS65_LH_OAI22X6 U1124 ( .A(n225), .B(n6217), .C(n815), .D(n6221), .Z(n1689)
         );
  HS65_LH_OAI22X6 U1125 ( .A(n216), .B(n6223), .C(n838), .D(n6225), .Z(n1698)
         );
  HS65_LH_OAI22X6 U1126 ( .A(n215), .B(n6223), .C(n837), .D(n6225), .Z(n1699)
         );
  HS65_LH_OAI22X6 U1127 ( .A(n214), .B(n6223), .C(n836), .D(n6225), .Z(n1700)
         );
  HS65_LH_OAI22X6 U1128 ( .A(n213), .B(n6223), .C(n835), .D(n6225), .Z(n1701)
         );
  HS65_LH_OAI22X6 U1129 ( .A(n212), .B(n6223), .C(n834), .D(n6225), .Z(n1702)
         );
  HS65_LH_OAI22X6 U1130 ( .A(n211), .B(n6223), .C(n833), .D(n6225), .Z(n1703)
         );
  HS65_LH_OAI22X6 U1131 ( .A(n210), .B(n6223), .C(n832), .D(n6225), .Z(n1704)
         );
  HS65_LH_OAI22X6 U1132 ( .A(n209), .B(n6223), .C(n831), .D(n6225), .Z(n1705)
         );
  HS65_LH_OAI22X6 U1133 ( .A(n208), .B(n6223), .C(n830), .D(n6225), .Z(n1706)
         );
  HS65_LH_OAI22X6 U1134 ( .A(n207), .B(n6223), .C(n829), .D(n6225), .Z(n1707)
         );
  HS65_LH_OAI22X6 U1135 ( .A(n206), .B(n6223), .C(n828), .D(n6225), .Z(n1708)
         );
  HS65_LH_OAI22X6 U1136 ( .A(n205), .B(n6223), .C(n827), .D(n6225), .Z(n1709)
         );
  HS65_LH_OAI22X6 U1137 ( .A(n204), .B(n6222), .C(n826), .D(n6226), .Z(n1710)
         );
  HS65_LH_OAI22X6 U1138 ( .A(n203), .B(n6222), .C(n825), .D(n6226), .Z(n1711)
         );
  HS65_LH_OAI22X6 U1139 ( .A(n202), .B(n6222), .C(n824), .D(n6226), .Z(n1712)
         );
  HS65_LH_OAI22X6 U1140 ( .A(n201), .B(n6222), .C(n823), .D(n6226), .Z(n1713)
         );
  HS65_LH_OAI22X6 U1141 ( .A(n200), .B(n6222), .C(n822), .D(n6226), .Z(n1714)
         );
  HS65_LH_OAI22X6 U1142 ( .A(n199), .B(n6222), .C(n821), .D(n6226), .Z(n1715)
         );
  HS65_LH_OAI22X6 U1143 ( .A(n198), .B(n6222), .C(n820), .D(n6226), .Z(n1716)
         );
  HS65_LH_OAI22X6 U1144 ( .A(n197), .B(n6222), .C(n819), .D(n6226), .Z(n1717)
         );
  HS65_LH_OAI22X6 U1145 ( .A(n196), .B(n6222), .C(n818), .D(n6226), .Z(n1718)
         );
  HS65_LH_OAI22X6 U1146 ( .A(n195), .B(n6222), .C(n817), .D(n6226), .Z(n1719)
         );
  HS65_LH_OAI22X6 U1147 ( .A(n194), .B(n6222), .C(n816), .D(n6226), .Z(n1720)
         );
  HS65_LH_OAI22X6 U1148 ( .A(n193), .B(n6222), .C(n815), .D(n6226), .Z(n1721)
         );
  HS65_LH_OAI22X6 U1149 ( .A(n184), .B(n6248), .C(n838), .D(n6250), .Z(n1858)
         );
  HS65_LH_OAI22X6 U1150 ( .A(n183), .B(n6248), .C(n837), .D(n6250), .Z(n1859)
         );
  HS65_LH_OAI22X6 U1151 ( .A(n182), .B(n6248), .C(n836), .D(n6250), .Z(n1860)
         );
  HS65_LH_OAI22X6 U1152 ( .A(n181), .B(n6248), .C(n835), .D(n6250), .Z(n1861)
         );
  HS65_LH_OAI22X6 U1153 ( .A(n180), .B(n6248), .C(n834), .D(n6250), .Z(n1862)
         );
  HS65_LH_OAI22X6 U1154 ( .A(n179), .B(n6248), .C(n833), .D(n6250), .Z(n1863)
         );
  HS65_LH_OAI22X6 U1155 ( .A(n178), .B(n6248), .C(n832), .D(n6250), .Z(n1864)
         );
  HS65_LH_OAI22X6 U1156 ( .A(n177), .B(n6248), .C(n831), .D(n6250), .Z(n1865)
         );
  HS65_LH_OAI22X6 U1157 ( .A(n176), .B(n6248), .C(n830), .D(n6250), .Z(n1866)
         );
  HS65_LH_OAI22X6 U1158 ( .A(n175), .B(n6248), .C(n829), .D(n6250), .Z(n1867)
         );
  HS65_LH_OAI22X6 U1159 ( .A(n174), .B(n6248), .C(n828), .D(n6250), .Z(n1868)
         );
  HS65_LH_OAI22X6 U1160 ( .A(n173), .B(n6248), .C(n827), .D(n6250), .Z(n1869)
         );
  HS65_LH_OAI22X6 U1161 ( .A(n172), .B(n6247), .C(n826), .D(n6251), .Z(n1870)
         );
  HS65_LH_OAI22X6 U1162 ( .A(n171), .B(n6247), .C(n825), .D(n6251), .Z(n1871)
         );
  HS65_LH_OAI22X6 U1163 ( .A(n170), .B(n6247), .C(n824), .D(n6251), .Z(n1872)
         );
  HS65_LH_OAI22X6 U1164 ( .A(n169), .B(n6247), .C(n823), .D(n6251), .Z(n1873)
         );
  HS65_LH_OAI22X6 U1165 ( .A(n168), .B(n6247), .C(n822), .D(n6251), .Z(n1874)
         );
  HS65_LH_OAI22X6 U1166 ( .A(n167), .B(n6247), .C(n821), .D(n6251), .Z(n1875)
         );
  HS65_LH_OAI22X6 U1167 ( .A(n166), .B(n6247), .C(n820), .D(n6251), .Z(n1876)
         );
  HS65_LH_OAI22X6 U1168 ( .A(n165), .B(n6247), .C(n819), .D(n6251), .Z(n1877)
         );
  HS65_LH_OAI22X6 U1169 ( .A(n164), .B(n6247), .C(n818), .D(n6251), .Z(n1878)
         );
  HS65_LH_OAI22X6 U1170 ( .A(n163), .B(n6247), .C(n817), .D(n6251), .Z(n1879)
         );
  HS65_LH_OAI22X6 U1171 ( .A(n162), .B(n6247), .C(n816), .D(n6251), .Z(n1880)
         );
  HS65_LH_OAI22X6 U1172 ( .A(n161), .B(n6247), .C(n815), .D(n6251), .Z(n1881)
         );
  HS65_LH_OAI22X6 U1173 ( .A(n152), .B(n6253), .C(n838), .D(n6255), .Z(n1890)
         );
  HS65_LH_OAI22X6 U1174 ( .A(n151), .B(n6253), .C(n837), .D(n6255), .Z(n1891)
         );
  HS65_LH_OAI22X6 U1175 ( .A(n150), .B(n6253), .C(n836), .D(n6255), .Z(n1892)
         );
  HS65_LH_OAI22X6 U1176 ( .A(n149), .B(n6253), .C(n835), .D(n6255), .Z(n1893)
         );
  HS65_LH_OAI22X6 U1177 ( .A(n148), .B(n6253), .C(n834), .D(n6255), .Z(n1894)
         );
  HS65_LH_OAI22X6 U1178 ( .A(n147), .B(n6253), .C(n833), .D(n6255), .Z(n1895)
         );
  HS65_LH_OAI22X6 U1179 ( .A(n146), .B(n6253), .C(n832), .D(n6255), .Z(n1896)
         );
  HS65_LH_OAI22X6 U1180 ( .A(n145), .B(n6253), .C(n831), .D(n6255), .Z(n1897)
         );
  HS65_LH_OAI22X6 U1181 ( .A(n144), .B(n6253), .C(n830), .D(n6255), .Z(n1898)
         );
  HS65_LH_OAI22X6 U1182 ( .A(n143), .B(n6253), .C(n829), .D(n6255), .Z(n1899)
         );
  HS65_LH_OAI22X6 U1183 ( .A(n142), .B(n6253), .C(n828), .D(n6255), .Z(n1900)
         );
  HS65_LH_OAI22X6 U1184 ( .A(n141), .B(n6253), .C(n827), .D(n6255), .Z(n1901)
         );
  HS65_LH_OAI22X6 U1185 ( .A(n140), .B(n6252), .C(n826), .D(n6256), .Z(n1902)
         );
  HS65_LH_OAI22X6 U1186 ( .A(n139), .B(n6252), .C(n825), .D(n6256), .Z(n1903)
         );
  HS65_LH_OAI22X6 U1187 ( .A(n138), .B(n6252), .C(n824), .D(n6256), .Z(n1904)
         );
  HS65_LH_OAI22X6 U1188 ( .A(n137), .B(n6252), .C(n823), .D(n6256), .Z(n1905)
         );
  HS65_LH_OAI22X6 U1189 ( .A(n136), .B(n6252), .C(n822), .D(n6256), .Z(n1906)
         );
  HS65_LH_OAI22X6 U1190 ( .A(n135), .B(n6252), .C(n821), .D(n6256), .Z(n1907)
         );
  HS65_LH_OAI22X6 U1191 ( .A(n134), .B(n6252), .C(n820), .D(n6256), .Z(n1908)
         );
  HS65_LH_OAI22X6 U1192 ( .A(n133), .B(n6252), .C(n819), .D(n6256), .Z(n1909)
         );
  HS65_LH_OAI22X6 U1193 ( .A(n132), .B(n6252), .C(n818), .D(n6256), .Z(n1910)
         );
  HS65_LH_OAI22X6 U1194 ( .A(n131), .B(n6252), .C(n817), .D(n6256), .Z(n1911)
         );
  HS65_LH_OAI22X6 U1195 ( .A(n130), .B(n6252), .C(n816), .D(n6256), .Z(n1912)
         );
  HS65_LH_OAI22X6 U1196 ( .A(n129), .B(n6252), .C(n815), .D(n6256), .Z(n1913)
         );
  HS65_LH_OAI22X6 U1197 ( .A(n24), .B(n6323), .C(n838), .D(n6325), .Z(n2338)
         );
  HS65_LH_OAI22X6 U1198 ( .A(n23), .B(n6323), .C(n837), .D(n6325), .Z(n2339)
         );
  HS65_LH_OAI22X6 U1199 ( .A(n22), .B(n6323), .C(n836), .D(n6325), .Z(n2340)
         );
  HS65_LH_OAI22X6 U1200 ( .A(n21), .B(n6323), .C(n835), .D(n6325), .Z(n2341)
         );
  HS65_LH_OAI22X6 U1201 ( .A(n20), .B(n6323), .C(n834), .D(n6325), .Z(n2342)
         );
  HS65_LH_OAI22X6 U1202 ( .A(n19), .B(n6323), .C(n833), .D(n6325), .Z(n2343)
         );
  HS65_LH_OAI22X6 U1203 ( .A(n18), .B(n6323), .C(n832), .D(n6325), .Z(n2344)
         );
  HS65_LH_OAI22X6 U1204 ( .A(n17), .B(n6323), .C(n831), .D(n6325), .Z(n2345)
         );
  HS65_LH_OAI22X6 U1205 ( .A(n16), .B(n6323), .C(n830), .D(n6325), .Z(n2346)
         );
  HS65_LH_OAI22X6 U1206 ( .A(n15), .B(n6323), .C(n829), .D(n6325), .Z(n2347)
         );
  HS65_LH_OAI22X6 U1207 ( .A(n14), .B(n6323), .C(n828), .D(n6325), .Z(n2348)
         );
  HS65_LH_OAI22X6 U1208 ( .A(n13), .B(n6323), .C(n827), .D(n6325), .Z(n2349)
         );
  HS65_LH_OAI22X6 U1209 ( .A(n12), .B(n6322), .C(n826), .D(n6326), .Z(n2350)
         );
  HS65_LH_OAI22X6 U1210 ( .A(n11), .B(n6322), .C(n825), .D(n6326), .Z(n2351)
         );
  HS65_LH_OAI22X6 U1211 ( .A(n10), .B(n6322), .C(n824), .D(n6326), .Z(n2352)
         );
  HS65_LH_OAI22X6 U1212 ( .A(n9), .B(n6322), .C(n823), .D(n6326), .Z(n2353) );
  HS65_LH_OAI22X6 U1213 ( .A(n8), .B(n6322), .C(n822), .D(n6326), .Z(n2354) );
  HS65_LH_OAI22X6 U1214 ( .A(n7), .B(n6322), .C(n821), .D(n6326), .Z(n2355) );
  HS65_LH_OAI22X6 U1215 ( .A(n6), .B(n6322), .C(n820), .D(n6326), .Z(n2356) );
  HS65_LH_OAI22X6 U1216 ( .A(n5), .B(n6322), .C(n819), .D(n6326), .Z(n2357) );
  HS65_LH_OAI22X6 U1217 ( .A(n4), .B(n6322), .C(n818), .D(n6326), .Z(n2358) );
  HS65_LH_OAI22X6 U1218 ( .A(n3), .B(n6322), .C(n817), .D(n6326), .Z(n2359) );
  HS65_LH_OAI22X6 U1219 ( .A(n2), .B(n6322), .C(n816), .D(n6326), .Z(n2360) );
  HS65_LH_OAI22X6 U1220 ( .A(n1), .B(n6322), .C(n815), .D(n6326), .Z(n2361) );
  HS65_LH_OAI22X6 U1221 ( .A(n120), .B(n6308), .C(n838), .D(n6310), .Z(n2242)
         );
  HS65_LH_OAI22X6 U1222 ( .A(n119), .B(n6308), .C(n837), .D(n6310), .Z(n2243)
         );
  HS65_LH_OAI22X6 U1223 ( .A(n118), .B(n6308), .C(n836), .D(n6310), .Z(n2244)
         );
  HS65_LH_OAI22X6 U1224 ( .A(n117), .B(n6308), .C(n835), .D(n6310), .Z(n2245)
         );
  HS65_LH_OAI22X6 U1225 ( .A(n116), .B(n6308), .C(n834), .D(n6310), .Z(n2246)
         );
  HS65_LH_OAI22X6 U1226 ( .A(n115), .B(n6308), .C(n833), .D(n6310), .Z(n2247)
         );
  HS65_LH_OAI22X6 U1227 ( .A(n114), .B(n6308), .C(n832), .D(n6310), .Z(n2248)
         );
  HS65_LH_OAI22X6 U1228 ( .A(n113), .B(n6308), .C(n831), .D(n6310), .Z(n2249)
         );
  HS65_LH_OAI22X6 U1229 ( .A(n112), .B(n6308), .C(n830), .D(n6310), .Z(n2250)
         );
  HS65_LH_OAI22X6 U1230 ( .A(n111), .B(n6308), .C(n829), .D(n6310), .Z(n2251)
         );
  HS65_LH_OAI22X6 U1231 ( .A(n110), .B(n6308), .C(n828), .D(n6310), .Z(n2252)
         );
  HS65_LH_OAI22X6 U1232 ( .A(n109), .B(n6308), .C(n827), .D(n6310), .Z(n2253)
         );
  HS65_LH_OAI22X6 U1233 ( .A(n108), .B(n6307), .C(n826), .D(n6311), .Z(n2254)
         );
  HS65_LH_OAI22X6 U1234 ( .A(n107), .B(n6307), .C(n825), .D(n6311), .Z(n2255)
         );
  HS65_LH_OAI22X6 U1235 ( .A(n106), .B(n6307), .C(n824), .D(n6311), .Z(n2256)
         );
  HS65_LH_OAI22X6 U1236 ( .A(n105), .B(n6307), .C(n823), .D(n6311), .Z(n2257)
         );
  HS65_LH_OAI22X6 U1237 ( .A(n104), .B(n6307), .C(n822), .D(n6311), .Z(n2258)
         );
  HS65_LH_OAI22X6 U1238 ( .A(n103), .B(n6307), .C(n821), .D(n6311), .Z(n2259)
         );
  HS65_LH_OAI22X6 U1239 ( .A(n102), .B(n6307), .C(n820), .D(n6311), .Z(n2260)
         );
  HS65_LH_OAI22X6 U1240 ( .A(n101), .B(n6307), .C(n819), .D(n6311), .Z(n2261)
         );
  HS65_LH_OAI22X6 U1241 ( .A(n100), .B(n6307), .C(n818), .D(n6311), .Z(n2262)
         );
  HS65_LH_OAI22X6 U1242 ( .A(n99), .B(n6307), .C(n817), .D(n6311), .Z(n2263)
         );
  HS65_LH_OAI22X6 U1243 ( .A(n98), .B(n6307), .C(n816), .D(n6311), .Z(n2264)
         );
  HS65_LH_OAI22X6 U1244 ( .A(n97), .B(n6307), .C(n815), .D(n6311), .Z(n2265)
         );
  HS65_LH_OAI22X6 U1245 ( .A(n56), .B(n6318), .C(n838), .D(n6320), .Z(n2306)
         );
  HS65_LH_OAI22X6 U1246 ( .A(n55), .B(n6318), .C(n837), .D(n6320), .Z(n2307)
         );
  HS65_LH_OAI22X6 U1247 ( .A(n54), .B(n6318), .C(n836), .D(n6320), .Z(n2308)
         );
  HS65_LH_OAI22X6 U1248 ( .A(n53), .B(n6318), .C(n835), .D(n6320), .Z(n2309)
         );
  HS65_LH_OAI22X6 U1249 ( .A(n52), .B(n6318), .C(n834), .D(n6320), .Z(n2310)
         );
  HS65_LH_OAI22X6 U1250 ( .A(n51), .B(n6318), .C(n833), .D(n6320), .Z(n2311)
         );
  HS65_LH_OAI22X6 U1251 ( .A(n50), .B(n6318), .C(n832), .D(n6320), .Z(n2312)
         );
  HS65_LH_OAI22X6 U1252 ( .A(n49), .B(n6318), .C(n831), .D(n6320), .Z(n2313)
         );
  HS65_LH_OAI22X6 U1253 ( .A(n48), .B(n6318), .C(n830), .D(n6320), .Z(n2314)
         );
  HS65_LH_OAI22X6 U1254 ( .A(n47), .B(n6318), .C(n829), .D(n6320), .Z(n2315)
         );
  HS65_LH_OAI22X6 U1255 ( .A(n46), .B(n6318), .C(n828), .D(n6320), .Z(n2316)
         );
  HS65_LH_OAI22X6 U1256 ( .A(n45), .B(n6318), .C(n827), .D(n6320), .Z(n2317)
         );
  HS65_LH_OAI22X6 U1257 ( .A(n44), .B(n6317), .C(n826), .D(n6321), .Z(n2318)
         );
  HS65_LH_OAI22X6 U1258 ( .A(n43), .B(n6317), .C(n825), .D(n6321), .Z(n2319)
         );
  HS65_LH_OAI22X6 U1259 ( .A(n42), .B(n6317), .C(n824), .D(n6321), .Z(n2320)
         );
  HS65_LH_OAI22X6 U1260 ( .A(n41), .B(n6317), .C(n823), .D(n6321), .Z(n2321)
         );
  HS65_LH_OAI22X6 U1261 ( .A(n40), .B(n6317), .C(n822), .D(n6321), .Z(n2322)
         );
  HS65_LH_OAI22X6 U1262 ( .A(n39), .B(n6317), .C(n821), .D(n6321), .Z(n2323)
         );
  HS65_LH_OAI22X6 U1263 ( .A(n38), .B(n6317), .C(n820), .D(n6321), .Z(n2324)
         );
  HS65_LH_OAI22X6 U1264 ( .A(n37), .B(n6317), .C(n819), .D(n6321), .Z(n2325)
         );
  HS65_LH_OAI22X6 U1265 ( .A(n36), .B(n6317), .C(n818), .D(n6321), .Z(n2326)
         );
  HS65_LH_OAI22X6 U1266 ( .A(n35), .B(n6317), .C(n817), .D(n6321), .Z(n2327)
         );
  HS65_LH_OAI22X6 U1267 ( .A(n34), .B(n6317), .C(n816), .D(n6321), .Z(n2328)
         );
  HS65_LH_OAI22X6 U1268 ( .A(n33), .B(n6317), .C(n815), .D(n6321), .Z(n2329)
         );
  HS65_LH_OAI22X6 U1269 ( .A(n88), .B(n6313), .C(n838), .D(n6315), .Z(n2274)
         );
  HS65_LH_OAI22X6 U1270 ( .A(n87), .B(n6313), .C(n837), .D(n6315), .Z(n2275)
         );
  HS65_LH_OAI22X6 U1271 ( .A(n86), .B(n6313), .C(n836), .D(n6315), .Z(n2276)
         );
  HS65_LH_OAI22X6 U1272 ( .A(n85), .B(n6313), .C(n835), .D(n6315), .Z(n2277)
         );
  HS65_LH_OAI22X6 U1273 ( .A(n84), .B(n6313), .C(n834), .D(n6315), .Z(n2278)
         );
  HS65_LH_OAI22X6 U1274 ( .A(n83), .B(n6313), .C(n833), .D(n6315), .Z(n2279)
         );
  HS65_LH_OAI22X6 U1275 ( .A(n82), .B(n6313), .C(n832), .D(n6315), .Z(n2280)
         );
  HS65_LH_OAI22X6 U1276 ( .A(n81), .B(n6313), .C(n831), .D(n6315), .Z(n2281)
         );
  HS65_LH_OAI22X6 U1277 ( .A(n80), .B(n6313), .C(n830), .D(n6315), .Z(n2282)
         );
  HS65_LH_OAI22X6 U1278 ( .A(n79), .B(n6313), .C(n829), .D(n6315), .Z(n2283)
         );
  HS65_LH_OAI22X6 U1279 ( .A(n78), .B(n6313), .C(n828), .D(n6315), .Z(n2284)
         );
  HS65_LH_OAI22X6 U1280 ( .A(n77), .B(n6313), .C(n827), .D(n6315), .Z(n2285)
         );
  HS65_LH_OAI22X6 U1281 ( .A(n76), .B(n6312), .C(n826), .D(n6316), .Z(n2286)
         );
  HS65_LH_OAI22X6 U1282 ( .A(n75), .B(n6312), .C(n825), .D(n6316), .Z(n2287)
         );
  HS65_LH_OAI22X6 U1283 ( .A(n74), .B(n6312), .C(n824), .D(n6316), .Z(n2288)
         );
  HS65_LH_OAI22X6 U1284 ( .A(n73), .B(n6312), .C(n823), .D(n6316), .Z(n2289)
         );
  HS65_LH_OAI22X6 U1285 ( .A(n72), .B(n6312), .C(n822), .D(n6316), .Z(n2290)
         );
  HS65_LH_OAI22X6 U1286 ( .A(n71), .B(n6312), .C(n821), .D(n6316), .Z(n2291)
         );
  HS65_LH_OAI22X6 U1287 ( .A(n70), .B(n6312), .C(n820), .D(n6316), .Z(n2292)
         );
  HS65_LH_OAI22X6 U1288 ( .A(n69), .B(n6312), .C(n819), .D(n6316), .Z(n2293)
         );
  HS65_LH_OAI22X6 U1289 ( .A(n68), .B(n6312), .C(n818), .D(n6316), .Z(n2294)
         );
  HS65_LH_OAI22X6 U1290 ( .A(n67), .B(n6312), .C(n817), .D(n6316), .Z(n2295)
         );
  HS65_LH_OAI22X6 U1291 ( .A(n66), .B(n6312), .C(n816), .D(n6316), .Z(n2296)
         );
  HS65_LH_OAI22X6 U1292 ( .A(n65), .B(n6312), .C(n815), .D(n6316), .Z(n2297)
         );
  HS65_LH_OAI22X6 U1293 ( .A(n256), .B(n6218), .C(n846), .D(n6219), .Z(n1658)
         );
  HS65_LH_OAI22X6 U1294 ( .A(n255), .B(n6217), .C(n845), .D(n6220), .Z(n1659)
         );
  HS65_LH_OAI22X6 U1295 ( .A(n254), .B(n6218), .C(n844), .D(n6220), .Z(n1660)
         );
  HS65_LH_OAI22X6 U1296 ( .A(n253), .B(n6217), .C(n843), .D(n6220), .Z(n1661)
         );
  HS65_LH_OAI22X6 U1297 ( .A(n252), .B(n6218), .C(n842), .D(n6220), .Z(n1662)
         );
  HS65_LH_OAI22X6 U1298 ( .A(n251), .B(n6217), .C(n841), .D(n6220), .Z(n1663)
         );
  HS65_LH_OAI22X6 U1299 ( .A(n250), .B(n6218), .C(n840), .D(n6220), .Z(n1664)
         );
  HS65_LH_OAI22X6 U1300 ( .A(n249), .B(n6217), .C(n839), .D(n6220), .Z(n1665)
         );
  HS65_LH_OAI22X6 U1301 ( .A(n224), .B(n6223), .C(n846), .D(n6224), .Z(n1690)
         );
  HS65_LH_OAI22X6 U1302 ( .A(n223), .B(n6222), .C(n845), .D(n6225), .Z(n1691)
         );
  HS65_LH_OAI22X6 U1303 ( .A(n222), .B(n6223), .C(n844), .D(n6225), .Z(n1692)
         );
  HS65_LH_OAI22X6 U1304 ( .A(n221), .B(n6222), .C(n843), .D(n6225), .Z(n1693)
         );
  HS65_LH_OAI22X6 U1305 ( .A(n220), .B(n6223), .C(n842), .D(n6225), .Z(n1694)
         );
  HS65_LH_OAI22X6 U1306 ( .A(n219), .B(n6222), .C(n841), .D(n6225), .Z(n1695)
         );
  HS65_LH_OAI22X6 U1307 ( .A(n218), .B(n6223), .C(n840), .D(n6225), .Z(n1696)
         );
  HS65_LH_OAI22X6 U1308 ( .A(n217), .B(n6222), .C(n839), .D(n6225), .Z(n1697)
         );
  HS65_LH_OAI22X6 U1309 ( .A(n192), .B(n6248), .C(n846), .D(n6249), .Z(n1850)
         );
  HS65_LH_OAI22X6 U1310 ( .A(n191), .B(n6247), .C(n845), .D(n6250), .Z(n1851)
         );
  HS65_LH_OAI22X6 U1311 ( .A(n190), .B(n6248), .C(n844), .D(n6250), .Z(n1852)
         );
  HS65_LH_OAI22X6 U1312 ( .A(n189), .B(n6247), .C(n843), .D(n6250), .Z(n1853)
         );
  HS65_LH_OAI22X6 U1313 ( .A(n188), .B(n6248), .C(n842), .D(n6250), .Z(n1854)
         );
  HS65_LH_OAI22X6 U1314 ( .A(n187), .B(n6247), .C(n841), .D(n6250), .Z(n1855)
         );
  HS65_LH_OAI22X6 U1315 ( .A(n186), .B(n6248), .C(n840), .D(n6250), .Z(n1856)
         );
  HS65_LH_OAI22X6 U1316 ( .A(n185), .B(n6247), .C(n839), .D(n6250), .Z(n1857)
         );
  HS65_LH_OAI22X6 U1317 ( .A(n160), .B(n6253), .C(n846), .D(n6254), .Z(n1882)
         );
  HS65_LH_OAI22X6 U1318 ( .A(n159), .B(n6252), .C(n845), .D(n6255), .Z(n1883)
         );
  HS65_LH_OAI22X6 U1319 ( .A(n158), .B(n6253), .C(n844), .D(n6255), .Z(n1884)
         );
  HS65_LH_OAI22X6 U1320 ( .A(n157), .B(n6252), .C(n843), .D(n6255), .Z(n1885)
         );
  HS65_LH_OAI22X6 U1321 ( .A(n156), .B(n6253), .C(n842), .D(n6255), .Z(n1886)
         );
  HS65_LH_OAI22X6 U1322 ( .A(n155), .B(n6252), .C(n841), .D(n6255), .Z(n1887)
         );
  HS65_LH_OAI22X6 U1323 ( .A(n154), .B(n6253), .C(n840), .D(n6255), .Z(n1888)
         );
  HS65_LH_OAI22X6 U1324 ( .A(n153), .B(n6252), .C(n839), .D(n6255), .Z(n1889)
         );
  HS65_LH_OAI22X6 U1325 ( .A(n32), .B(n6323), .C(n846), .D(n6324), .Z(n2330)
         );
  HS65_LH_OAI22X6 U1326 ( .A(n31), .B(n6322), .C(n845), .D(n6325), .Z(n2331)
         );
  HS65_LH_OAI22X6 U1327 ( .A(n30), .B(n6323), .C(n844), .D(n6325), .Z(n2332)
         );
  HS65_LH_OAI22X6 U1328 ( .A(n29), .B(n6322), .C(n843), .D(n6325), .Z(n2333)
         );
  HS65_LH_OAI22X6 U1329 ( .A(n28), .B(n6323), .C(n842), .D(n6325), .Z(n2334)
         );
  HS65_LH_OAI22X6 U1330 ( .A(n27), .B(n6322), .C(n841), .D(n6325), .Z(n2335)
         );
  HS65_LH_OAI22X6 U1331 ( .A(n26), .B(n6323), .C(n840), .D(n6325), .Z(n2336)
         );
  HS65_LH_OAI22X6 U1332 ( .A(n25), .B(n6322), .C(n839), .D(n6325), .Z(n2337)
         );
  HS65_LH_OAI22X6 U1333 ( .A(n128), .B(n6308), .C(n846), .D(n6309), .Z(n2234)
         );
  HS65_LH_OAI22X6 U1334 ( .A(n127), .B(n6307), .C(n845), .D(n6310), .Z(n2235)
         );
  HS65_LH_OAI22X6 U1335 ( .A(n126), .B(n6308), .C(n844), .D(n6310), .Z(n2236)
         );
  HS65_LH_OAI22X6 U1336 ( .A(n125), .B(n6307), .C(n843), .D(n6310), .Z(n2237)
         );
  HS65_LH_OAI22X6 U1337 ( .A(n124), .B(n6308), .C(n842), .D(n6310), .Z(n2238)
         );
  HS65_LH_OAI22X6 U1338 ( .A(n123), .B(n6307), .C(n841), .D(n6310), .Z(n2239)
         );
  HS65_LH_OAI22X6 U1339 ( .A(n122), .B(n6308), .C(n840), .D(n6310), .Z(n2240)
         );
  HS65_LH_OAI22X6 U1340 ( .A(n121), .B(n6307), .C(n839), .D(n6310), .Z(n2241)
         );
  HS65_LH_OAI22X6 U1341 ( .A(n64), .B(n6318), .C(n846), .D(n6319), .Z(n2298)
         );
  HS65_LH_OAI22X6 U1342 ( .A(n63), .B(n6317), .C(n845), .D(n6320), .Z(n2299)
         );
  HS65_LH_OAI22X6 U1343 ( .A(n62), .B(n6318), .C(n844), .D(n6320), .Z(n2300)
         );
  HS65_LH_OAI22X6 U1344 ( .A(n61), .B(n6317), .C(n843), .D(n6320), .Z(n2301)
         );
  HS65_LH_OAI22X6 U1345 ( .A(n60), .B(n6318), .C(n842), .D(n6320), .Z(n2302)
         );
  HS65_LH_OAI22X6 U1346 ( .A(n59), .B(n6317), .C(n841), .D(n6320), .Z(n2303)
         );
  HS65_LH_OAI22X6 U1347 ( .A(n58), .B(n6318), .C(n840), .D(n6320), .Z(n2304)
         );
  HS65_LH_OAI22X6 U1348 ( .A(n57), .B(n6317), .C(n839), .D(n6320), .Z(n2305)
         );
  HS65_LH_OAI22X6 U1349 ( .A(n96), .B(n6313), .C(n846), .D(n6314), .Z(n2266)
         );
  HS65_LH_OAI22X6 U1350 ( .A(n95), .B(n6312), .C(n845), .D(n6315), .Z(n2267)
         );
  HS65_LH_OAI22X6 U1351 ( .A(n94), .B(n6313), .C(n844), .D(n6315), .Z(n2268)
         );
  HS65_LH_OAI22X6 U1352 ( .A(n93), .B(n6312), .C(n843), .D(n6315), .Z(n2269)
         );
  HS65_LH_OAI22X6 U1353 ( .A(n92), .B(n6313), .C(n842), .D(n6315), .Z(n2270)
         );
  HS65_LH_OAI22X6 U1354 ( .A(n91), .B(n6312), .C(n841), .D(n6315), .Z(n2271)
         );
  HS65_LH_OAI22X6 U1355 ( .A(n90), .B(n6313), .C(n840), .D(n6315), .Z(n2272)
         );
  HS65_LH_OAI22X6 U1356 ( .A(n89), .B(n6312), .C(n839), .D(n6315), .Z(n2273)
         );
  HS65_LH_IVX9 U1357 ( .A(\registers[25][0] ), .Z(n288) );
  HS65_LH_IVX9 U1358 ( .A(\registers[25][1] ), .Z(n287) );
  HS65_LH_IVX9 U1359 ( .A(\registers[25][2] ), .Z(n286) );
  HS65_LH_IVX9 U1360 ( .A(\registers[25][3] ), .Z(n285) );
  HS65_LH_IVX9 U1361 ( .A(\registers[25][4] ), .Z(n284) );
  HS65_LH_IVX9 U1362 ( .A(\registers[25][5] ), .Z(n283) );
  HS65_LH_IVX9 U1363 ( .A(\registers[25][6] ), .Z(n282) );
  HS65_LH_IVX9 U1364 ( .A(\registers[25][7] ), .Z(n281) );
  HS65_LH_IVX9 U1365 ( .A(\registers[25][8] ), .Z(n280) );
  HS65_LH_IVX9 U1366 ( .A(\registers[25][9] ), .Z(n279) );
  HS65_LH_IVX9 U1367 ( .A(\registers[25][10] ), .Z(n278) );
  HS65_LH_IVX9 U1368 ( .A(\registers[25][11] ), .Z(n277) );
  HS65_LH_IVX9 U1369 ( .A(\registers[25][12] ), .Z(n276) );
  HS65_LH_IVX9 U1370 ( .A(\registers[25][13] ), .Z(n275) );
  HS65_LH_IVX9 U1371 ( .A(\registers[25][14] ), .Z(n274) );
  HS65_LH_IVX9 U1372 ( .A(\registers[25][15] ), .Z(n273) );
  HS65_LH_IVX9 U1373 ( .A(\registers[25][16] ), .Z(n272) );
  HS65_LH_IVX9 U1374 ( .A(\registers[25][17] ), .Z(n271) );
  HS65_LH_IVX9 U1375 ( .A(\registers[25][18] ), .Z(n270) );
  HS65_LH_IVX9 U1376 ( .A(\registers[25][19] ), .Z(n269) );
  HS65_LH_IVX9 U1377 ( .A(\registers[25][20] ), .Z(n268) );
  HS65_LH_IVX9 U1378 ( .A(\registers[25][21] ), .Z(n267) );
  HS65_LH_IVX9 U1379 ( .A(\registers[25][22] ), .Z(n266) );
  HS65_LH_IVX9 U1380 ( .A(\registers[25][23] ), .Z(n265) );
  HS65_LH_IVX9 U1381 ( .A(\registers[25][24] ), .Z(n264) );
  HS65_LH_IVX9 U1382 ( .A(\registers[25][25] ), .Z(n263) );
  HS65_LH_IVX9 U1383 ( .A(\registers[25][26] ), .Z(n262) );
  HS65_LH_IVX9 U1384 ( .A(\registers[25][27] ), .Z(n261) );
  HS65_LH_IVX9 U1385 ( .A(\registers[25][28] ), .Z(n260) );
  HS65_LH_IVX9 U1386 ( .A(\registers[25][29] ), .Z(n259) );
  HS65_LH_IVX9 U1387 ( .A(\registers[25][30] ), .Z(n258) );
  HS65_LH_IVX9 U1388 ( .A(\registers[25][31] ), .Z(n257) );
  HS65_LH_IVX9 U1389 ( .A(\registers[16][0] ), .Z(n416) );
  HS65_LH_IVX9 U1390 ( .A(\registers[16][1] ), .Z(n415) );
  HS65_LH_IVX9 U1391 ( .A(\registers[16][2] ), .Z(n414) );
  HS65_LH_IVX9 U1392 ( .A(\registers[16][3] ), .Z(n413) );
  HS65_LH_IVX9 U1393 ( .A(\registers[16][4] ), .Z(n412) );
  HS65_LH_IVX9 U1394 ( .A(\registers[16][5] ), .Z(n411) );
  HS65_LH_IVX9 U1395 ( .A(\registers[16][6] ), .Z(n410) );
  HS65_LH_IVX9 U1396 ( .A(\registers[16][7] ), .Z(n409) );
  HS65_LH_IVX9 U1397 ( .A(\registers[16][8] ), .Z(n408) );
  HS65_LH_IVX9 U1398 ( .A(\registers[16][9] ), .Z(n407) );
  HS65_LH_IVX9 U1399 ( .A(\registers[16][10] ), .Z(n406) );
  HS65_LH_IVX9 U1400 ( .A(\registers[16][11] ), .Z(n405) );
  HS65_LH_IVX9 U1401 ( .A(\registers[16][12] ), .Z(n404) );
  HS65_LH_IVX9 U1402 ( .A(\registers[16][13] ), .Z(n403) );
  HS65_LH_IVX9 U1403 ( .A(\registers[16][14] ), .Z(n402) );
  HS65_LH_IVX9 U1404 ( .A(\registers[16][15] ), .Z(n401) );
  HS65_LH_IVX9 U1405 ( .A(\registers[16][16] ), .Z(n400) );
  HS65_LH_IVX9 U1406 ( .A(\registers[16][17] ), .Z(n399) );
  HS65_LH_IVX9 U1407 ( .A(\registers[16][18] ), .Z(n398) );
  HS65_LH_IVX9 U1408 ( .A(\registers[16][19] ), .Z(n397) );
  HS65_LH_IVX9 U1409 ( .A(\registers[16][20] ), .Z(n396) );
  HS65_LH_IVX9 U1410 ( .A(\registers[16][21] ), .Z(n395) );
  HS65_LH_IVX9 U1411 ( .A(\registers[16][22] ), .Z(n394) );
  HS65_LH_IVX9 U1412 ( .A(\registers[16][23] ), .Z(n393) );
  HS65_LH_IVX9 U1413 ( .A(\registers[16][24] ), .Z(n392) );
  HS65_LH_IVX9 U1414 ( .A(\registers[16][25] ), .Z(n391) );
  HS65_LH_IVX9 U1415 ( .A(\registers[16][26] ), .Z(n390) );
  HS65_LH_IVX9 U1416 ( .A(\registers[16][27] ), .Z(n389) );
  HS65_LH_IVX9 U1417 ( .A(\registers[16][28] ), .Z(n388) );
  HS65_LH_IVX9 U1418 ( .A(\registers[16][29] ), .Z(n387) );
  HS65_LH_IVX9 U1419 ( .A(\registers[16][30] ), .Z(n386) );
  HS65_LH_IVX9 U1420 ( .A(\registers[16][31] ), .Z(n385) );
  HS65_LH_IVX9 U1421 ( .A(\registers[10][0] ), .Z(n480) );
  HS65_LH_IVX9 U1422 ( .A(\registers[10][1] ), .Z(n479) );
  HS65_LH_IVX9 U1423 ( .A(\registers[10][2] ), .Z(n478) );
  HS65_LH_IVX9 U1424 ( .A(\registers[10][3] ), .Z(n477) );
  HS65_LH_IVX9 U1425 ( .A(\registers[10][4] ), .Z(n476) );
  HS65_LH_IVX9 U1426 ( .A(\registers[10][5] ), .Z(n475) );
  HS65_LH_IVX9 U1427 ( .A(\registers[10][6] ), .Z(n474) );
  HS65_LH_IVX9 U1428 ( .A(\registers[10][7] ), .Z(n473) );
  HS65_LH_IVX9 U1429 ( .A(\registers[10][8] ), .Z(n472) );
  HS65_LH_IVX9 U1430 ( .A(\registers[10][9] ), .Z(n471) );
  HS65_LH_IVX9 U1431 ( .A(\registers[10][10] ), .Z(n470) );
  HS65_LH_IVX9 U1432 ( .A(\registers[10][11] ), .Z(n469) );
  HS65_LH_IVX9 U1433 ( .A(\registers[10][12] ), .Z(n468) );
  HS65_LH_IVX9 U1434 ( .A(\registers[10][13] ), .Z(n467) );
  HS65_LH_IVX9 U1435 ( .A(\registers[10][14] ), .Z(n466) );
  HS65_LH_IVX9 U1436 ( .A(\registers[10][15] ), .Z(n465) );
  HS65_LH_IVX9 U1437 ( .A(\registers[10][16] ), .Z(n464) );
  HS65_LH_IVX9 U1438 ( .A(\registers[10][17] ), .Z(n463) );
  HS65_LH_IVX9 U1439 ( .A(\registers[10][18] ), .Z(n462) );
  HS65_LH_IVX9 U1440 ( .A(\registers[10][19] ), .Z(n461) );
  HS65_LH_IVX9 U1441 ( .A(\registers[10][20] ), .Z(n460) );
  HS65_LH_IVX9 U1442 ( .A(\registers[10][21] ), .Z(n459) );
  HS65_LH_IVX9 U1443 ( .A(\registers[10][22] ), .Z(n458) );
  HS65_LH_IVX9 U1444 ( .A(\registers[10][23] ), .Z(n457) );
  HS65_LH_IVX9 U1445 ( .A(\registers[10][24] ), .Z(n456) );
  HS65_LH_IVX9 U1446 ( .A(\registers[10][25] ), .Z(n455) );
  HS65_LH_IVX9 U1447 ( .A(\registers[10][26] ), .Z(n454) );
  HS65_LH_IVX9 U1448 ( .A(\registers[10][27] ), .Z(n453) );
  HS65_LH_IVX9 U1449 ( .A(\registers[10][28] ), .Z(n452) );
  HS65_LH_IVX9 U1450 ( .A(\registers[10][29] ), .Z(n451) );
  HS65_LH_IVX9 U1451 ( .A(\registers[10][30] ), .Z(n450) );
  HS65_LH_IVX9 U1452 ( .A(\registers[10][31] ), .Z(n449) );
  HS65_LH_IVX9 U1453 ( .A(\registers[18][0] ), .Z(n352) );
  HS65_LH_IVX9 U1454 ( .A(\registers[18][1] ), .Z(n351) );
  HS65_LH_IVX9 U1455 ( .A(\registers[18][2] ), .Z(n350) );
  HS65_LH_IVX9 U1456 ( .A(\registers[18][3] ), .Z(n349) );
  HS65_LH_IVX9 U1457 ( .A(\registers[18][4] ), .Z(n348) );
  HS65_LH_IVX9 U1458 ( .A(\registers[18][5] ), .Z(n347) );
  HS65_LH_IVX9 U1459 ( .A(\registers[18][6] ), .Z(n346) );
  HS65_LH_IVX9 U1460 ( .A(\registers[18][7] ), .Z(n345) );
  HS65_LH_IVX9 U1461 ( .A(\registers[18][8] ), .Z(n344) );
  HS65_LH_IVX9 U1462 ( .A(\registers[18][9] ), .Z(n343) );
  HS65_LH_IVX9 U1463 ( .A(\registers[18][10] ), .Z(n342) );
  HS65_LH_IVX9 U1464 ( .A(\registers[18][11] ), .Z(n341) );
  HS65_LH_IVX9 U1465 ( .A(\registers[18][12] ), .Z(n340) );
  HS65_LH_IVX9 U1466 ( .A(\registers[18][13] ), .Z(n339) );
  HS65_LH_IVX9 U1467 ( .A(\registers[18][14] ), .Z(n338) );
  HS65_LH_IVX9 U1468 ( .A(\registers[18][15] ), .Z(n337) );
  HS65_LH_IVX9 U1469 ( .A(\registers[18][16] ), .Z(n336) );
  HS65_LH_IVX9 U1470 ( .A(\registers[18][17] ), .Z(n335) );
  HS65_LH_IVX9 U1471 ( .A(\registers[18][18] ), .Z(n334) );
  HS65_LH_IVX9 U1472 ( .A(\registers[18][19] ), .Z(n333) );
  HS65_LH_IVX9 U1473 ( .A(\registers[18][20] ), .Z(n332) );
  HS65_LH_IVX9 U1474 ( .A(\registers[18][21] ), .Z(n331) );
  HS65_LH_IVX9 U1475 ( .A(\registers[18][22] ), .Z(n330) );
  HS65_LH_IVX9 U1476 ( .A(\registers[18][23] ), .Z(n329) );
  HS65_LH_IVX9 U1477 ( .A(\registers[18][24] ), .Z(n328) );
  HS65_LH_IVX9 U1478 ( .A(\registers[18][25] ), .Z(n327) );
  HS65_LH_IVX9 U1479 ( .A(\registers[18][26] ), .Z(n326) );
  HS65_LH_IVX9 U1480 ( .A(\registers[18][27] ), .Z(n325) );
  HS65_LH_IVX9 U1481 ( .A(\registers[18][28] ), .Z(n324) );
  HS65_LH_IVX9 U1482 ( .A(\registers[18][29] ), .Z(n323) );
  HS65_LH_IVX9 U1483 ( .A(\registers[18][30] ), .Z(n322) );
  HS65_LH_IVX9 U1484 ( .A(\registers[18][31] ), .Z(n321) );
  HS65_LH_IVX9 U1485 ( .A(\registers[24][0] ), .Z(n320) );
  HS65_LH_IVX9 U1486 ( .A(\registers[24][1] ), .Z(n319) );
  HS65_LH_IVX9 U1487 ( .A(\registers[24][2] ), .Z(n318) );
  HS65_LH_IVX9 U1488 ( .A(\registers[24][3] ), .Z(n317) );
  HS65_LH_IVX9 U1489 ( .A(\registers[24][4] ), .Z(n316) );
  HS65_LH_IVX9 U1490 ( .A(\registers[24][5] ), .Z(n315) );
  HS65_LH_IVX9 U1491 ( .A(\registers[24][6] ), .Z(n314) );
  HS65_LH_IVX9 U1492 ( .A(\registers[24][7] ), .Z(n313) );
  HS65_LH_IVX9 U1493 ( .A(\registers[24][8] ), .Z(n312) );
  HS65_LH_IVX9 U1494 ( .A(\registers[24][9] ), .Z(n311) );
  HS65_LH_IVX9 U1495 ( .A(\registers[24][10] ), .Z(n310) );
  HS65_LH_IVX9 U1496 ( .A(\registers[24][11] ), .Z(n309) );
  HS65_LH_IVX9 U1497 ( .A(\registers[24][12] ), .Z(n308) );
  HS65_LH_IVX9 U1498 ( .A(\registers[24][13] ), .Z(n307) );
  HS65_LH_IVX9 U1499 ( .A(\registers[24][14] ), .Z(n306) );
  HS65_LH_IVX9 U1500 ( .A(\registers[24][15] ), .Z(n305) );
  HS65_LH_IVX9 U1501 ( .A(\registers[24][16] ), .Z(n304) );
  HS65_LH_IVX9 U1502 ( .A(\registers[24][17] ), .Z(n303) );
  HS65_LH_IVX9 U1503 ( .A(\registers[24][18] ), .Z(n302) );
  HS65_LH_IVX9 U1504 ( .A(\registers[24][19] ), .Z(n301) );
  HS65_LH_IVX9 U1505 ( .A(\registers[24][20] ), .Z(n300) );
  HS65_LH_IVX9 U1506 ( .A(\registers[24][21] ), .Z(n299) );
  HS65_LH_IVX9 U1507 ( .A(\registers[24][22] ), .Z(n298) );
  HS65_LH_IVX9 U1508 ( .A(\registers[24][23] ), .Z(n297) );
  HS65_LH_IVX9 U1509 ( .A(\registers[24][24] ), .Z(n296) );
  HS65_LH_IVX9 U1510 ( .A(\registers[24][25] ), .Z(n295) );
  HS65_LH_IVX9 U1511 ( .A(\registers[24][26] ), .Z(n294) );
  HS65_LH_IVX9 U1512 ( .A(\registers[24][27] ), .Z(n293) );
  HS65_LH_IVX9 U1513 ( .A(\registers[24][28] ), .Z(n292) );
  HS65_LH_IVX9 U1514 ( .A(\registers[24][29] ), .Z(n291) );
  HS65_LH_IVX9 U1515 ( .A(\registers[24][30] ), .Z(n290) );
  HS65_LH_IVX9 U1516 ( .A(\registers[24][31] ), .Z(n289) );
  HS65_LH_IVX9 U1517 ( .A(\registers[6][0] ), .Z(n512) );
  HS65_LH_IVX9 U1518 ( .A(\registers[6][1] ), .Z(n511) );
  HS65_LH_IVX9 U1519 ( .A(\registers[6][2] ), .Z(n510) );
  HS65_LH_IVX9 U1520 ( .A(\registers[6][3] ), .Z(n509) );
  HS65_LH_IVX9 U1521 ( .A(\registers[6][4] ), .Z(n508) );
  HS65_LH_IVX9 U1522 ( .A(\registers[6][5] ), .Z(n507) );
  HS65_LH_IVX9 U1523 ( .A(\registers[6][6] ), .Z(n506) );
  HS65_LH_IVX9 U1524 ( .A(\registers[6][7] ), .Z(n505) );
  HS65_LH_IVX9 U1525 ( .A(\registers[6][8] ), .Z(n504) );
  HS65_LH_IVX9 U1526 ( .A(\registers[6][9] ), .Z(n503) );
  HS65_LH_IVX9 U1527 ( .A(\registers[6][10] ), .Z(n502) );
  HS65_LH_IVX9 U1528 ( .A(\registers[6][11] ), .Z(n501) );
  HS65_LH_IVX9 U1529 ( .A(\registers[6][12] ), .Z(n500) );
  HS65_LH_IVX9 U1530 ( .A(\registers[6][13] ), .Z(n499) );
  HS65_LH_IVX9 U1531 ( .A(\registers[6][14] ), .Z(n498) );
  HS65_LH_IVX9 U1532 ( .A(\registers[6][15] ), .Z(n497) );
  HS65_LH_IVX9 U1533 ( .A(\registers[6][16] ), .Z(n496) );
  HS65_LH_IVX9 U1534 ( .A(\registers[6][17] ), .Z(n495) );
  HS65_LH_IVX9 U1535 ( .A(\registers[6][18] ), .Z(n494) );
  HS65_LH_IVX9 U1536 ( .A(\registers[6][19] ), .Z(n493) );
  HS65_LH_IVX9 U1537 ( .A(\registers[6][20] ), .Z(n492) );
  HS65_LH_IVX9 U1538 ( .A(\registers[6][21] ), .Z(n491) );
  HS65_LH_IVX9 U1539 ( .A(\registers[6][22] ), .Z(n490) );
  HS65_LH_IVX9 U1540 ( .A(\registers[6][23] ), .Z(n489) );
  HS65_LH_IVX9 U1541 ( .A(\registers[6][24] ), .Z(n488) );
  HS65_LH_IVX9 U1542 ( .A(\registers[6][25] ), .Z(n487) );
  HS65_LH_IVX9 U1543 ( .A(\registers[6][26] ), .Z(n486) );
  HS65_LH_IVX9 U1544 ( .A(\registers[6][27] ), .Z(n485) );
  HS65_LH_IVX9 U1545 ( .A(\registers[6][28] ), .Z(n484) );
  HS65_LH_IVX9 U1546 ( .A(\registers[6][29] ), .Z(n483) );
  HS65_LH_IVX9 U1547 ( .A(\registers[6][30] ), .Z(n482) );
  HS65_LH_IVX9 U1548 ( .A(\registers[6][31] ), .Z(n481) );
  HS65_LH_IVX9 U1549 ( .A(\registers[17][0] ), .Z(n384) );
  HS65_LH_IVX9 U1550 ( .A(\registers[17][1] ), .Z(n383) );
  HS65_LH_IVX9 U1551 ( .A(\registers[17][2] ), .Z(n382) );
  HS65_LH_IVX9 U1552 ( .A(\registers[17][3] ), .Z(n381) );
  HS65_LH_IVX9 U1553 ( .A(\registers[17][4] ), .Z(n380) );
  HS65_LH_IVX9 U1554 ( .A(\registers[17][5] ), .Z(n379) );
  HS65_LH_IVX9 U1555 ( .A(\registers[17][6] ), .Z(n378) );
  HS65_LH_IVX9 U1556 ( .A(\registers[17][7] ), .Z(n377) );
  HS65_LH_IVX9 U1557 ( .A(\registers[17][8] ), .Z(n376) );
  HS65_LH_IVX9 U1558 ( .A(\registers[17][9] ), .Z(n375) );
  HS65_LH_IVX9 U1559 ( .A(\registers[17][10] ), .Z(n374) );
  HS65_LH_IVX9 U1560 ( .A(\registers[17][11] ), .Z(n373) );
  HS65_LH_IVX9 U1561 ( .A(\registers[17][12] ), .Z(n372) );
  HS65_LH_IVX9 U1562 ( .A(\registers[17][13] ), .Z(n371) );
  HS65_LH_IVX9 U1563 ( .A(\registers[17][14] ), .Z(n370) );
  HS65_LH_IVX9 U1564 ( .A(\registers[17][15] ), .Z(n369) );
  HS65_LH_IVX9 U1565 ( .A(\registers[17][16] ), .Z(n368) );
  HS65_LH_IVX9 U1566 ( .A(\registers[17][17] ), .Z(n367) );
  HS65_LH_IVX9 U1567 ( .A(\registers[17][18] ), .Z(n366) );
  HS65_LH_IVX9 U1568 ( .A(\registers[17][19] ), .Z(n365) );
  HS65_LH_IVX9 U1569 ( .A(\registers[17][20] ), .Z(n364) );
  HS65_LH_IVX9 U1570 ( .A(\registers[17][21] ), .Z(n363) );
  HS65_LH_IVX9 U1571 ( .A(\registers[17][22] ), .Z(n362) );
  HS65_LH_IVX9 U1572 ( .A(\registers[17][23] ), .Z(n361) );
  HS65_LH_IVX9 U1573 ( .A(\registers[17][24] ), .Z(n360) );
  HS65_LH_IVX9 U1574 ( .A(\registers[17][25] ), .Z(n359) );
  HS65_LH_IVX9 U1575 ( .A(\registers[17][26] ), .Z(n358) );
  HS65_LH_IVX9 U1576 ( .A(\registers[17][27] ), .Z(n357) );
  HS65_LH_IVX9 U1577 ( .A(\registers[17][28] ), .Z(n356) );
  HS65_LH_IVX9 U1578 ( .A(\registers[17][29] ), .Z(n355) );
  HS65_LH_IVX9 U1579 ( .A(\registers[17][30] ), .Z(n354) );
  HS65_LH_IVX9 U1580 ( .A(\registers[17][31] ), .Z(n353) );
  HS65_LH_IVX9 U1581 ( .A(\registers[12][0] ), .Z(n448) );
  HS65_LH_IVX9 U1582 ( .A(\registers[12][1] ), .Z(n447) );
  HS65_LH_IVX9 U1583 ( .A(\registers[12][2] ), .Z(n446) );
  HS65_LH_IVX9 U1584 ( .A(\registers[12][3] ), .Z(n445) );
  HS65_LH_IVX9 U1585 ( .A(\registers[12][4] ), .Z(n444) );
  HS65_LH_IVX9 U1586 ( .A(\registers[12][5] ), .Z(n443) );
  HS65_LH_IVX9 U1587 ( .A(\registers[12][6] ), .Z(n442) );
  HS65_LH_IVX9 U1588 ( .A(\registers[12][7] ), .Z(n441) );
  HS65_LH_IVX9 U1589 ( .A(\registers[12][8] ), .Z(n440) );
  HS65_LH_IVX9 U1590 ( .A(\registers[12][9] ), .Z(n439) );
  HS65_LH_IVX9 U1591 ( .A(\registers[12][10] ), .Z(n438) );
  HS65_LH_IVX9 U1592 ( .A(\registers[12][11] ), .Z(n437) );
  HS65_LH_IVX9 U1593 ( .A(\registers[12][12] ), .Z(n436) );
  HS65_LH_IVX9 U1594 ( .A(\registers[12][13] ), .Z(n435) );
  HS65_LH_IVX9 U1595 ( .A(\registers[12][14] ), .Z(n434) );
  HS65_LH_IVX9 U1596 ( .A(\registers[12][15] ), .Z(n433) );
  HS65_LH_IVX9 U1597 ( .A(\registers[12][16] ), .Z(n432) );
  HS65_LH_IVX9 U1598 ( .A(\registers[12][17] ), .Z(n431) );
  HS65_LH_IVX9 U1599 ( .A(\registers[12][18] ), .Z(n430) );
  HS65_LH_IVX9 U1600 ( .A(\registers[12][19] ), .Z(n429) );
  HS65_LH_IVX9 U1601 ( .A(\registers[12][20] ), .Z(n428) );
  HS65_LH_IVX9 U1602 ( .A(\registers[12][21] ), .Z(n427) );
  HS65_LH_IVX9 U1603 ( .A(\registers[12][22] ), .Z(n426) );
  HS65_LH_IVX9 U1604 ( .A(\registers[12][23] ), .Z(n425) );
  HS65_LH_IVX9 U1605 ( .A(\registers[12][24] ), .Z(n424) );
  HS65_LH_IVX9 U1606 ( .A(\registers[12][25] ), .Z(n423) );
  HS65_LH_IVX9 U1607 ( .A(\registers[12][26] ), .Z(n422) );
  HS65_LH_IVX9 U1608 ( .A(\registers[12][27] ), .Z(n421) );
  HS65_LH_IVX9 U1609 ( .A(\registers[12][28] ), .Z(n420) );
  HS65_LH_IVX9 U1610 ( .A(\registers[12][29] ), .Z(n419) );
  HS65_LH_IVX9 U1611 ( .A(\registers[12][30] ), .Z(n418) );
  HS65_LH_IVX9 U1612 ( .A(\registers[12][31] ), .Z(n417) );
  HS65_LH_AO22X9 U1613 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6246), .C(n6242), 
        .D(\registers[13][0] ), .Z(n1818) );
  HS65_LH_AO22X9 U1614 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6246), .C(n6242), 
        .D(\registers[13][1] ), .Z(n1819) );
  HS65_LH_AO22X9 U1615 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6246), .C(n6242), 
        .D(\registers[13][2] ), .Z(n1820) );
  HS65_LH_AO22X9 U1616 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6246), .C(n6242), 
        .D(\registers[13][3] ), .Z(n1821) );
  HS65_LH_AO22X9 U1617 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6246), .C(n6242), 
        .D(\registers[13][4] ), .Z(n1822) );
  HS65_LH_AO22X9 U1618 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6246), .C(n6242), 
        .D(\registers[13][5] ), .Z(n1823) );
  HS65_LH_AO22X9 U1619 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6246), .C(n6242), 
        .D(\registers[13][6] ), .Z(n1824) );
  HS65_LH_AO22X9 U1620 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6246), .C(n6242), 
        .D(\registers[13][7] ), .Z(n1825) );
  HS65_LH_AO22X9 U1621 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6246), .C(n6242), 
        .D(\registers[13][8] ), .Z(n1826) );
  HS65_LH_AO22X9 U1622 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6246), .C(n6242), 
        .D(\registers[13][9] ), .Z(n1827) );
  HS65_LH_AO22X9 U1623 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6246), .C(n6242), 
        .D(\registers[13][10] ), .Z(n1828) );
  HS65_LH_AO22X9 U1624 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6245), .C(n6242), 
        .D(\registers[13][11] ), .Z(n1829) );
  HS65_LH_AO22X9 U1625 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6245), .C(n6242), 
        .D(\registers[13][12] ), .Z(n1830) );
  HS65_LH_AO22X9 U1626 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6245), .C(n6243), 
        .D(\registers[13][13] ), .Z(n1831) );
  HS65_LH_AO22X9 U1627 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6245), .C(n6243), 
        .D(\registers[13][14] ), .Z(n1832) );
  HS65_LH_AO22X9 U1628 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6245), .C(n6243), 
        .D(\registers[13][15] ), .Z(n1833) );
  HS65_LH_AO22X9 U1629 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6245), .C(n6243), 
        .D(\registers[13][16] ), .Z(n1834) );
  HS65_LH_AO22X9 U1630 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6245), .C(n6243), 
        .D(\registers[13][17] ), .Z(n1835) );
  HS65_LH_AO22X9 U1631 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6245), .C(n6243), 
        .D(\registers[13][18] ), .Z(n1836) );
  HS65_LH_AO22X9 U1632 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6245), .C(n6243), 
        .D(\registers[13][19] ), .Z(n1837) );
  HS65_LH_AO22X9 U1633 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6245), .C(n6243), 
        .D(\registers[13][20] ), .Z(n1838) );
  HS65_LH_AO22X9 U1634 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6245), .C(n6243), 
        .D(\registers[13][21] ), .Z(n1839) );
  HS65_LH_AO22X9 U1635 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6245), .C(n6243), 
        .D(\registers[13][22] ), .Z(n1840) );
  HS65_LH_AO22X9 U1636 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6245), .C(n6243), 
        .D(\registers[13][23] ), .Z(n1841) );
  HS65_LH_AO22X9 U1637 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6245), .C(n6243), 
        .D(\registers[13][24] ), .Z(n1842) );
  HS65_LH_AO22X9 U1638 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6245), .C(n6243), 
        .D(\registers[13][25] ), .Z(n1843) );
  HS65_LH_AO22X9 U1639 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6245), .C(n6242), 
        .D(\registers[13][26] ), .Z(n1844) );
  HS65_LH_AO22X9 U1640 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6245), .C(n6243), 
        .D(\registers[13][27] ), .Z(n1845) );
  HS65_LH_AO22X9 U1641 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6245), .C(n6242), 
        .D(\registers[13][28] ), .Z(n1846) );
  HS65_LH_AO22X9 U1642 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6245), .C(n6243), 
        .D(\registers[13][29] ), .Z(n1847) );
  HS65_LH_AO22X9 U1643 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6245), .C(n6242), 
        .D(\registers[13][30] ), .Z(n1848) );
  HS65_LH_AO22X9 U1644 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6244), .C(n6243), 
        .D(\registers[13][31] ), .Z(n1849) );
  HS65_LH_AO22X9 U1645 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6201), .C(n6197), 
        .D(\registers[4][0] ), .Z(n1530) );
  HS65_LH_AO22X9 U1646 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6201), .C(n6197), 
        .D(\registers[4][1] ), .Z(n1531) );
  HS65_LH_AO22X9 U1647 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6201), .C(n6197), 
        .D(\registers[4][2] ), .Z(n1532) );
  HS65_LH_AO22X9 U1648 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6201), .C(n6197), 
        .D(\registers[4][3] ), .Z(n1533) );
  HS65_LH_AO22X9 U1649 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6201), .C(n6197), 
        .D(\registers[4][4] ), .Z(n1534) );
  HS65_LH_AO22X9 U1650 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6201), .C(n6197), 
        .D(\registers[4][5] ), .Z(n1535) );
  HS65_LH_AO22X9 U1651 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6201), .C(n6197), 
        .D(\registers[4][6] ), .Z(n1536) );
  HS65_LH_AO22X9 U1652 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6201), .C(n6197), 
        .D(\registers[4][7] ), .Z(n1537) );
  HS65_LH_AO22X9 U1653 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6201), .C(n6197), 
        .D(\registers[4][8] ), .Z(n1538) );
  HS65_LH_AO22X9 U1654 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6201), .C(n6197), 
        .D(\registers[4][9] ), .Z(n1539) );
  HS65_LH_AO22X9 U1655 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6201), .C(n6197), 
        .D(\registers[4][10] ), .Z(n1540) );
  HS65_LH_AO22X9 U1656 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6200), .C(n6197), 
        .D(\registers[4][11] ), .Z(n1541) );
  HS65_LH_AO22X9 U1657 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6200), .C(n6197), 
        .D(\registers[4][12] ), .Z(n1542) );
  HS65_LH_AO22X9 U1658 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6200), .C(n6198), 
        .D(\registers[4][13] ), .Z(n1543) );
  HS65_LH_AO22X9 U1659 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6200), .C(n6198), 
        .D(\registers[4][14] ), .Z(n1544) );
  HS65_LH_AO22X9 U1660 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6200), .C(n6198), 
        .D(\registers[4][15] ), .Z(n1545) );
  HS65_LH_AO22X9 U1661 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6200), .C(n6198), 
        .D(\registers[4][16] ), .Z(n1546) );
  HS65_LH_AO22X9 U1662 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6200), .C(n6198), 
        .D(\registers[4][17] ), .Z(n1547) );
  HS65_LH_AO22X9 U1663 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6200), .C(n6198), 
        .D(\registers[4][18] ), .Z(n1548) );
  HS65_LH_AO22X9 U1664 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6200), .C(n6198), 
        .D(\registers[4][19] ), .Z(n1549) );
  HS65_LH_AO22X9 U1665 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6200), .C(n6198), 
        .D(\registers[4][20] ), .Z(n1550) );
  HS65_LH_AO22X9 U1666 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6200), .C(n6198), 
        .D(\registers[4][21] ), .Z(n1551) );
  HS65_LH_AO22X9 U1667 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6200), .C(n6198), 
        .D(\registers[4][22] ), .Z(n1552) );
  HS65_LH_AO22X9 U1668 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6200), .C(n6198), 
        .D(\registers[4][23] ), .Z(n1553) );
  HS65_LH_AO22X9 U1669 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6200), .C(n6198), 
        .D(\registers[4][24] ), .Z(n1554) );
  HS65_LH_AO22X9 U1670 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6200), .C(n6198), 
        .D(\registers[4][25] ), .Z(n1555) );
  HS65_LH_AO22X9 U1671 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6200), .C(n6197), 
        .D(\registers[4][26] ), .Z(n1556) );
  HS65_LH_AO22X9 U1672 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6200), .C(n6198), 
        .D(\registers[4][27] ), .Z(n1557) );
  HS65_LH_AO22X9 U1673 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6200), .C(n6197), 
        .D(\registers[4][28] ), .Z(n1558) );
  HS65_LH_AO22X9 U1674 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6200), .C(n6198), 
        .D(\registers[4][29] ), .Z(n1559) );
  HS65_LH_AO22X9 U1675 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6200), .C(n6197), 
        .D(\registers[4][30] ), .Z(n1560) );
  HS65_LH_AO22X9 U1676 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6199), .C(n6198), 
        .D(\registers[4][31] ), .Z(n1561) );
  HS65_LH_AO22X9 U1677 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6236), .C(n6232), 
        .D(\registers[11][0] ), .Z(n1754) );
  HS65_LH_AO22X9 U1678 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6236), .C(n6232), 
        .D(\registers[11][1] ), .Z(n1755) );
  HS65_LH_AO22X9 U1679 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6236), .C(n6232), 
        .D(\registers[11][2] ), .Z(n1756) );
  HS65_LH_AO22X9 U1680 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6236), .C(n6232), 
        .D(\registers[11][3] ), .Z(n1757) );
  HS65_LH_AO22X9 U1681 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6236), .C(n6232), 
        .D(\registers[11][4] ), .Z(n1758) );
  HS65_LH_AO22X9 U1682 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6236), .C(n6232), 
        .D(\registers[11][5] ), .Z(n1759) );
  HS65_LH_AO22X9 U1683 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6236), .C(n6232), 
        .D(\registers[11][6] ), .Z(n1760) );
  HS65_LH_AO22X9 U1684 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6236), .C(n6232), 
        .D(\registers[11][7] ), .Z(n1761) );
  HS65_LH_AO22X9 U1685 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6236), .C(n6232), 
        .D(\registers[11][8] ), .Z(n1762) );
  HS65_LH_AO22X9 U1686 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6236), .C(n6232), 
        .D(\registers[11][9] ), .Z(n1763) );
  HS65_LH_AO22X9 U1687 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6236), .C(n6232), 
        .D(\registers[11][10] ), .Z(n1764) );
  HS65_LH_AO22X9 U1688 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6235), .C(n6232), 
        .D(\registers[11][11] ), .Z(n1765) );
  HS65_LH_AO22X9 U1689 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6235), .C(n6232), 
        .D(\registers[11][12] ), .Z(n1766) );
  HS65_LH_AO22X9 U1690 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6235), .C(n6233), 
        .D(\registers[11][13] ), .Z(n1767) );
  HS65_LH_AO22X9 U1691 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6235), .C(n6233), 
        .D(\registers[11][14] ), .Z(n1768) );
  HS65_LH_AO22X9 U1692 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6235), .C(n6233), 
        .D(\registers[11][15] ), .Z(n1769) );
  HS65_LH_AO22X9 U1693 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6235), .C(n6233), 
        .D(\registers[11][16] ), .Z(n1770) );
  HS65_LH_AO22X9 U1694 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6235), .C(n6233), 
        .D(\registers[11][17] ), .Z(n1771) );
  HS65_LH_AO22X9 U1695 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6235), .C(n6233), 
        .D(\registers[11][18] ), .Z(n1772) );
  HS65_LH_AO22X9 U1696 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6235), .C(n6233), 
        .D(\registers[11][19] ), .Z(n1773) );
  HS65_LH_AO22X9 U1697 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6235), .C(n6233), 
        .D(\registers[11][20] ), .Z(n1774) );
  HS65_LH_AO22X9 U1698 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6235), .C(n6233), 
        .D(\registers[11][21] ), .Z(n1775) );
  HS65_LH_AO22X9 U1699 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6235), .C(n6233), 
        .D(\registers[11][22] ), .Z(n1776) );
  HS65_LH_AO22X9 U1700 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6235), .C(n6233), 
        .D(\registers[11][23] ), .Z(n1777) );
  HS65_LH_AO22X9 U1701 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6235), .C(n6233), 
        .D(\registers[11][24] ), .Z(n1778) );
  HS65_LH_AO22X9 U1702 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6235), .C(n6233), 
        .D(\registers[11][25] ), .Z(n1779) );
  HS65_LH_AO22X9 U1703 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6235), .C(n6232), 
        .D(\registers[11][26] ), .Z(n1780) );
  HS65_LH_AO22X9 U1704 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6235), .C(n6233), 
        .D(\registers[11][27] ), .Z(n1781) );
  HS65_LH_AO22X9 U1705 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6235), .C(n6232), 
        .D(\registers[11][28] ), .Z(n1782) );
  HS65_LH_AO22X9 U1706 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6235), .C(n6233), 
        .D(\registers[11][29] ), .Z(n1783) );
  HS65_LH_AO22X9 U1707 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6235), .C(n6232), 
        .D(\registers[11][30] ), .Z(n1784) );
  HS65_LH_AO22X9 U1708 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6234), .C(n6233), 
        .D(\registers[11][31] ), .Z(n1785) );
  HS65_LH_AO22X9 U1709 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6196), .C(n6192), 
        .D(\registers[3][0] ), .Z(n1498) );
  HS65_LH_AO22X9 U1710 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6196), .C(n6192), 
        .D(\registers[3][1] ), .Z(n1499) );
  HS65_LH_AO22X9 U1711 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6196), .C(n6192), 
        .D(\registers[3][2] ), .Z(n1500) );
  HS65_LH_AO22X9 U1712 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6196), .C(n6192), 
        .D(\registers[3][3] ), .Z(n1501) );
  HS65_LH_AO22X9 U1713 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6196), .C(n6192), 
        .D(\registers[3][4] ), .Z(n1502) );
  HS65_LH_AO22X9 U1714 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6196), .C(n6192), 
        .D(\registers[3][5] ), .Z(n1503) );
  HS65_LH_AO22X9 U1715 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6196), .C(n6192), 
        .D(\registers[3][6] ), .Z(n1504) );
  HS65_LH_AO22X9 U1716 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6196), .C(n6192), 
        .D(\registers[3][7] ), .Z(n1505) );
  HS65_LH_AO22X9 U1717 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6196), .C(n6192), 
        .D(\registers[3][8] ), .Z(n1506) );
  HS65_LH_AO22X9 U1718 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6196), .C(n6192), 
        .D(\registers[3][9] ), .Z(n1507) );
  HS65_LH_AO22X9 U1719 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6196), .C(n6192), 
        .D(\registers[3][10] ), .Z(n1508) );
  HS65_LH_AO22X9 U1720 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6195), .C(n6192), 
        .D(\registers[3][11] ), .Z(n1509) );
  HS65_LH_AO22X9 U1721 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6195), .C(n6192), 
        .D(\registers[3][12] ), .Z(n1510) );
  HS65_LH_AO22X9 U1722 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6195), .C(n6193), 
        .D(\registers[3][13] ), .Z(n1511) );
  HS65_LH_AO22X9 U1723 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6195), .C(n6193), 
        .D(\registers[3][14] ), .Z(n1512) );
  HS65_LH_AO22X9 U1724 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6195), .C(n6193), 
        .D(\registers[3][15] ), .Z(n1513) );
  HS65_LH_AO22X9 U1725 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6195), .C(n6193), 
        .D(\registers[3][16] ), .Z(n1514) );
  HS65_LH_AO22X9 U1726 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6195), .C(n6193), 
        .D(\registers[3][17] ), .Z(n1515) );
  HS65_LH_AO22X9 U1727 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6195), .C(n6193), 
        .D(\registers[3][18] ), .Z(n1516) );
  HS65_LH_AO22X9 U1728 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6195), .C(n6193), 
        .D(\registers[3][19] ), .Z(n1517) );
  HS65_LH_AO22X9 U1729 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6195), .C(n6193), 
        .D(\registers[3][20] ), .Z(n1518) );
  HS65_LH_AO22X9 U1730 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6195), .C(n6193), 
        .D(\registers[3][21] ), .Z(n1519) );
  HS65_LH_AO22X9 U1731 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6195), .C(n6193), 
        .D(\registers[3][22] ), .Z(n1520) );
  HS65_LH_AO22X9 U1732 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6195), .C(n6193), 
        .D(\registers[3][23] ), .Z(n1521) );
  HS65_LH_AO22X9 U1733 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6195), .C(n6193), 
        .D(\registers[3][24] ), .Z(n1522) );
  HS65_LH_AO22X9 U1734 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6195), .C(n6193), 
        .D(\registers[3][25] ), .Z(n1523) );
  HS65_LH_AO22X9 U1735 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6195), .C(n6192), 
        .D(\registers[3][26] ), .Z(n1524) );
  HS65_LH_AO22X9 U1736 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6195), .C(n6193), 
        .D(\registers[3][27] ), .Z(n1525) );
  HS65_LH_AO22X9 U1737 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6195), .C(n6192), 
        .D(\registers[3][28] ), .Z(n1526) );
  HS65_LH_AO22X9 U1738 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6195), .C(n6193), 
        .D(\registers[3][29] ), .Z(n1527) );
  HS65_LH_AO22X9 U1739 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6195), .C(n6192), 
        .D(\registers[3][30] ), .Z(n1528) );
  HS65_LH_AO22X9 U1740 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6194), .C(n6193), 
        .D(\registers[3][31] ), .Z(n1529) );
  HS65_LH_AO22X9 U1741 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6191), .C(n6187), 
        .D(\registers[2][0] ), .Z(n1466) );
  HS65_LH_AO22X9 U1742 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6191), .C(n6187), 
        .D(\registers[2][1] ), .Z(n1467) );
  HS65_LH_AO22X9 U1743 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6191), .C(n6187), 
        .D(\registers[2][2] ), .Z(n1468) );
  HS65_LH_AO22X9 U1744 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6191), .C(n6187), 
        .D(\registers[2][3] ), .Z(n1469) );
  HS65_LH_AO22X9 U1745 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6191), .C(n6187), 
        .D(\registers[2][4] ), .Z(n1470) );
  HS65_LH_AO22X9 U1746 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6191), .C(n6187), 
        .D(\registers[2][5] ), .Z(n1471) );
  HS65_LH_AO22X9 U1747 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6191), .C(n6187), 
        .D(\registers[2][6] ), .Z(n1472) );
  HS65_LH_AO22X9 U1748 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6191), .C(n6187), 
        .D(\registers[2][7] ), .Z(n1473) );
  HS65_LH_AO22X9 U1749 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6191), .C(n6187), 
        .D(\registers[2][8] ), .Z(n1474) );
  HS65_LH_AO22X9 U1750 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6191), .C(n6187), 
        .D(\registers[2][9] ), .Z(n1475) );
  HS65_LH_AO22X9 U1751 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6191), .C(n6187), 
        .D(\registers[2][10] ), .Z(n1476) );
  HS65_LH_AO22X9 U1752 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6190), .C(n6187), 
        .D(\registers[2][11] ), .Z(n1477) );
  HS65_LH_AO22X9 U1753 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6190), .C(n6187), 
        .D(\registers[2][12] ), .Z(n1478) );
  HS65_LH_AO22X9 U1754 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6190), .C(n6188), 
        .D(\registers[2][13] ), .Z(n1479) );
  HS65_LH_AO22X9 U1755 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6190), .C(n6188), 
        .D(\registers[2][14] ), .Z(n1480) );
  HS65_LH_AO22X9 U1756 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6190), .C(n6188), 
        .D(\registers[2][15] ), .Z(n1481) );
  HS65_LH_AO22X9 U1757 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6190), .C(n6188), 
        .D(\registers[2][16] ), .Z(n1482) );
  HS65_LH_AO22X9 U1758 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6190), .C(n6188), 
        .D(\registers[2][17] ), .Z(n1483) );
  HS65_LH_AO22X9 U1759 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6190), .C(n6188), 
        .D(\registers[2][18] ), .Z(n1484) );
  HS65_LH_AO22X9 U1760 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6190), .C(n6188), 
        .D(\registers[2][19] ), .Z(n1485) );
  HS65_LH_AO22X9 U1761 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6190), .C(n6188), 
        .D(\registers[2][20] ), .Z(n1486) );
  HS65_LH_AO22X9 U1762 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6190), .C(n6188), 
        .D(\registers[2][21] ), .Z(n1487) );
  HS65_LH_AO22X9 U1763 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6190), .C(n6188), 
        .D(\registers[2][22] ), .Z(n1488) );
  HS65_LH_AO22X9 U1764 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6190), .C(n6188), 
        .D(\registers[2][23] ), .Z(n1489) );
  HS65_LH_AO22X9 U1765 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6190), .C(n6188), 
        .D(\registers[2][24] ), .Z(n1490) );
  HS65_LH_AO22X9 U1766 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6190), .C(n6188), 
        .D(\registers[2][25] ), .Z(n1491) );
  HS65_LH_AO22X9 U1767 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6190), .C(n6187), 
        .D(\registers[2][26] ), .Z(n1492) );
  HS65_LH_AO22X9 U1768 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6190), .C(n6188), 
        .D(\registers[2][27] ), .Z(n1493) );
  HS65_LH_AO22X9 U1769 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6190), .C(n6187), 
        .D(\registers[2][28] ), .Z(n1494) );
  HS65_LH_AO22X9 U1770 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6190), .C(n6188), 
        .D(\registers[2][29] ), .Z(n1495) );
  HS65_LH_AO22X9 U1771 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6190), .C(n6187), 
        .D(\registers[2][30] ), .Z(n1496) );
  HS65_LH_AO22X9 U1772 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6189), .C(n6188), 
        .D(\registers[2][31] ), .Z(n1497) );
  HS65_LH_AO22X9 U1773 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n6206), .C(n6202), 
        .D(\registers[5][0] ), .Z(n1562) );
  HS65_LH_AO22X9 U1774 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n6206), .C(n6202), 
        .D(\registers[5][1] ), .Z(n1563) );
  HS65_LH_AO22X9 U1775 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n6206), .C(n6202), 
        .D(\registers[5][2] ), .Z(n1564) );
  HS65_LH_AO22X9 U1776 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n6206), .C(n6202), 
        .D(\registers[5][3] ), .Z(n1565) );
  HS65_LH_AO22X9 U1777 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n6206), .C(n6202), 
        .D(\registers[5][4] ), .Z(n1566) );
  HS65_LH_AO22X9 U1778 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n6206), .C(n6202), 
        .D(\registers[5][5] ), .Z(n1567) );
  HS65_LH_AO22X9 U1779 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n6206), .C(n6202), 
        .D(\registers[5][6] ), .Z(n1568) );
  HS65_LH_AO22X9 U1780 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n6206), .C(n6202), 
        .D(\registers[5][7] ), .Z(n1569) );
  HS65_LH_AO22X9 U1781 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n6206), .C(n6202), 
        .D(\registers[5][8] ), .Z(n1570) );
  HS65_LH_AO22X9 U1782 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n6206), .C(n6202), 
        .D(\registers[5][9] ), .Z(n1571) );
  HS65_LH_AO22X9 U1783 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n6206), .C(n6202), 
        .D(\registers[5][10] ), .Z(n1572) );
  HS65_LH_AO22X9 U1784 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n6205), .C(n6202), 
        .D(\registers[5][11] ), .Z(n1573) );
  HS65_LH_AO22X9 U1785 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n6205), .C(n6202), 
        .D(\registers[5][12] ), .Z(n1574) );
  HS65_LH_AO22X9 U1786 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n6205), .C(n6203), 
        .D(\registers[5][13] ), .Z(n1575) );
  HS65_LH_AO22X9 U1787 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n6205), .C(n6203), 
        .D(\registers[5][14] ), .Z(n1576) );
  HS65_LH_AO22X9 U1788 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n6205), .C(n6203), 
        .D(\registers[5][15] ), .Z(n1577) );
  HS65_LH_AO22X9 U1789 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n6205), .C(n6203), 
        .D(\registers[5][16] ), .Z(n1578) );
  HS65_LH_AO22X9 U1790 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n6205), .C(n6203), 
        .D(\registers[5][17] ), .Z(n1579) );
  HS65_LH_AO22X9 U1791 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n6205), .C(n6203), 
        .D(\registers[5][18] ), .Z(n1580) );
  HS65_LH_AO22X9 U1792 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n6205), .C(n6203), 
        .D(\registers[5][19] ), .Z(n1581) );
  HS65_LH_AO22X9 U1793 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n6205), .C(n6203), 
        .D(\registers[5][20] ), .Z(n1582) );
  HS65_LH_AO22X9 U1794 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n6205), .C(n6203), 
        .D(\registers[5][21] ), .Z(n1583) );
  HS65_LH_AO22X9 U1795 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n6205), .C(n6203), 
        .D(\registers[5][22] ), .Z(n1584) );
  HS65_LH_AO22X9 U1796 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n6205), .C(n6203), 
        .D(\registers[5][23] ), .Z(n1585) );
  HS65_LH_AO22X9 U1797 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n6205), .C(n6203), 
        .D(\registers[5][24] ), .Z(n1586) );
  HS65_LH_AO22X9 U1798 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n6205), .C(n6203), 
        .D(\registers[5][25] ), .Z(n1587) );
  HS65_LH_AO22X9 U1799 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n6205), .C(n6202), 
        .D(\registers[5][26] ), .Z(n1588) );
  HS65_LH_AO22X9 U1800 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n6205), .C(n6203), 
        .D(\registers[5][27] ), .Z(n1589) );
  HS65_LH_AO22X9 U1801 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n6205), .C(n6202), 
        .D(\registers[5][28] ), .Z(n1590) );
  HS65_LH_AO22X9 U1802 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n6205), .C(n6203), 
        .D(\registers[5][29] ), .Z(n1591) );
  HS65_LH_AO22X9 U1803 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n6205), .C(n6202), 
        .D(\registers[5][30] ), .Z(n1592) );
  HS65_LH_AO22X9 U1804 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n6204), .C(n6203), 
        .D(\registers[5][31] ), .Z(n1593) );
  HS65_LH_AO22X9 U1805 ( .A(n6182), .B(\registers[1][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6186), .Z(n1434) );
  HS65_LH_AO22X9 U1806 ( .A(n6182), .B(\registers[1][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6186), .Z(n1435) );
  HS65_LH_AO22X9 U1807 ( .A(n6182), .B(\registers[1][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6186), .Z(n1436) );
  HS65_LH_AO22X9 U1808 ( .A(n6182), .B(\registers[1][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6186), .Z(n1437) );
  HS65_LH_AO22X9 U1809 ( .A(n6182), .B(\registers[1][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6186), .Z(n1438) );
  HS65_LH_AO22X9 U1810 ( .A(n6182), .B(\registers[1][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6186), .Z(n1439) );
  HS65_LH_AO22X9 U1811 ( .A(n6182), .B(\registers[1][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6186), .Z(n1440) );
  HS65_LH_AO22X9 U1812 ( .A(n6182), .B(\registers[1][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6186), .Z(n1441) );
  HS65_LH_AO22X9 U1813 ( .A(n6182), .B(\registers[1][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6186), .Z(n1442) );
  HS65_LH_AO22X9 U1814 ( .A(n6182), .B(\registers[1][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6186), .Z(n1443) );
  HS65_LH_AO22X9 U1815 ( .A(n6182), .B(\registers[1][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6186), .Z(n1444) );
  HS65_LH_AO22X9 U1816 ( .A(n6182), .B(\registers[1][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6185), .Z(n1445) );
  HS65_LH_AO22X9 U1817 ( .A(n6183), .B(\registers[1][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6185), .Z(n1446) );
  HS65_LH_AO22X9 U1818 ( .A(n6183), .B(\registers[1][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6185), .Z(n1447) );
  HS65_LH_AO22X9 U1819 ( .A(n6183), .B(\registers[1][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6185), .Z(n1448) );
  HS65_LH_AO22X9 U1820 ( .A(n6183), .B(\registers[1][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6185), .Z(n1449) );
  HS65_LH_AO22X9 U1821 ( .A(n6183), .B(\registers[1][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6185), .Z(n1450) );
  HS65_LH_AO22X9 U1822 ( .A(n6183), .B(\registers[1][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6185), .Z(n1451) );
  HS65_LH_AO22X9 U1823 ( .A(n6183), .B(\registers[1][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6185), .Z(n1452) );
  HS65_LH_AO22X9 U1824 ( .A(n6183), .B(\registers[1][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6185), .Z(n1453) );
  HS65_LH_AO22X9 U1825 ( .A(n6183), .B(\registers[1][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6185), .Z(n1454) );
  HS65_LH_AO22X9 U1826 ( .A(n6183), .B(\registers[1][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6185), .Z(n1455) );
  HS65_LH_AO22X9 U1827 ( .A(n6183), .B(\registers[1][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6185), .Z(n1456) );
  HS65_LH_AO22X9 U1828 ( .A(n6183), .B(\registers[1][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6185), .Z(n1457) );
  HS65_LH_AO22X9 U1829 ( .A(n6182), .B(\registers[1][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6185), .Z(n1458) );
  HS65_LH_AO22X9 U1830 ( .A(n6183), .B(\registers[1][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6185), .Z(n1459) );
  HS65_LH_AO22X9 U1831 ( .A(n6182), .B(\registers[1][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6185), .Z(n1460) );
  HS65_LH_AO22X9 U1832 ( .A(n6183), .B(\registers[1][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6185), .Z(n1461) );
  HS65_LH_AO22X9 U1833 ( .A(n6182), .B(\registers[1][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6185), .Z(n1462) );
  HS65_LH_AO22X9 U1834 ( .A(n6183), .B(\registers[1][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6185), .Z(n1463) );
  HS65_LH_AO22X9 U1835 ( .A(n6182), .B(\registers[1][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6185), .Z(n1464) );
  HS65_LH_AO22X9 U1836 ( .A(n6183), .B(\registers[1][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6184), .Z(n1465) );
  HS65_LH_AO22X9 U1837 ( .A(n6332), .B(\registers[31][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6336), .Z(n2394) );
  HS65_LH_AO22X9 U1838 ( .A(n6332), .B(\registers[31][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6336), .Z(n2395) );
  HS65_LH_AO22X9 U1839 ( .A(n6332), .B(\registers[31][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6336), .Z(n2396) );
  HS65_LH_AO22X9 U1840 ( .A(n6332), .B(\registers[31][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6336), .Z(n2397) );
  HS65_LH_AO22X9 U1841 ( .A(n6332), .B(\registers[31][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6336), .Z(n2398) );
  HS65_LH_AO22X9 U1842 ( .A(n6332), .B(\registers[31][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6336), .Z(n2399) );
  HS65_LH_AO22X9 U1843 ( .A(n6332), .B(\registers[31][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6336), .Z(n2400) );
  HS65_LH_AO22X9 U1844 ( .A(n6332), .B(\registers[31][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6336), .Z(n2401) );
  HS65_LH_AO22X9 U1845 ( .A(n6332), .B(\registers[31][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6336), .Z(n2402) );
  HS65_LH_AO22X9 U1846 ( .A(n6332), .B(\registers[31][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6336), .Z(n2403) );
  HS65_LH_AO22X9 U1847 ( .A(n6332), .B(\registers[31][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6336), .Z(n2404) );
  HS65_LH_AO22X9 U1848 ( .A(n6332), .B(\registers[31][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6335), .Z(n2405) );
  HS65_LH_AO22X9 U1849 ( .A(n6333), .B(\registers[31][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6335), .Z(n2406) );
  HS65_LH_AO22X9 U1850 ( .A(n6333), .B(\registers[31][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6335), .Z(n2407) );
  HS65_LH_AO22X9 U1851 ( .A(n6333), .B(\registers[31][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6335), .Z(n2408) );
  HS65_LH_AO22X9 U1852 ( .A(n6333), .B(\registers[31][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6335), .Z(n2409) );
  HS65_LH_AO22X9 U1853 ( .A(n6333), .B(\registers[31][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6335), .Z(n2410) );
  HS65_LH_AO22X9 U1854 ( .A(n6333), .B(\registers[31][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6335), .Z(n2411) );
  HS65_LH_AO22X9 U1855 ( .A(n6333), .B(\registers[31][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6335), .Z(n2412) );
  HS65_LH_AO22X9 U1856 ( .A(n6333), .B(\registers[31][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6335), .Z(n2413) );
  HS65_LH_AO22X9 U1857 ( .A(n6333), .B(\registers[31][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6335), .Z(n2414) );
  HS65_LH_AO22X9 U1858 ( .A(n6333), .B(\registers[31][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6335), .Z(n2415) );
  HS65_LH_AO22X9 U1859 ( .A(n6333), .B(\registers[31][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6335), .Z(n2416) );
  HS65_LH_AO22X9 U1860 ( .A(n6333), .B(\registers[31][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6335), .Z(n2417) );
  HS65_LH_AO22X9 U1861 ( .A(n6332), .B(\registers[31][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6335), .Z(n2418) );
  HS65_LH_AO22X9 U1862 ( .A(n6333), .B(\registers[31][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6335), .Z(n2419) );
  HS65_LH_AO22X9 U1863 ( .A(n6332), .B(\registers[31][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6335), .Z(n2420) );
  HS65_LH_AO22X9 U1864 ( .A(n6333), .B(\registers[31][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6335), .Z(n2421) );
  HS65_LH_AO22X9 U1865 ( .A(n6332), .B(\registers[31][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6335), .Z(n2422) );
  HS65_LH_AO22X9 U1866 ( .A(n6333), .B(\registers[31][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6335), .Z(n2423) );
  HS65_LH_AO22X9 U1867 ( .A(n6332), .B(\registers[31][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6335), .Z(n2424) );
  HS65_LH_AO22X9 U1868 ( .A(n6333), .B(\registers[31][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6334), .Z(n2425) );
  HS65_LH_AO22X9 U1869 ( .A(n6272), .B(\registers[19][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6276), .Z(n2010) );
  HS65_LH_AO22X9 U1870 ( .A(n6272), .B(\registers[19][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6276), .Z(n2011) );
  HS65_LH_AO22X9 U1871 ( .A(n6272), .B(\registers[19][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6276), .Z(n2012) );
  HS65_LH_AO22X9 U1872 ( .A(n6272), .B(\registers[19][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6276), .Z(n2013) );
  HS65_LH_AO22X9 U1873 ( .A(n6272), .B(\registers[19][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6276), .Z(n2014) );
  HS65_LH_AO22X9 U1874 ( .A(n6272), .B(\registers[19][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6276), .Z(n2015) );
  HS65_LH_AO22X9 U1875 ( .A(n6272), .B(\registers[19][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6276), .Z(n2016) );
  HS65_LH_AO22X9 U1876 ( .A(n6272), .B(\registers[19][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6276), .Z(n2017) );
  HS65_LH_AO22X9 U1877 ( .A(n6272), .B(\registers[19][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6276), .Z(n2018) );
  HS65_LH_AO22X9 U1878 ( .A(n6272), .B(\registers[19][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6276), .Z(n2019) );
  HS65_LH_AO22X9 U1879 ( .A(n6272), .B(\registers[19][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6276), .Z(n2020) );
  HS65_LH_AO22X9 U1880 ( .A(n6272), .B(\registers[19][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6275), .Z(n2021) );
  HS65_LH_AO22X9 U1881 ( .A(n6273), .B(\registers[19][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6275), .Z(n2022) );
  HS65_LH_AO22X9 U1882 ( .A(n6273), .B(\registers[19][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6275), .Z(n2023) );
  HS65_LH_AO22X9 U1883 ( .A(n6273), .B(\registers[19][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6275), .Z(n2024) );
  HS65_LH_AO22X9 U1884 ( .A(n6273), .B(\registers[19][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6275), .Z(n2025) );
  HS65_LH_AO22X9 U1885 ( .A(n6273), .B(\registers[19][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6275), .Z(n2026) );
  HS65_LH_AO22X9 U1886 ( .A(n6273), .B(\registers[19][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6275), .Z(n2027) );
  HS65_LH_AO22X9 U1887 ( .A(n6273), .B(\registers[19][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6275), .Z(n2028) );
  HS65_LH_AO22X9 U1888 ( .A(n6273), .B(\registers[19][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6275), .Z(n2029) );
  HS65_LH_AO22X9 U1889 ( .A(n6273), .B(\registers[19][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6275), .Z(n2030) );
  HS65_LH_AO22X9 U1890 ( .A(n6273), .B(\registers[19][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6275), .Z(n2031) );
  HS65_LH_AO22X9 U1891 ( .A(n6273), .B(\registers[19][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6275), .Z(n2032) );
  HS65_LH_AO22X9 U1892 ( .A(n6273), .B(\registers[19][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6275), .Z(n2033) );
  HS65_LH_AO22X9 U1893 ( .A(n6272), .B(\registers[19][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6275), .Z(n2034) );
  HS65_LH_AO22X9 U1894 ( .A(n6273), .B(\registers[19][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6275), .Z(n2035) );
  HS65_LH_AO22X9 U1895 ( .A(n6272), .B(\registers[19][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6275), .Z(n2036) );
  HS65_LH_AO22X9 U1896 ( .A(n6273), .B(\registers[19][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6275), .Z(n2037) );
  HS65_LH_AO22X9 U1897 ( .A(n6272), .B(\registers[19][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6275), .Z(n2038) );
  HS65_LH_AO22X9 U1898 ( .A(n6273), .B(\registers[19][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6275), .Z(n2039) );
  HS65_LH_AO22X9 U1899 ( .A(n6272), .B(\registers[19][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6275), .Z(n2040) );
  HS65_LH_AO22X9 U1900 ( .A(n6273), .B(\registers[19][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6274), .Z(n2041) );
  HS65_LH_AO22X9 U1901 ( .A(n6212), .B(\registers[7][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6216), .Z(n1626) );
  HS65_LH_AO22X9 U1902 ( .A(n6212), .B(\registers[7][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6216), .Z(n1627) );
  HS65_LH_AO22X9 U1903 ( .A(n6212), .B(\registers[7][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6216), .Z(n1628) );
  HS65_LH_AO22X9 U1904 ( .A(n6212), .B(\registers[7][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6216), .Z(n1629) );
  HS65_LH_AO22X9 U1905 ( .A(n6212), .B(\registers[7][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6216), .Z(n1630) );
  HS65_LH_AO22X9 U1906 ( .A(n6212), .B(\registers[7][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6216), .Z(n1631) );
  HS65_LH_AO22X9 U1907 ( .A(n6212), .B(\registers[7][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6216), .Z(n1632) );
  HS65_LH_AO22X9 U1908 ( .A(n6212), .B(\registers[7][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6216), .Z(n1633) );
  HS65_LH_AO22X9 U1909 ( .A(n6212), .B(\registers[7][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6216), .Z(n1634) );
  HS65_LH_AO22X9 U1910 ( .A(n6212), .B(\registers[7][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6216), .Z(n1635) );
  HS65_LH_AO22X9 U1911 ( .A(n6212), .B(\registers[7][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6216), .Z(n1636) );
  HS65_LH_AO22X9 U1912 ( .A(n6212), .B(\registers[7][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6215), .Z(n1637) );
  HS65_LH_AO22X9 U1913 ( .A(n6213), .B(\registers[7][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6215), .Z(n1638) );
  HS65_LH_AO22X9 U1914 ( .A(n6213), .B(\registers[7][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6215), .Z(n1639) );
  HS65_LH_AO22X9 U1915 ( .A(n6213), .B(\registers[7][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6215), .Z(n1640) );
  HS65_LH_AO22X9 U1916 ( .A(n6213), .B(\registers[7][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6215), .Z(n1641) );
  HS65_LH_AO22X9 U1917 ( .A(n6213), .B(\registers[7][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6215), .Z(n1642) );
  HS65_LH_AO22X9 U1918 ( .A(n6213), .B(\registers[7][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6215), .Z(n1643) );
  HS65_LH_AO22X9 U1919 ( .A(n6213), .B(\registers[7][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6215), .Z(n1644) );
  HS65_LH_AO22X9 U1920 ( .A(n6213), .B(\registers[7][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6215), .Z(n1645) );
  HS65_LH_AO22X9 U1921 ( .A(n6213), .B(\registers[7][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6215), .Z(n1646) );
  HS65_LH_AO22X9 U1922 ( .A(n6213), .B(\registers[7][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6215), .Z(n1647) );
  HS65_LH_AO22X9 U1923 ( .A(n6213), .B(\registers[7][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6215), .Z(n1648) );
  HS65_LH_AO22X9 U1924 ( .A(n6213), .B(\registers[7][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6215), .Z(n1649) );
  HS65_LH_AO22X9 U1925 ( .A(n6212), .B(\registers[7][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6215), .Z(n1650) );
  HS65_LH_AO22X9 U1926 ( .A(n6213), .B(\registers[7][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6215), .Z(n1651) );
  HS65_LH_AO22X9 U1927 ( .A(n6212), .B(\registers[7][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6215), .Z(n1652) );
  HS65_LH_AO22X9 U1928 ( .A(n6213), .B(\registers[7][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6215), .Z(n1653) );
  HS65_LH_AO22X9 U1929 ( .A(n6212), .B(\registers[7][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6215), .Z(n1654) );
  HS65_LH_AO22X9 U1930 ( .A(n6213), .B(\registers[7][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6215), .Z(n1655) );
  HS65_LH_AO22X9 U1931 ( .A(n6212), .B(\registers[7][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6215), .Z(n1656) );
  HS65_LH_AO22X9 U1932 ( .A(n6213), .B(\registers[7][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6214), .Z(n1657) );
  HS65_LH_AO22X9 U1933 ( .A(n6277), .B(\registers[20][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6281), .Z(n2042) );
  HS65_LH_AO22X9 U1934 ( .A(n6277), .B(\registers[20][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6281), .Z(n2043) );
  HS65_LH_AO22X9 U1935 ( .A(n6277), .B(\registers[20][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6281), .Z(n2044) );
  HS65_LH_AO22X9 U1936 ( .A(n6277), .B(\registers[20][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6281), .Z(n2045) );
  HS65_LH_AO22X9 U1937 ( .A(n6277), .B(\registers[20][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6281), .Z(n2046) );
  HS65_LH_AO22X9 U1938 ( .A(n6277), .B(\registers[20][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6281), .Z(n2047) );
  HS65_LH_AO22X9 U1939 ( .A(n6277), .B(\registers[20][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6281), .Z(n2048) );
  HS65_LH_AO22X9 U1940 ( .A(n6277), .B(\registers[20][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6281), .Z(n2049) );
  HS65_LH_AO22X9 U1941 ( .A(n6277), .B(\registers[20][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6281), .Z(n2050) );
  HS65_LH_AO22X9 U1942 ( .A(n6277), .B(\registers[20][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6281), .Z(n2051) );
  HS65_LH_AO22X9 U1943 ( .A(n6277), .B(\registers[20][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6281), .Z(n2052) );
  HS65_LH_AO22X9 U1944 ( .A(n6277), .B(\registers[20][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6280), .Z(n2053) );
  HS65_LH_AO22X9 U1945 ( .A(n6278), .B(\registers[20][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6280), .Z(n2054) );
  HS65_LH_AO22X9 U1946 ( .A(n6278), .B(\registers[20][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6280), .Z(n2055) );
  HS65_LH_AO22X9 U1947 ( .A(n6278), .B(\registers[20][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6280), .Z(n2056) );
  HS65_LH_AO22X9 U1948 ( .A(n6278), .B(\registers[20][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6280), .Z(n2057) );
  HS65_LH_AO22X9 U1949 ( .A(n6278), .B(\registers[20][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6280), .Z(n2058) );
  HS65_LH_AO22X9 U1950 ( .A(n6278), .B(\registers[20][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6280), .Z(n2059) );
  HS65_LH_AO22X9 U1951 ( .A(n6278), .B(\registers[20][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6280), .Z(n2060) );
  HS65_LH_AO22X9 U1952 ( .A(n6278), .B(\registers[20][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6280), .Z(n2061) );
  HS65_LH_AO22X9 U1953 ( .A(n6278), .B(\registers[20][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6280), .Z(n2062) );
  HS65_LH_AO22X9 U1954 ( .A(n6278), .B(\registers[20][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6280), .Z(n2063) );
  HS65_LH_AO22X9 U1955 ( .A(n6278), .B(\registers[20][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6280), .Z(n2064) );
  HS65_LH_AO22X9 U1956 ( .A(n6278), .B(\registers[20][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6280), .Z(n2065) );
  HS65_LH_AO22X9 U1957 ( .A(n6277), .B(\registers[20][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6280), .Z(n2066) );
  HS65_LH_AO22X9 U1958 ( .A(n6278), .B(\registers[20][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6280), .Z(n2067) );
  HS65_LH_AO22X9 U1959 ( .A(n6277), .B(\registers[20][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6280), .Z(n2068) );
  HS65_LH_AO22X9 U1960 ( .A(n6278), .B(\registers[20][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6280), .Z(n2069) );
  HS65_LH_AO22X9 U1961 ( .A(n6277), .B(\registers[20][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6280), .Z(n2070) );
  HS65_LH_AO22X9 U1962 ( .A(n6278), .B(\registers[20][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6280), .Z(n2071) );
  HS65_LH_AO22X9 U1963 ( .A(n6277), .B(\registers[20][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6280), .Z(n2072) );
  HS65_LH_AO22X9 U1964 ( .A(n6278), .B(\registers[20][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6279), .Z(n2073) );
  HS65_LH_AO22X9 U1965 ( .A(n6282), .B(\registers[21][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6286), .Z(n2074) );
  HS65_LH_AO22X9 U1966 ( .A(n6282), .B(\registers[21][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6286), .Z(n2075) );
  HS65_LH_AO22X9 U1967 ( .A(n6282), .B(\registers[21][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6286), .Z(n2076) );
  HS65_LH_AO22X9 U1968 ( .A(n6282), .B(\registers[21][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6286), .Z(n2077) );
  HS65_LH_AO22X9 U1969 ( .A(n6282), .B(\registers[21][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6286), .Z(n2078) );
  HS65_LH_AO22X9 U1970 ( .A(n6282), .B(\registers[21][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6286), .Z(n2079) );
  HS65_LH_AO22X9 U1971 ( .A(n6282), .B(\registers[21][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6286), .Z(n2080) );
  HS65_LH_AO22X9 U1972 ( .A(n6282), .B(\registers[21][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6286), .Z(n2081) );
  HS65_LH_AO22X9 U1973 ( .A(n6282), .B(\registers[21][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6286), .Z(n2082) );
  HS65_LH_AO22X9 U1974 ( .A(n6282), .B(\registers[21][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6286), .Z(n2083) );
  HS65_LH_AO22X9 U1975 ( .A(n6282), .B(\registers[21][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6286), .Z(n2084) );
  HS65_LH_AO22X9 U1976 ( .A(n6282), .B(\registers[21][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6285), .Z(n2085) );
  HS65_LH_AO22X9 U1977 ( .A(n6283), .B(\registers[21][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6285), .Z(n2086) );
  HS65_LH_AO22X9 U1978 ( .A(n6283), .B(\registers[21][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6285), .Z(n2087) );
  HS65_LH_AO22X9 U1979 ( .A(n6283), .B(\registers[21][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6285), .Z(n2088) );
  HS65_LH_AO22X9 U1980 ( .A(n6283), .B(\registers[21][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6285), .Z(n2089) );
  HS65_LH_AO22X9 U1981 ( .A(n6283), .B(\registers[21][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6285), .Z(n2090) );
  HS65_LH_AO22X9 U1982 ( .A(n6283), .B(\registers[21][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6285), .Z(n2091) );
  HS65_LH_AO22X9 U1983 ( .A(n6283), .B(\registers[21][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6285), .Z(n2092) );
  HS65_LH_AO22X9 U1984 ( .A(n6283), .B(\registers[21][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6285), .Z(n2093) );
  HS65_LH_AO22X9 U1985 ( .A(n6283), .B(\registers[21][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6285), .Z(n2094) );
  HS65_LH_AO22X9 U1986 ( .A(n6283), .B(\registers[21][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6285), .Z(n2095) );
  HS65_LH_AO22X9 U1987 ( .A(n6283), .B(\registers[21][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6285), .Z(n2096) );
  HS65_LH_AO22X9 U1988 ( .A(n6283), .B(\registers[21][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6285), .Z(n2097) );
  HS65_LH_AO22X9 U1989 ( .A(n6282), .B(\registers[21][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6285), .Z(n2098) );
  HS65_LH_AO22X9 U1990 ( .A(n6283), .B(\registers[21][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6285), .Z(n2099) );
  HS65_LH_AO22X9 U1991 ( .A(n6282), .B(\registers[21][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6285), .Z(n2100) );
  HS65_LH_AO22X9 U1992 ( .A(n6283), .B(\registers[21][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6285), .Z(n2101) );
  HS65_LH_AO22X9 U1993 ( .A(n6282), .B(\registers[21][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6285), .Z(n2102) );
  HS65_LH_AO22X9 U1994 ( .A(n6283), .B(\registers[21][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6285), .Z(n2103) );
  HS65_LH_AO22X9 U1995 ( .A(n6282), .B(\registers[21][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6285), .Z(n2104) );
  HS65_LH_AO22X9 U1996 ( .A(n6283), .B(\registers[21][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6284), .Z(n2105) );
  HS65_LH_AO22X9 U1997 ( .A(n6327), .B(\registers[30][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6331), .Z(n2362) );
  HS65_LH_AO22X9 U1998 ( .A(n6327), .B(\registers[30][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6331), .Z(n2363) );
  HS65_LH_AO22X9 U1999 ( .A(n6327), .B(\registers[30][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6331), .Z(n2364) );
  HS65_LH_AO22X9 U2000 ( .A(n6327), .B(\registers[30][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6331), .Z(n2365) );
  HS65_LH_AO22X9 U2001 ( .A(n6327), .B(\registers[30][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6331), .Z(n2366) );
  HS65_LH_AO22X9 U2002 ( .A(n6327), .B(\registers[30][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6331), .Z(n2367) );
  HS65_LH_AO22X9 U2003 ( .A(n6327), .B(\registers[30][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6331), .Z(n2368) );
  HS65_LH_AO22X9 U2004 ( .A(n6327), .B(\registers[30][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6331), .Z(n2369) );
  HS65_LH_AO22X9 U2005 ( .A(n6327), .B(\registers[30][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6331), .Z(n2370) );
  HS65_LH_AO22X9 U2006 ( .A(n6327), .B(\registers[30][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6331), .Z(n2371) );
  HS65_LH_AO22X9 U2007 ( .A(n6327), .B(\registers[30][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6331), .Z(n2372) );
  HS65_LH_AO22X9 U2008 ( .A(n6327), .B(\registers[30][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6330), .Z(n2373) );
  HS65_LH_AO22X9 U2009 ( .A(n6328), .B(\registers[30][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6330), .Z(n2374) );
  HS65_LH_AO22X9 U2010 ( .A(n6328), .B(\registers[30][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6330), .Z(n2375) );
  HS65_LH_AO22X9 U2011 ( .A(n6328), .B(\registers[30][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6330), .Z(n2376) );
  HS65_LH_AO22X9 U2012 ( .A(n6328), .B(\registers[30][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6330), .Z(n2377) );
  HS65_LH_AO22X9 U2013 ( .A(n6328), .B(\registers[30][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6330), .Z(n2378) );
  HS65_LH_AO22X9 U2014 ( .A(n6328), .B(\registers[30][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6330), .Z(n2379) );
  HS65_LH_AO22X9 U2015 ( .A(n6328), .B(\registers[30][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6330), .Z(n2380) );
  HS65_LH_AO22X9 U2016 ( .A(n6328), .B(\registers[30][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6330), .Z(n2381) );
  HS65_LH_AO22X9 U2017 ( .A(n6328), .B(\registers[30][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6330), .Z(n2382) );
  HS65_LH_AO22X9 U2018 ( .A(n6328), .B(\registers[30][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6330), .Z(n2383) );
  HS65_LH_AO22X9 U2019 ( .A(n6328), .B(\registers[30][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6330), .Z(n2384) );
  HS65_LH_AO22X9 U2020 ( .A(n6328), .B(\registers[30][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6330), .Z(n2385) );
  HS65_LH_AO22X9 U2021 ( .A(n6327), .B(\registers[30][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6330), .Z(n2386) );
  HS65_LH_AO22X9 U2022 ( .A(n6328), .B(\registers[30][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6330), .Z(n2387) );
  HS65_LH_AO22X9 U2023 ( .A(n6327), .B(\registers[30][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6330), .Z(n2388) );
  HS65_LH_AO22X9 U2024 ( .A(n6328), .B(\registers[30][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6330), .Z(n2389) );
  HS65_LH_AO22X9 U2025 ( .A(n6327), .B(\registers[30][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6330), .Z(n2390) );
  HS65_LH_AO22X9 U2026 ( .A(n6328), .B(\registers[30][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6330), .Z(n2391) );
  HS65_LH_AO22X9 U2027 ( .A(n6327), .B(\registers[30][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6330), .Z(n2392) );
  HS65_LH_AO22X9 U2028 ( .A(n6328), .B(\registers[30][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6329), .Z(n2393) );
  HS65_LH_AO22X9 U2029 ( .A(n6292), .B(\registers[23][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6296), .Z(n2138) );
  HS65_LH_AO22X9 U2030 ( .A(n6292), .B(\registers[23][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6296), .Z(n2139) );
  HS65_LH_AO22X9 U2031 ( .A(n6292), .B(\registers[23][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6296), .Z(n2140) );
  HS65_LH_AO22X9 U2032 ( .A(n6292), .B(\registers[23][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6296), .Z(n2141) );
  HS65_LH_AO22X9 U2033 ( .A(n6292), .B(\registers[23][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6296), .Z(n2142) );
  HS65_LH_AO22X9 U2034 ( .A(n6292), .B(\registers[23][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6296), .Z(n2143) );
  HS65_LH_AO22X9 U2035 ( .A(n6292), .B(\registers[23][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6296), .Z(n2144) );
  HS65_LH_AO22X9 U2036 ( .A(n6292), .B(\registers[23][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6296), .Z(n2145) );
  HS65_LH_AO22X9 U2037 ( .A(n6292), .B(\registers[23][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6296), .Z(n2146) );
  HS65_LH_AO22X9 U2038 ( .A(n6292), .B(\registers[23][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6296), .Z(n2147) );
  HS65_LH_AO22X9 U2039 ( .A(n6292), .B(\registers[23][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6296), .Z(n2148) );
  HS65_LH_AO22X9 U2040 ( .A(n6292), .B(\registers[23][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6295), .Z(n2149) );
  HS65_LH_AO22X9 U2041 ( .A(n6293), .B(\registers[23][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6295), .Z(n2150) );
  HS65_LH_AO22X9 U2042 ( .A(n6293), .B(\registers[23][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6295), .Z(n2151) );
  HS65_LH_AO22X9 U2043 ( .A(n6293), .B(\registers[23][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6295), .Z(n2152) );
  HS65_LH_AO22X9 U2044 ( .A(n6293), .B(\registers[23][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6295), .Z(n2153) );
  HS65_LH_AO22X9 U2045 ( .A(n6293), .B(\registers[23][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6295), .Z(n2154) );
  HS65_LH_AO22X9 U2046 ( .A(n6293), .B(\registers[23][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6295), .Z(n2155) );
  HS65_LH_AO22X9 U2047 ( .A(n6293), .B(\registers[23][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6295), .Z(n2156) );
  HS65_LH_AO22X9 U2048 ( .A(n6293), .B(\registers[23][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6295), .Z(n2157) );
  HS65_LH_AO22X9 U2049 ( .A(n6293), .B(\registers[23][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6295), .Z(n2158) );
  HS65_LH_AO22X9 U2050 ( .A(n6293), .B(\registers[23][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6295), .Z(n2159) );
  HS65_LH_AO22X9 U2051 ( .A(n6293), .B(\registers[23][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6295), .Z(n2160) );
  HS65_LH_AO22X9 U2052 ( .A(n6293), .B(\registers[23][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6295), .Z(n2161) );
  HS65_LH_AO22X9 U2053 ( .A(n6292), .B(\registers[23][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6295), .Z(n2162) );
  HS65_LH_AO22X9 U2054 ( .A(n6293), .B(\registers[23][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6295), .Z(n2163) );
  HS65_LH_AO22X9 U2055 ( .A(n6292), .B(\registers[23][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6295), .Z(n2164) );
  HS65_LH_AO22X9 U2056 ( .A(n6293), .B(\registers[23][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6295), .Z(n2165) );
  HS65_LH_AO22X9 U2057 ( .A(n6292), .B(\registers[23][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6295), .Z(n2166) );
  HS65_LH_AO22X9 U2058 ( .A(n6293), .B(\registers[23][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6295), .Z(n2167) );
  HS65_LH_AO22X9 U2059 ( .A(n6292), .B(\registers[23][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6295), .Z(n2168) );
  HS65_LH_AO22X9 U2060 ( .A(n6293), .B(\registers[23][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6294), .Z(n2169) );
  HS65_LH_AO22X9 U2061 ( .A(n6287), .B(\registers[22][0] ), .C(
        \regfile_i[WRITE_DATA][0] ), .D(n6291), .Z(n2106) );
  HS65_LH_AO22X9 U2062 ( .A(n6287), .B(\registers[22][1] ), .C(
        \regfile_i[WRITE_DATA][1] ), .D(n6291), .Z(n2107) );
  HS65_LH_AO22X9 U2063 ( .A(n6287), .B(\registers[22][2] ), .C(
        \regfile_i[WRITE_DATA][2] ), .D(n6291), .Z(n2108) );
  HS65_LH_AO22X9 U2064 ( .A(n6287), .B(\registers[22][3] ), .C(
        \regfile_i[WRITE_DATA][3] ), .D(n6291), .Z(n2109) );
  HS65_LH_AO22X9 U2065 ( .A(n6287), .B(\registers[22][4] ), .C(
        \regfile_i[WRITE_DATA][4] ), .D(n6291), .Z(n2110) );
  HS65_LH_AO22X9 U2066 ( .A(n6287), .B(\registers[22][5] ), .C(
        \regfile_i[WRITE_DATA][5] ), .D(n6291), .Z(n2111) );
  HS65_LH_AO22X9 U2067 ( .A(n6287), .B(\registers[22][6] ), .C(
        \regfile_i[WRITE_DATA][6] ), .D(n6291), .Z(n2112) );
  HS65_LH_AO22X9 U2068 ( .A(n6287), .B(\registers[22][7] ), .C(
        \regfile_i[WRITE_DATA][7] ), .D(n6291), .Z(n2113) );
  HS65_LH_AO22X9 U2069 ( .A(n6287), .B(\registers[22][8] ), .C(
        \regfile_i[WRITE_DATA][8] ), .D(n6291), .Z(n2114) );
  HS65_LH_AO22X9 U2070 ( .A(n6287), .B(\registers[22][9] ), .C(
        \regfile_i[WRITE_DATA][9] ), .D(n6291), .Z(n2115) );
  HS65_LH_AO22X9 U2071 ( .A(n6287), .B(\registers[22][10] ), .C(
        \regfile_i[WRITE_DATA][10] ), .D(n6291), .Z(n2116) );
  HS65_LH_AO22X9 U2072 ( .A(n6287), .B(\registers[22][11] ), .C(
        \regfile_i[WRITE_DATA][11] ), .D(n6290), .Z(n2117) );
  HS65_LH_AO22X9 U2073 ( .A(n6288), .B(\registers[22][12] ), .C(
        \regfile_i[WRITE_DATA][12] ), .D(n6290), .Z(n2118) );
  HS65_LH_AO22X9 U2074 ( .A(n6288), .B(\registers[22][13] ), .C(
        \regfile_i[WRITE_DATA][13] ), .D(n6290), .Z(n2119) );
  HS65_LH_AO22X9 U2075 ( .A(n6288), .B(\registers[22][14] ), .C(
        \regfile_i[WRITE_DATA][14] ), .D(n6290), .Z(n2120) );
  HS65_LH_AO22X9 U2076 ( .A(n6288), .B(\registers[22][15] ), .C(
        \regfile_i[WRITE_DATA][15] ), .D(n6290), .Z(n2121) );
  HS65_LH_AO22X9 U2077 ( .A(n6288), .B(\registers[22][16] ), .C(
        \regfile_i[WRITE_DATA][16] ), .D(n6290), .Z(n2122) );
  HS65_LH_AO22X9 U2078 ( .A(n6288), .B(\registers[22][17] ), .C(
        \regfile_i[WRITE_DATA][17] ), .D(n6290), .Z(n2123) );
  HS65_LH_AO22X9 U2079 ( .A(n6288), .B(\registers[22][18] ), .C(
        \regfile_i[WRITE_DATA][18] ), .D(n6290), .Z(n2124) );
  HS65_LH_AO22X9 U2080 ( .A(n6288), .B(\registers[22][19] ), .C(
        \regfile_i[WRITE_DATA][19] ), .D(n6290), .Z(n2125) );
  HS65_LH_AO22X9 U2081 ( .A(n6288), .B(\registers[22][20] ), .C(
        \regfile_i[WRITE_DATA][20] ), .D(n6290), .Z(n2126) );
  HS65_LH_AO22X9 U2082 ( .A(n6288), .B(\registers[22][21] ), .C(
        \regfile_i[WRITE_DATA][21] ), .D(n6290), .Z(n2127) );
  HS65_LH_AO22X9 U2083 ( .A(n6288), .B(\registers[22][22] ), .C(
        \regfile_i[WRITE_DATA][22] ), .D(n6290), .Z(n2128) );
  HS65_LH_AO22X9 U2084 ( .A(n6288), .B(\registers[22][23] ), .C(
        \regfile_i[WRITE_DATA][23] ), .D(n6290), .Z(n2129) );
  HS65_LH_AO22X9 U2085 ( .A(n6287), .B(\registers[22][24] ), .C(
        \regfile_i[WRITE_DATA][24] ), .D(n6290), .Z(n2130) );
  HS65_LH_AO22X9 U2086 ( .A(n6288), .B(\registers[22][25] ), .C(
        \regfile_i[WRITE_DATA][25] ), .D(n6290), .Z(n2131) );
  HS65_LH_AO22X9 U2087 ( .A(n6287), .B(\registers[22][26] ), .C(
        \regfile_i[WRITE_DATA][26] ), .D(n6290), .Z(n2132) );
  HS65_LH_AO22X9 U2088 ( .A(n6288), .B(\registers[22][27] ), .C(
        \regfile_i[WRITE_DATA][27] ), .D(n6290), .Z(n2133) );
  HS65_LH_AO22X9 U2089 ( .A(n6287), .B(\registers[22][28] ), .C(
        \regfile_i[WRITE_DATA][28] ), .D(n6290), .Z(n2134) );
  HS65_LH_AO22X9 U2090 ( .A(n6288), .B(\registers[22][29] ), .C(
        \regfile_i[WRITE_DATA][29] ), .D(n6290), .Z(n2135) );
  HS65_LH_AO22X9 U2091 ( .A(n6287), .B(\registers[22][30] ), .C(
        \regfile_i[WRITE_DATA][30] ), .D(n6290), .Z(n2136) );
  HS65_LH_AO22X9 U2092 ( .A(n6288), .B(\registers[22][31] ), .C(
        \regfile_i[WRITE_DATA][31] ), .D(n6289), .Z(n2137) );
  HS65_LH_NOR3X4 U2093 ( .A(\regfile_i[ADRWRITE][1] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(n814), .Z(n2837) );
  HS65_LH_NOR3X4 U2094 ( .A(\regfile_i[ADRWRITE][0] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(n813), .Z(n2835) );
  HS65_LH_NOR3X4 U2095 ( .A(n814), .B(\regfile_i[ADRWRITE][2] ), .C(n813), .Z(
        n2833) );
  HS65_LH_NOR3X4 U2096 ( .A(\regfile_i[ADRWRITE][0] ), .B(
        \regfile_i[ADRWRITE][1] ), .C(n812), .Z(n2831) );
  HS65_LH_NOR3X4 U2097 ( .A(n814), .B(\regfile_i[ADRWRITE][1] ), .C(n812), .Z(
        n2829) );
  HS65_LH_NOR3X4 U2098 ( .A(n813), .B(\regfile_i[ADRWRITE][0] ), .C(n812), .Z(
        n2827) );
  HS65_LH_NOR3X4 U2099 ( .A(n770), .B(\regfile_i[ADRREAD0][4] ), .C(n773), .Z(
        n2805) );
  HS65_LH_NOR3X4 U2100 ( .A(\regfile_i[ADRREAD0][0] ), .B(
        \regfile_i[ADRREAD0][3] ), .C(n769), .Z(n2822) );
  HS65_LH_NOR3X4 U2101 ( .A(\regfile_i[ADRREAD1][0] ), .B(
        \regfile_i[ADRREAD1][4] ), .C(n775), .Z(n1324) );
  HS65_LH_NOR3X4 U2102 ( .A(n774), .B(\regfile_i[ADRREAD1][3] ), .C(n778), .Z(
        n1331) );
  HS65_LH_NOR3X4 U2103 ( .A(n770), .B(\regfile_i[ADRREAD0][0] ), .C(n769), .Z(
        n2809) );
  HS65_LH_NOR3X4 U2104 ( .A(\regfile_i[ADRWRITE][1] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(\regfile_i[ADRWRITE][0] ), .Z(n2839) );
  HS65_LH_NOR3X4 U2105 ( .A(\regfile_i[ADRREAD1][0] ), .B(
        \regfile_i[ADRREAD1][3] ), .C(n774), .Z(n1337) );
  HS65_LH_NOR3X4 U2106 ( .A(\regfile_i[ADRREAD1][3] ), .B(
        \regfile_i[ADRREAD1][4] ), .C(n778), .Z(n1329) );
  HS65_LH_NOR3X4 U2107 ( .A(n775), .B(\regfile_i[ADRREAD1][4] ), .C(n778), .Z(
        n1326) );
  HS65_LH_NOR3X4 U2108 ( .A(\regfile_i[ADRREAD0][3] ), .B(
        \regfile_i[ADRREAD0][4] ), .C(n773), .Z(n2813) );
  HS65_LH_NOR3X4 U2109 ( .A(\regfile_i[ADRREAD0][0] ), .B(
        \regfile_i[ADRREAD0][4] ), .C(n770), .Z(n2811) );
  HS65_LH_NOR3X4 U2110 ( .A(n774), .B(\regfile_i[ADRREAD1][0] ), .C(n775), .Z(
        n1338) );
  HS65_LH_NOR3X4 U2111 ( .A(n769), .B(\regfile_i[ADRREAD0][3] ), .C(n773), .Z(
        n2820) );
  HS65_LH_NOR2X6 U2112 ( .A(\regfile_i[ADRREAD0][1] ), .B(
        \regfile_i[ADRREAD0][2] ), .Z(n2807) );
  HS65_LH_AOI222X2 U2113 ( .A(n6508), .B(n704), .C(\registers[4][0] ), .D(
        n6505), .E(\registers[1][0] ), .F(n6502), .Z(n1319) );
  HS65_LH_AOI222X2 U2114 ( .A(n6508), .B(n703), .C(\registers[4][1] ), .D(
        n6505), .E(\registers[1][1] ), .F(n6502), .Z(n1165) );
  HS65_LH_AOI222X2 U2115 ( .A(n6509), .B(n702), .C(\registers[4][2] ), .D(
        n6506), .E(\registers[1][2] ), .F(n6503), .Z(n1011) );
  HS65_LH_AOI222X2 U2116 ( .A(n6510), .B(n701), .C(\registers[4][3] ), .D(
        n6507), .E(\registers[1][3] ), .F(n6504), .Z(n969) );
  HS65_LH_AOI222X2 U2117 ( .A(n6510), .B(n700), .C(\registers[4][4] ), .D(
        n6507), .E(\registers[1][4] ), .F(n6504), .Z(n955) );
  HS65_LH_AOI222X2 U2118 ( .A(n6510), .B(n699), .C(\registers[4][5] ), .D(
        n6507), .E(\registers[1][5] ), .F(n6504), .Z(n941) );
  HS65_LH_AOI222X2 U2119 ( .A(n6510), .B(n698), .C(\registers[4][6] ), .D(
        n6507), .E(\registers[1][6] ), .F(n6504), .Z(n927) );
  HS65_LH_AOI222X2 U2120 ( .A(n6510), .B(n697), .C(\registers[4][7] ), .D(
        n6507), .E(\registers[1][7] ), .F(n6504), .Z(n913) );
  HS65_LH_AOI222X2 U2121 ( .A(n6510), .B(n696), .C(\registers[4][8] ), .D(
        n6507), .E(\registers[1][8] ), .F(n6504), .Z(n899) );
  HS65_LH_AOI222X2 U2122 ( .A(n6510), .B(n695), .C(\registers[4][9] ), .D(
        n6507), .E(\registers[1][9] ), .F(n6504), .Z(n854) );
  HS65_LH_AOI222X2 U2123 ( .A(n6508), .B(n694), .C(\registers[4][10] ), .D(
        n6505), .E(\registers[1][10] ), .F(n6502), .Z(n1305) );
  HS65_LH_AOI222X2 U2124 ( .A(n6508), .B(n693), .C(\registers[4][11] ), .D(
        n6505), .E(\registers[1][11] ), .F(n6502), .Z(n1291) );
  HS65_LH_AOI222X2 U2125 ( .A(n6508), .B(n692), .C(\registers[4][12] ), .D(
        n6505), .E(\registers[1][12] ), .F(n6502), .Z(n1277) );
  HS65_LH_AOI222X2 U2126 ( .A(n6508), .B(n691), .C(\registers[4][13] ), .D(
        n6505), .E(\registers[1][13] ), .F(n6502), .Z(n1263) );
  HS65_LH_AOI222X2 U2127 ( .A(n6508), .B(n690), .C(\registers[4][14] ), .D(
        n6505), .E(\registers[1][14] ), .F(n6502), .Z(n1249) );
  HS65_LH_AOI222X2 U2128 ( .A(n6508), .B(n689), .C(\registers[4][15] ), .D(
        n6505), .E(\registers[1][15] ), .F(n6502), .Z(n1235) );
  HS65_LH_AOI222X2 U2129 ( .A(n6508), .B(n688), .C(\registers[4][16] ), .D(
        n6505), .E(\registers[1][16] ), .F(n6502), .Z(n1221) );
  HS65_LH_AOI222X2 U2130 ( .A(n6508), .B(n687), .C(\registers[4][17] ), .D(
        n6505), .E(\registers[1][17] ), .F(n6502), .Z(n1207) );
  HS65_LH_AOI222X2 U2131 ( .A(n6508), .B(n686), .C(\registers[4][18] ), .D(
        n6505), .E(\registers[1][18] ), .F(n6502), .Z(n1193) );
  HS65_LH_AOI222X2 U2132 ( .A(n6508), .B(n685), .C(\registers[4][19] ), .D(
        n6505), .E(\registers[1][19] ), .F(n6502), .Z(n1179) );
  HS65_LH_AOI222X2 U2133 ( .A(n6509), .B(n684), .C(\registers[4][20] ), .D(
        n6506), .E(\registers[1][20] ), .F(n6503), .Z(n1151) );
  HS65_LH_AOI222X2 U2134 ( .A(n6509), .B(n683), .C(\registers[4][21] ), .D(
        n6506), .E(\registers[1][21] ), .F(n6503), .Z(n1137) );
  HS65_LH_AOI222X2 U2135 ( .A(n6509), .B(n682), .C(\registers[4][22] ), .D(
        n6506), .E(\registers[1][22] ), .F(n6503), .Z(n1123) );
  HS65_LH_AOI222X2 U2136 ( .A(n6509), .B(n681), .C(\registers[4][23] ), .D(
        n6506), .E(\registers[1][23] ), .F(n6503), .Z(n1109) );
  HS65_LH_AOI222X2 U2137 ( .A(n6509), .B(n680), .C(\registers[4][24] ), .D(
        n6506), .E(\registers[1][24] ), .F(n6503), .Z(n1095) );
  HS65_LH_AOI222X2 U2138 ( .A(n6509), .B(n679), .C(\registers[4][25] ), .D(
        n6506), .E(\registers[1][25] ), .F(n6503), .Z(n1081) );
  HS65_LH_AOI222X2 U2139 ( .A(n6509), .B(n678), .C(\registers[4][26] ), .D(
        n6506), .E(\registers[1][26] ), .F(n6503), .Z(n1067) );
  HS65_LH_AOI222X2 U2140 ( .A(n6509), .B(n677), .C(\registers[4][27] ), .D(
        n6506), .E(\registers[1][27] ), .F(n6503), .Z(n1053) );
  HS65_LH_AOI222X2 U2141 ( .A(n6509), .B(n676), .C(\registers[4][28] ), .D(
        n6506), .E(\registers[1][28] ), .F(n6503), .Z(n1039) );
  HS65_LH_AOI222X2 U2142 ( .A(n6509), .B(n675), .C(\registers[4][29] ), .D(
        n6506), .E(\registers[1][29] ), .F(n6503), .Z(n1025) );
  HS65_LH_AOI222X2 U2143 ( .A(n6509), .B(n674), .C(\registers[4][30] ), .D(
        n6506), .E(\registers[1][30] ), .F(n6503), .Z(n997) );
  HS65_LH_AOI222X2 U2144 ( .A(n6510), .B(n673), .C(\registers[4][31] ), .D(
        n6507), .E(\registers[1][31] ), .F(n6504), .Z(n983) );
  HS65_LH_NOR2X6 U2145 ( .A(n776), .B(\regfile_i[ADRREAD1][1] ), .Z(n1327) );
  HS65_LH_NOR2X6 U2146 ( .A(n772), .B(\regfile_i[ADRREAD0][2] ), .Z(n2808) );
  HS65_LH_NOR2X6 U2147 ( .A(\regfile_i[ADRREAD1][1] ), .B(
        \regfile_i[ADRREAD1][2] ), .Z(n1328) );
  HS65_LH_AOI222X2 U2148 ( .A(n6415), .B(\registers[13][0] ), .C(n6412), .D(
        \registers[10][0] ), .E(n6409), .F(\registers[6][0] ), .Z(n2802) );
  HS65_LH_AOI222X2 U2149 ( .A(n6415), .B(\registers[13][1] ), .C(n6412), .D(
        \registers[10][1] ), .E(n6409), .F(\registers[6][1] ), .Z(n2648) );
  HS65_LH_AOI222X2 U2150 ( .A(n6416), .B(\registers[13][2] ), .C(n6413), .D(
        \registers[10][2] ), .E(n6410), .F(\registers[6][2] ), .Z(n2494) );
  HS65_LH_AOI222X2 U2151 ( .A(n6417), .B(\registers[13][3] ), .C(n6414), .D(
        \registers[10][3] ), .E(n6410), .F(\registers[6][3] ), .Z(n2452) );
  HS65_LH_AOI222X2 U2152 ( .A(n6415), .B(\registers[13][10] ), .C(n6412), .D(
        \registers[10][10] ), .E(n6409), .F(\registers[6][10] ), .Z(n2788) );
  HS65_LH_AOI222X2 U2153 ( .A(n6415), .B(\registers[13][11] ), .C(n6412), .D(
        \registers[10][11] ), .E(n6409), .F(\registers[6][11] ), .Z(n2774) );
  HS65_LH_AOI222X2 U2154 ( .A(n6415), .B(\registers[13][12] ), .C(n6412), .D(
        \registers[10][12] ), .E(n6409), .F(\registers[6][12] ), .Z(n2760) );
  HS65_LH_AOI222X2 U2155 ( .A(n6415), .B(\registers[13][13] ), .C(n6412), .D(
        \registers[10][13] ), .E(n6409), .F(\registers[6][13] ), .Z(n2746) );
  HS65_LH_AOI222X2 U2156 ( .A(n6415), .B(\registers[13][14] ), .C(n6412), .D(
        \registers[10][14] ), .E(n6409), .F(\registers[6][14] ), .Z(n2732) );
  HS65_LH_AOI222X2 U2157 ( .A(n6415), .B(\registers[13][15] ), .C(n6412), .D(
        \registers[10][15] ), .E(n6409), .F(\registers[6][15] ), .Z(n2718) );
  HS65_LH_AOI222X2 U2158 ( .A(n6415), .B(\registers[13][16] ), .C(n6412), .D(
        \registers[10][16] ), .E(n6409), .F(\registers[6][16] ), .Z(n2704) );
  HS65_LH_AOI222X2 U2159 ( .A(n6415), .B(\registers[13][17] ), .C(n6412), .D(
        \registers[10][17] ), .E(n6409), .F(\registers[6][17] ), .Z(n2690) );
  HS65_LH_AOI222X2 U2160 ( .A(n6415), .B(\registers[13][18] ), .C(n6412), .D(
        \registers[10][18] ), .E(n6409), .F(\registers[6][18] ), .Z(n2676) );
  HS65_LH_AOI222X2 U2161 ( .A(n6415), .B(\registers[13][19] ), .C(n6412), .D(
        \registers[10][19] ), .E(n6409), .F(\registers[6][19] ), .Z(n2662) );
  HS65_LH_AOI222X2 U2162 ( .A(n6416), .B(\registers[13][20] ), .C(n6413), .D(
        \registers[10][20] ), .E(n6409), .F(\registers[6][20] ), .Z(n2634) );
  HS65_LH_AOI222X2 U2163 ( .A(n6416), .B(\registers[13][21] ), .C(n6413), .D(
        \registers[10][21] ), .E(n6410), .F(\registers[6][21] ), .Z(n2620) );
  HS65_LH_AOI222X2 U2164 ( .A(n6416), .B(\registers[13][22] ), .C(n6413), .D(
        \registers[10][22] ), .E(n6410), .F(\registers[6][22] ), .Z(n2606) );
  HS65_LH_AOI222X2 U2165 ( .A(n6416), .B(\registers[13][23] ), .C(n6413), .D(
        \registers[10][23] ), .E(n6410), .F(\registers[6][23] ), .Z(n2592) );
  HS65_LH_AOI222X2 U2166 ( .A(n6416), .B(\registers[13][24] ), .C(n6413), .D(
        \registers[10][24] ), .E(n6410), .F(\registers[6][24] ), .Z(n2578) );
  HS65_LH_AOI222X2 U2167 ( .A(n6416), .B(\registers[13][25] ), .C(n6413), .D(
        \registers[10][25] ), .E(n6410), .F(\registers[6][25] ), .Z(n2564) );
  HS65_LH_AOI222X2 U2168 ( .A(n6416), .B(\registers[13][26] ), .C(n6413), .D(
        \registers[10][26] ), .E(n6410), .F(\registers[6][26] ), .Z(n2550) );
  HS65_LH_AOI222X2 U2169 ( .A(n6416), .B(\registers[13][27] ), .C(n6413), .D(
        \registers[10][27] ), .E(n6410), .F(\registers[6][27] ), .Z(n2536) );
  HS65_LH_AOI222X2 U2170 ( .A(n6416), .B(\registers[13][28] ), .C(n6413), .D(
        \registers[10][28] ), .E(n6410), .F(\registers[6][28] ), .Z(n2522) );
  HS65_LH_AOI222X2 U2171 ( .A(n6416), .B(\registers[13][29] ), .C(n6413), .D(
        \registers[10][29] ), .E(n6410), .F(\registers[6][29] ), .Z(n2508) );
  HS65_LH_AOI222X2 U2172 ( .A(n6416), .B(\registers[13][30] ), .C(n6413), .D(
        \registers[10][30] ), .E(n6410), .F(\registers[6][30] ), .Z(n2480) );
  HS65_LH_AOI222X2 U2173 ( .A(n6417), .B(\registers[13][31] ), .C(n6414), .D(
        \registers[10][31] ), .E(n6410), .F(\registers[6][31] ), .Z(n2466) );
  HS65_LH_AOI222X2 U2174 ( .A(n6417), .B(\registers[13][4] ), .C(n6414), .D(
        \registers[10][4] ), .E(n6411), .F(\registers[6][4] ), .Z(n2438) );
  HS65_LH_AOI222X2 U2175 ( .A(n6417), .B(\registers[13][5] ), .C(n6414), .D(
        \registers[10][5] ), .E(n6411), .F(\registers[6][5] ), .Z(n1432) );
  HS65_LH_AOI222X2 U2176 ( .A(n6417), .B(\registers[13][6] ), .C(n6414), .D(
        \registers[10][6] ), .E(n6411), .F(\registers[6][6] ), .Z(n1418) );
  HS65_LH_AOI222X2 U2177 ( .A(n6417), .B(\registers[13][7] ), .C(n6414), .D(
        \registers[10][7] ), .E(n6411), .F(\registers[6][7] ), .Z(n1404) );
  HS65_LH_AOI222X2 U2178 ( .A(n6417), .B(\registers[13][8] ), .C(n6414), .D(
        \registers[10][8] ), .E(n6411), .F(\registers[6][8] ), .Z(n1390) );
  HS65_LH_AOI222X2 U2179 ( .A(n6417), .B(\registers[13][9] ), .C(n6414), .D(
        \registers[10][9] ), .E(n6411), .F(\registers[6][9] ), .Z(n1345) );
  HS65_LH_NOR2X6 U2180 ( .A(n777), .B(\regfile_i[ADRREAD1][2] ), .Z(n1325) );
  HS65_LH_AOI212X4 U2181 ( .A(n6463), .B(n544), .C(\registers[31][0] ), .D(
        n6460), .E(n1339), .Z(n1334) );
  HS65_LH_OAI22X6 U2182 ( .A(n6457), .B(n288), .C(n6454), .D(n448), .Z(n1339)
         );
  HS65_LH_AOI212X4 U2183 ( .A(n6463), .B(n543), .C(\registers[31][1] ), .D(
        n6460), .E(n1173), .Z(n1170) );
  HS65_LH_OAI22X6 U2184 ( .A(n6457), .B(n287), .C(n6454), .D(n447), .Z(n1173)
         );
  HS65_LH_AOI212X4 U2185 ( .A(n6464), .B(n542), .C(\registers[31][2] ), .D(
        n6461), .E(n1019), .Z(n1016) );
  HS65_LH_OAI22X6 U2186 ( .A(n6458), .B(n286), .C(n6455), .D(n446), .Z(n1019)
         );
  HS65_LH_AOI212X4 U2187 ( .A(n6464), .B(n541), .C(\registers[31][3] ), .D(
        n6461), .E(n977), .Z(n974) );
  HS65_LH_OAI22X6 U2188 ( .A(n6459), .B(n285), .C(n6455), .D(n445), .Z(n977)
         );
  HS65_LH_AOI212X4 U2189 ( .A(n6465), .B(n540), .C(\registers[31][4] ), .D(
        n6462), .E(n963), .Z(n960) );
  HS65_LH_OAI22X6 U2190 ( .A(n6459), .B(n284), .C(n6456), .D(n444), .Z(n963)
         );
  HS65_LH_AOI212X4 U2191 ( .A(n6465), .B(n539), .C(\registers[31][5] ), .D(
        n6462), .E(n949), .Z(n946) );
  HS65_LH_OAI22X6 U2192 ( .A(n6459), .B(n283), .C(n6456), .D(n443), .Z(n949)
         );
  HS65_LH_AOI212X4 U2193 ( .A(n6465), .B(n538), .C(\registers[31][6] ), .D(
        n6462), .E(n935), .Z(n932) );
  HS65_LH_OAI22X6 U2194 ( .A(n6459), .B(n282), .C(n6456), .D(n442), .Z(n935)
         );
  HS65_LH_AOI212X4 U2195 ( .A(n6465), .B(n537), .C(\registers[31][7] ), .D(
        n6462), .E(n921), .Z(n918) );
  HS65_LH_OAI22X6 U2196 ( .A(n6459), .B(n281), .C(n6456), .D(n441), .Z(n921)
         );
  HS65_LH_AOI212X4 U2197 ( .A(n6465), .B(n536), .C(\registers[31][8] ), .D(
        n6462), .E(n907), .Z(n904) );
  HS65_LH_OAI22X6 U2198 ( .A(n6459), .B(n280), .C(n6456), .D(n440), .Z(n907)
         );
  HS65_LH_AOI212X4 U2199 ( .A(n6465), .B(n535), .C(\registers[31][9] ), .D(
        n6462), .E(n883), .Z(n874) );
  HS65_LH_OAI22X6 U2200 ( .A(n6459), .B(n279), .C(n6456), .D(n439), .Z(n883)
         );
  HS65_LH_AOI212X4 U2201 ( .A(n6463), .B(n534), .C(\registers[31][10] ), .D(
        n6460), .E(n1313), .Z(n1310) );
  HS65_LH_OAI22X6 U2202 ( .A(n6457), .B(n278), .C(n6454), .D(n438), .Z(n1313)
         );
  HS65_LH_AOI212X4 U2203 ( .A(n6463), .B(n533), .C(\registers[31][11] ), .D(
        n6460), .E(n1299), .Z(n1296) );
  HS65_LH_OAI22X6 U2204 ( .A(n6457), .B(n277), .C(n6454), .D(n437), .Z(n1299)
         );
  HS65_LH_AOI212X4 U2205 ( .A(n6463), .B(n532), .C(\registers[31][12] ), .D(
        n6460), .E(n1285), .Z(n1282) );
  HS65_LH_OAI22X6 U2206 ( .A(n6457), .B(n276), .C(n6454), .D(n436), .Z(n1285)
         );
  HS65_LH_AOI212X4 U2207 ( .A(n6463), .B(n531), .C(\registers[31][13] ), .D(
        n6460), .E(n1271), .Z(n1268) );
  HS65_LH_OAI22X6 U2208 ( .A(n6457), .B(n275), .C(n6454), .D(n435), .Z(n1271)
         );
  HS65_LH_AOI212X4 U2209 ( .A(n6463), .B(n530), .C(\registers[31][14] ), .D(
        n6460), .E(n1257), .Z(n1254) );
  HS65_LH_OAI22X6 U2210 ( .A(n6457), .B(n274), .C(n6454), .D(n434), .Z(n1257)
         );
  HS65_LH_AOI212X4 U2211 ( .A(n6463), .B(n529), .C(\registers[31][15] ), .D(
        n6460), .E(n1243), .Z(n1240) );
  HS65_LH_OAI22X6 U2212 ( .A(n6457), .B(n273), .C(n6454), .D(n433), .Z(n1243)
         );
  HS65_LH_AOI212X4 U2213 ( .A(n6463), .B(n528), .C(\registers[31][16] ), .D(
        n6460), .E(n1229), .Z(n1226) );
  HS65_LH_OAI22X6 U2214 ( .A(n6457), .B(n272), .C(n6454), .D(n432), .Z(n1229)
         );
  HS65_LH_AOI212X4 U2215 ( .A(n6463), .B(n527), .C(\registers[31][17] ), .D(
        n6460), .E(n1215), .Z(n1212) );
  HS65_LH_OAI22X6 U2216 ( .A(n6457), .B(n271), .C(n6454), .D(n431), .Z(n1215)
         );
  HS65_LH_AOI212X4 U2217 ( .A(n6463), .B(n526), .C(\registers[31][18] ), .D(
        n6460), .E(n1201), .Z(n1198) );
  HS65_LH_OAI22X6 U2218 ( .A(n6457), .B(n270), .C(n6454), .D(n430), .Z(n1201)
         );
  HS65_LH_AOI212X4 U2219 ( .A(n6463), .B(n525), .C(\registers[31][19] ), .D(
        n6460), .E(n1187), .Z(n1184) );
  HS65_LH_OAI22X6 U2220 ( .A(n6457), .B(n269), .C(n6454), .D(n429), .Z(n1187)
         );
  HS65_LH_AOI212X4 U2221 ( .A(n6463), .B(n524), .C(\registers[31][20] ), .D(
        n6460), .E(n1159), .Z(n1156) );
  HS65_LH_OAI22X6 U2222 ( .A(n6458), .B(n268), .C(n6454), .D(n428), .Z(n1159)
         );
  HS65_LH_AOI212X4 U2223 ( .A(n6464), .B(n523), .C(\registers[31][21] ), .D(
        n6461), .E(n1145), .Z(n1142) );
  HS65_LH_OAI22X6 U2224 ( .A(n6458), .B(n267), .C(n6455), .D(n427), .Z(n1145)
         );
  HS65_LH_AOI212X4 U2225 ( .A(n6464), .B(n522), .C(\registers[31][22] ), .D(
        n6461), .E(n1131), .Z(n1128) );
  HS65_LH_OAI22X6 U2226 ( .A(n6458), .B(n266), .C(n6455), .D(n426), .Z(n1131)
         );
  HS65_LH_AOI212X4 U2227 ( .A(n6464), .B(n521), .C(\registers[31][23] ), .D(
        n6461), .E(n1117), .Z(n1114) );
  HS65_LH_OAI22X6 U2228 ( .A(n6458), .B(n265), .C(n6455), .D(n425), .Z(n1117)
         );
  HS65_LH_AOI212X4 U2229 ( .A(n6464), .B(n520), .C(\registers[31][24] ), .D(
        n6461), .E(n1103), .Z(n1100) );
  HS65_LH_OAI22X6 U2230 ( .A(n6458), .B(n264), .C(n6455), .D(n424), .Z(n1103)
         );
  HS65_LH_AOI212X4 U2231 ( .A(n6464), .B(n519), .C(\registers[31][25] ), .D(
        n6461), .E(n1089), .Z(n1086) );
  HS65_LH_OAI22X6 U2232 ( .A(n6458), .B(n263), .C(n6455), .D(n423), .Z(n1089)
         );
  HS65_LH_AOI212X4 U2233 ( .A(n6464), .B(n518), .C(\registers[31][26] ), .D(
        n6461), .E(n1075), .Z(n1072) );
  HS65_LH_OAI22X6 U2234 ( .A(n6458), .B(n262), .C(n6455), .D(n422), .Z(n1075)
         );
  HS65_LH_AOI212X4 U2235 ( .A(n6464), .B(n517), .C(\registers[31][27] ), .D(
        n6461), .E(n1061), .Z(n1058) );
  HS65_LH_OAI22X6 U2236 ( .A(n6458), .B(n261), .C(n6455), .D(n421), .Z(n1061)
         );
  HS65_LH_AOI212X4 U2237 ( .A(n6464), .B(n516), .C(\registers[31][28] ), .D(
        n6461), .E(n1047), .Z(n1044) );
  HS65_LH_OAI22X6 U2238 ( .A(n6458), .B(n260), .C(n6455), .D(n420), .Z(n1047)
         );
  HS65_LH_AOI212X4 U2239 ( .A(n6464), .B(n515), .C(\registers[31][29] ), .D(
        n6461), .E(n1033), .Z(n1030) );
  HS65_LH_OAI22X6 U2240 ( .A(n6458), .B(n259), .C(n6455), .D(n419), .Z(n1033)
         );
  HS65_LH_AOI212X4 U2241 ( .A(n6464), .B(n514), .C(\registers[31][30] ), .D(
        n6461), .E(n1005), .Z(n1002) );
  HS65_LH_OAI22X6 U2242 ( .A(n6458), .B(n258), .C(n6455), .D(n418), .Z(n1005)
         );
  HS65_LH_AOI212X4 U2243 ( .A(n6464), .B(n513), .C(\registers[31][31] ), .D(
        n6461), .E(n991), .Z(n988) );
  HS65_LH_OAI22X6 U2244 ( .A(n6459), .B(n257), .C(n6455), .D(n417), .Z(n991)
         );
  HS65_LH_AOI212X4 U2245 ( .A(n6520), .B(n736), .C(\registers[13][0] ), .D(
        n6517), .E(n1321), .Z(n1320) );
  HS65_LH_IVX9 U2246 ( .A(n224), .Z(n736) );
  HS65_LH_OAI22X6 U2247 ( .A(n6514), .B(n480), .C(n6511), .D(n512), .Z(n1321)
         );
  HS65_LH_AOI212X4 U2248 ( .A(n6520), .B(n735), .C(\registers[13][1] ), .D(
        n6517), .E(n1167), .Z(n1166) );
  HS65_LH_IVX9 U2249 ( .A(n223), .Z(n735) );
  HS65_LH_OAI22X6 U2250 ( .A(n6514), .B(n479), .C(n6511), .D(n511), .Z(n1167)
         );
  HS65_LH_AOI212X4 U2251 ( .A(n6521), .B(n734), .C(\registers[13][2] ), .D(
        n6518), .E(n1013), .Z(n1012) );
  HS65_LH_IVX9 U2252 ( .A(n222), .Z(n734) );
  HS65_LH_OAI22X6 U2253 ( .A(n6515), .B(n478), .C(n6512), .D(n510), .Z(n1013)
         );
  HS65_LH_AOI212X4 U2254 ( .A(n6521), .B(n733), .C(\registers[13][3] ), .D(
        n6518), .E(n971), .Z(n970) );
  HS65_LH_IVX9 U2255 ( .A(n221), .Z(n733) );
  HS65_LH_OAI22X6 U2256 ( .A(n6516), .B(n477), .C(n6512), .D(n509), .Z(n971)
         );
  HS65_LH_AOI212X4 U2257 ( .A(n6522), .B(n732), .C(\registers[13][4] ), .D(
        n6519), .E(n957), .Z(n956) );
  HS65_LH_IVX9 U2258 ( .A(n220), .Z(n732) );
  HS65_LH_OAI22X6 U2259 ( .A(n6516), .B(n476), .C(n6513), .D(n508), .Z(n957)
         );
  HS65_LH_AOI212X4 U2260 ( .A(n6522), .B(n731), .C(\registers[13][5] ), .D(
        n6519), .E(n943), .Z(n942) );
  HS65_LH_IVX9 U2261 ( .A(n219), .Z(n731) );
  HS65_LH_OAI22X6 U2262 ( .A(n6516), .B(n475), .C(n6513), .D(n507), .Z(n943)
         );
  HS65_LH_AOI212X4 U2263 ( .A(n6522), .B(n730), .C(\registers[13][6] ), .D(
        n6519), .E(n929), .Z(n928) );
  HS65_LH_IVX9 U2264 ( .A(n218), .Z(n730) );
  HS65_LH_OAI22X6 U2265 ( .A(n6516), .B(n474), .C(n6513), .D(n506), .Z(n929)
         );
  HS65_LH_AOI212X4 U2266 ( .A(n6522), .B(n729), .C(\registers[13][7] ), .D(
        n6519), .E(n915), .Z(n914) );
  HS65_LH_IVX9 U2267 ( .A(n217), .Z(n729) );
  HS65_LH_OAI22X6 U2268 ( .A(n6516), .B(n473), .C(n6513), .D(n505), .Z(n915)
         );
  HS65_LH_AOI212X4 U2269 ( .A(n6522), .B(n728), .C(\registers[13][8] ), .D(
        n6519), .E(n901), .Z(n900) );
  HS65_LH_IVX9 U2270 ( .A(n216), .Z(n728) );
  HS65_LH_OAI22X6 U2271 ( .A(n6516), .B(n472), .C(n6513), .D(n504), .Z(n901)
         );
  HS65_LH_AOI212X4 U2272 ( .A(n6522), .B(n727), .C(\registers[13][9] ), .D(
        n6519), .E(n858), .Z(n855) );
  HS65_LH_IVX9 U2273 ( .A(n215), .Z(n727) );
  HS65_LH_OAI22X6 U2274 ( .A(n6516), .B(n471), .C(n6513), .D(n503), .Z(n858)
         );
  HS65_LH_AOI212X4 U2275 ( .A(n6520), .B(n726), .C(\registers[13][10] ), .D(
        n6517), .E(n1307), .Z(n1306) );
  HS65_LH_IVX9 U2276 ( .A(n214), .Z(n726) );
  HS65_LH_OAI22X6 U2277 ( .A(n6514), .B(n470), .C(n6511), .D(n502), .Z(n1307)
         );
  HS65_LH_AOI212X4 U2278 ( .A(n6520), .B(n725), .C(\registers[13][11] ), .D(
        n6517), .E(n1293), .Z(n1292) );
  HS65_LH_IVX9 U2279 ( .A(n213), .Z(n725) );
  HS65_LH_OAI22X6 U2280 ( .A(n6514), .B(n469), .C(n6511), .D(n501), .Z(n1293)
         );
  HS65_LH_AOI212X4 U2281 ( .A(n6520), .B(n724), .C(\registers[13][12] ), .D(
        n6517), .E(n1279), .Z(n1278) );
  HS65_LH_IVX9 U2282 ( .A(n212), .Z(n724) );
  HS65_LH_OAI22X6 U2283 ( .A(n6514), .B(n468), .C(n6511), .D(n500), .Z(n1279)
         );
  HS65_LH_AOI212X4 U2284 ( .A(n6520), .B(n723), .C(\registers[13][13] ), .D(
        n6517), .E(n1265), .Z(n1264) );
  HS65_LH_IVX9 U2285 ( .A(n211), .Z(n723) );
  HS65_LH_OAI22X6 U2286 ( .A(n6514), .B(n467), .C(n6511), .D(n499), .Z(n1265)
         );
  HS65_LH_AOI212X4 U2287 ( .A(n6520), .B(n722), .C(\registers[13][14] ), .D(
        n6517), .E(n1251), .Z(n1250) );
  HS65_LH_IVX9 U2288 ( .A(n210), .Z(n722) );
  HS65_LH_OAI22X6 U2289 ( .A(n6514), .B(n466), .C(n6511), .D(n498), .Z(n1251)
         );
  HS65_LH_AOI212X4 U2290 ( .A(n6520), .B(n721), .C(\registers[13][15] ), .D(
        n6517), .E(n1237), .Z(n1236) );
  HS65_LH_IVX9 U2291 ( .A(n209), .Z(n721) );
  HS65_LH_OAI22X6 U2292 ( .A(n6514), .B(n465), .C(n6511), .D(n497), .Z(n1237)
         );
  HS65_LH_AOI212X4 U2293 ( .A(n6520), .B(n720), .C(\registers[13][16] ), .D(
        n6517), .E(n1223), .Z(n1222) );
  HS65_LH_IVX9 U2294 ( .A(n208), .Z(n720) );
  HS65_LH_OAI22X6 U2295 ( .A(n6514), .B(n464), .C(n6511), .D(n496), .Z(n1223)
         );
  HS65_LH_AOI212X4 U2296 ( .A(n6520), .B(n719), .C(\registers[13][17] ), .D(
        n6517), .E(n1209), .Z(n1208) );
  HS65_LH_IVX9 U2297 ( .A(n207), .Z(n719) );
  HS65_LH_OAI22X6 U2298 ( .A(n6514), .B(n463), .C(n6511), .D(n495), .Z(n1209)
         );
  HS65_LH_AOI212X4 U2299 ( .A(n6520), .B(n718), .C(\registers[13][18] ), .D(
        n6517), .E(n1195), .Z(n1194) );
  HS65_LH_IVX9 U2300 ( .A(n206), .Z(n718) );
  HS65_LH_OAI22X6 U2301 ( .A(n6514), .B(n462), .C(n6511), .D(n494), .Z(n1195)
         );
  HS65_LH_AOI212X4 U2302 ( .A(n6520), .B(n717), .C(\registers[13][19] ), .D(
        n6517), .E(n1181), .Z(n1180) );
  HS65_LH_IVX9 U2303 ( .A(n205), .Z(n717) );
  HS65_LH_OAI22X6 U2304 ( .A(n6514), .B(n461), .C(n6511), .D(n493), .Z(n1181)
         );
  HS65_LH_AOI212X4 U2305 ( .A(n6520), .B(n716), .C(\registers[13][20] ), .D(
        n6517), .E(n1153), .Z(n1152) );
  HS65_LH_IVX9 U2306 ( .A(n204), .Z(n716) );
  HS65_LH_OAI22X6 U2307 ( .A(n6515), .B(n460), .C(n6511), .D(n492), .Z(n1153)
         );
  HS65_LH_AOI212X4 U2308 ( .A(n6521), .B(n715), .C(\registers[13][21] ), .D(
        n6518), .E(n1139), .Z(n1138) );
  HS65_LH_IVX9 U2309 ( .A(n203), .Z(n715) );
  HS65_LH_OAI22X6 U2310 ( .A(n6515), .B(n459), .C(n6512), .D(n491), .Z(n1139)
         );
  HS65_LH_AOI212X4 U2311 ( .A(n6521), .B(n714), .C(\registers[13][22] ), .D(
        n6518), .E(n1125), .Z(n1124) );
  HS65_LH_IVX9 U2312 ( .A(n202), .Z(n714) );
  HS65_LH_OAI22X6 U2313 ( .A(n6515), .B(n458), .C(n6512), .D(n490), .Z(n1125)
         );
  HS65_LH_AOI212X4 U2314 ( .A(n6521), .B(n713), .C(\registers[13][23] ), .D(
        n6518), .E(n1111), .Z(n1110) );
  HS65_LH_IVX9 U2315 ( .A(n201), .Z(n713) );
  HS65_LH_OAI22X6 U2316 ( .A(n6515), .B(n457), .C(n6512), .D(n489), .Z(n1111)
         );
  HS65_LH_AOI212X4 U2317 ( .A(n6521), .B(n712), .C(\registers[13][24] ), .D(
        n6518), .E(n1097), .Z(n1096) );
  HS65_LH_IVX9 U2318 ( .A(n200), .Z(n712) );
  HS65_LH_OAI22X6 U2319 ( .A(n6515), .B(n456), .C(n6512), .D(n488), .Z(n1097)
         );
  HS65_LH_AOI212X4 U2320 ( .A(n6521), .B(n711), .C(\registers[13][25] ), .D(
        n6518), .E(n1083), .Z(n1082) );
  HS65_LH_IVX9 U2321 ( .A(n199), .Z(n711) );
  HS65_LH_OAI22X6 U2322 ( .A(n6515), .B(n455), .C(n6512), .D(n487), .Z(n1083)
         );
  HS65_LH_AOI212X4 U2323 ( .A(n6521), .B(n710), .C(\registers[13][26] ), .D(
        n6518), .E(n1069), .Z(n1068) );
  HS65_LH_IVX9 U2324 ( .A(n198), .Z(n710) );
  HS65_LH_OAI22X6 U2325 ( .A(n6515), .B(n454), .C(n6512), .D(n486), .Z(n1069)
         );
  HS65_LH_AOI212X4 U2326 ( .A(n6521), .B(n709), .C(\registers[13][27] ), .D(
        n6518), .E(n1055), .Z(n1054) );
  HS65_LH_IVX9 U2327 ( .A(n197), .Z(n709) );
  HS65_LH_OAI22X6 U2328 ( .A(n6515), .B(n453), .C(n6512), .D(n485), .Z(n1055)
         );
  HS65_LH_AOI212X4 U2329 ( .A(n6521), .B(n708), .C(\registers[13][28] ), .D(
        n6518), .E(n1041), .Z(n1040) );
  HS65_LH_IVX9 U2330 ( .A(n196), .Z(n708) );
  HS65_LH_OAI22X6 U2331 ( .A(n6515), .B(n452), .C(n6512), .D(n484), .Z(n1041)
         );
  HS65_LH_AOI212X4 U2332 ( .A(n6521), .B(n707), .C(\registers[13][29] ), .D(
        n6518), .E(n1027), .Z(n1026) );
  HS65_LH_IVX9 U2333 ( .A(n195), .Z(n707) );
  HS65_LH_OAI22X6 U2334 ( .A(n6515), .B(n451), .C(n6512), .D(n483), .Z(n1027)
         );
  HS65_LH_AOI212X4 U2335 ( .A(n6521), .B(n706), .C(\registers[13][30] ), .D(
        n6518), .E(n999), .Z(n998) );
  HS65_LH_IVX9 U2336 ( .A(n194), .Z(n706) );
  HS65_LH_OAI22X6 U2337 ( .A(n6515), .B(n450), .C(n6512), .D(n482), .Z(n999)
         );
  HS65_LH_AOI212X4 U2338 ( .A(n6521), .B(n705), .C(\registers[13][31] ), .D(
        n6518), .E(n985), .Z(n984) );
  HS65_LH_IVX9 U2339 ( .A(n193), .Z(n705) );
  HS65_LH_OAI22X6 U2340 ( .A(n6516), .B(n449), .C(n6512), .D(n481), .Z(n985)
         );
  HS65_LH_NOR3X4 U2341 ( .A(\regfile_i[ADRREAD1][3] ), .B(
        \regfile_i[ADRREAD1][4] ), .C(\regfile_i[ADRREAD1][0] ), .Z(n1322) );
  HS65_LH_AOI212X4 U2342 ( .A(\registers[18][0] ), .B(n6475), .C(
        \registers[24][0] ), .D(n6472), .E(n1336), .Z(n1335) );
  HS65_LH_OAI22X6 U2343 ( .A(n6469), .B(n416), .C(n6466), .D(n384), .Z(n1336)
         );
  HS65_LH_AOI212X4 U2344 ( .A(\registers[18][1] ), .B(n6475), .C(
        \registers[24][1] ), .D(n6472), .E(n1172), .Z(n1171) );
  HS65_LH_OAI22X6 U2345 ( .A(n6469), .B(n415), .C(n6466), .D(n383), .Z(n1172)
         );
  HS65_LH_AOI212X4 U2346 ( .A(\registers[18][2] ), .B(n6476), .C(
        \registers[24][2] ), .D(n6473), .E(n1018), .Z(n1017) );
  HS65_LH_OAI22X6 U2347 ( .A(n6470), .B(n414), .C(n6467), .D(n382), .Z(n1018)
         );
  HS65_LH_AOI212X4 U2348 ( .A(\registers[18][3] ), .B(n6477), .C(
        \registers[24][3] ), .D(n6473), .E(n976), .Z(n975) );
  HS65_LH_OAI22X6 U2349 ( .A(n6471), .B(n413), .C(n6467), .D(n381), .Z(n976)
         );
  HS65_LH_AOI212X4 U2350 ( .A(\registers[18][4] ), .B(n6477), .C(
        \registers[24][4] ), .D(n6474), .E(n962), .Z(n961) );
  HS65_LH_OAI22X6 U2351 ( .A(n6471), .B(n412), .C(n6468), .D(n380), .Z(n962)
         );
  HS65_LH_AOI212X4 U2352 ( .A(\registers[18][5] ), .B(n6477), .C(
        \registers[24][5] ), .D(n6474), .E(n948), .Z(n947) );
  HS65_LH_OAI22X6 U2353 ( .A(n6471), .B(n411), .C(n6468), .D(n379), .Z(n948)
         );
  HS65_LH_AOI212X4 U2354 ( .A(\registers[18][6] ), .B(n6477), .C(
        \registers[24][6] ), .D(n6474), .E(n934), .Z(n933) );
  HS65_LH_OAI22X6 U2355 ( .A(n6471), .B(n410), .C(n6468), .D(n378), .Z(n934)
         );
  HS65_LH_AOI212X4 U2356 ( .A(\registers[18][7] ), .B(n6477), .C(
        \registers[24][7] ), .D(n6474), .E(n920), .Z(n919) );
  HS65_LH_OAI22X6 U2357 ( .A(n6471), .B(n409), .C(n6468), .D(n377), .Z(n920)
         );
  HS65_LH_AOI212X4 U2358 ( .A(\registers[18][8] ), .B(n6477), .C(
        \registers[24][8] ), .D(n6474), .E(n906), .Z(n905) );
  HS65_LH_OAI22X6 U2359 ( .A(n6471), .B(n408), .C(n6468), .D(n376), .Z(n906)
         );
  HS65_LH_AOI212X4 U2360 ( .A(\registers[18][9] ), .B(n6477), .C(
        \registers[24][9] ), .D(n6474), .E(n878), .Z(n875) );
  HS65_LH_OAI22X6 U2361 ( .A(n6471), .B(n407), .C(n6468), .D(n375), .Z(n878)
         );
  HS65_LH_AOI212X4 U2362 ( .A(\registers[18][11] ), .B(n6475), .C(
        \registers[24][11] ), .D(n6472), .E(n1298), .Z(n1297) );
  HS65_LH_OAI22X6 U2363 ( .A(n6469), .B(n405), .C(n6466), .D(n373), .Z(n1298)
         );
  HS65_LH_AOI212X4 U2364 ( .A(\registers[18][12] ), .B(n6475), .C(
        \registers[24][12] ), .D(n6472), .E(n1284), .Z(n1283) );
  HS65_LH_OAI22X6 U2365 ( .A(n6469), .B(n404), .C(n6466), .D(n372), .Z(n1284)
         );
  HS65_LH_AOI212X4 U2366 ( .A(\registers[18][13] ), .B(n6475), .C(
        \registers[24][13] ), .D(n6472), .E(n1270), .Z(n1269) );
  HS65_LH_OAI22X6 U2367 ( .A(n6469), .B(n403), .C(n6466), .D(n371), .Z(n1270)
         );
  HS65_LH_AOI212X4 U2368 ( .A(\registers[18][14] ), .B(n6475), .C(
        \registers[24][14] ), .D(n6472), .E(n1256), .Z(n1255) );
  HS65_LH_OAI22X6 U2369 ( .A(n6469), .B(n402), .C(n6466), .D(n370), .Z(n1256)
         );
  HS65_LH_AOI212X4 U2370 ( .A(\registers[18][15] ), .B(n6475), .C(
        \registers[24][15] ), .D(n6472), .E(n1242), .Z(n1241) );
  HS65_LH_OAI22X6 U2371 ( .A(n6469), .B(n401), .C(n6466), .D(n369), .Z(n1242)
         );
  HS65_LH_AOI212X4 U2372 ( .A(\registers[18][16] ), .B(n6475), .C(
        \registers[24][16] ), .D(n6472), .E(n1228), .Z(n1227) );
  HS65_LH_OAI22X6 U2373 ( .A(n6469), .B(n400), .C(n6466), .D(n368), .Z(n1228)
         );
  HS65_LH_AOI212X4 U2374 ( .A(\registers[18][17] ), .B(n6475), .C(
        \registers[24][17] ), .D(n6472), .E(n1214), .Z(n1213) );
  HS65_LH_OAI22X6 U2375 ( .A(n6469), .B(n399), .C(n6466), .D(n367), .Z(n1214)
         );
  HS65_LH_AOI212X4 U2376 ( .A(\registers[18][18] ), .B(n6475), .C(
        \registers[24][18] ), .D(n6472), .E(n1200), .Z(n1199) );
  HS65_LH_OAI22X6 U2377 ( .A(n6469), .B(n398), .C(n6466), .D(n366), .Z(n1200)
         );
  HS65_LH_AOI212X4 U2378 ( .A(\registers[18][19] ), .B(n6475), .C(
        \registers[24][19] ), .D(n6472), .E(n1186), .Z(n1185) );
  HS65_LH_OAI22X6 U2379 ( .A(n6469), .B(n397), .C(n6466), .D(n365), .Z(n1186)
         );
  HS65_LH_AOI212X4 U2380 ( .A(\registers[18][20] ), .B(n6476), .C(
        \registers[24][20] ), .D(n6472), .E(n1158), .Z(n1157) );
  HS65_LH_OAI22X6 U2381 ( .A(n6470), .B(n396), .C(n6466), .D(n364), .Z(n1158)
         );
  HS65_LH_AOI212X4 U2382 ( .A(\registers[18][21] ), .B(n6476), .C(
        \registers[24][21] ), .D(n6473), .E(n1144), .Z(n1143) );
  HS65_LH_OAI22X6 U2383 ( .A(n6470), .B(n395), .C(n6467), .D(n363), .Z(n1144)
         );
  HS65_LH_AOI212X4 U2384 ( .A(\registers[18][22] ), .B(n6476), .C(
        \registers[24][22] ), .D(n6473), .E(n1130), .Z(n1129) );
  HS65_LH_OAI22X6 U2385 ( .A(n6470), .B(n394), .C(n6467), .D(n362), .Z(n1130)
         );
  HS65_LH_AOI212X4 U2386 ( .A(\registers[18][23] ), .B(n6476), .C(
        \registers[24][23] ), .D(n6473), .E(n1116), .Z(n1115) );
  HS65_LH_OAI22X6 U2387 ( .A(n6470), .B(n393), .C(n6467), .D(n361), .Z(n1116)
         );
  HS65_LH_AOI212X4 U2388 ( .A(\registers[18][24] ), .B(n6476), .C(
        \registers[24][24] ), .D(n6473), .E(n1102), .Z(n1101) );
  HS65_LH_OAI22X6 U2389 ( .A(n6470), .B(n392), .C(n6467), .D(n360), .Z(n1102)
         );
  HS65_LH_AOI212X4 U2390 ( .A(\registers[18][25] ), .B(n6476), .C(
        \registers[24][25] ), .D(n6473), .E(n1088), .Z(n1087) );
  HS65_LH_OAI22X6 U2391 ( .A(n6470), .B(n391), .C(n6467), .D(n359), .Z(n1088)
         );
  HS65_LH_AOI212X4 U2392 ( .A(\registers[18][26] ), .B(n6476), .C(
        \registers[24][26] ), .D(n6473), .E(n1074), .Z(n1073) );
  HS65_LH_OAI22X6 U2393 ( .A(n6470), .B(n390), .C(n6467), .D(n358), .Z(n1074)
         );
  HS65_LH_AOI212X4 U2394 ( .A(\registers[18][27] ), .B(n6476), .C(
        \registers[24][27] ), .D(n6473), .E(n1060), .Z(n1059) );
  HS65_LH_OAI22X6 U2395 ( .A(n6470), .B(n389), .C(n6467), .D(n357), .Z(n1060)
         );
  HS65_LH_AOI212X4 U2396 ( .A(\registers[18][28] ), .B(n6476), .C(
        \registers[24][28] ), .D(n6473), .E(n1046), .Z(n1045) );
  HS65_LH_OAI22X6 U2397 ( .A(n6470), .B(n388), .C(n6467), .D(n356), .Z(n1046)
         );
  HS65_LH_AOI212X4 U2398 ( .A(\registers[18][29] ), .B(n6476), .C(
        \registers[24][29] ), .D(n6473), .E(n1032), .Z(n1031) );
  HS65_LH_OAI22X6 U2399 ( .A(n6470), .B(n387), .C(n6467), .D(n355), .Z(n1032)
         );
  HS65_LH_AOI212X4 U2400 ( .A(\registers[18][30] ), .B(n6476), .C(
        \registers[24][30] ), .D(n6473), .E(n1004), .Z(n1003) );
  HS65_LH_OAI22X6 U2401 ( .A(n6470), .B(n386), .C(n6467), .D(n354), .Z(n1004)
         );
  HS65_LH_AOI212X4 U2402 ( .A(\registers[18][31] ), .B(n6477), .C(
        \registers[24][31] ), .D(n6473), .E(n990), .Z(n989) );
  HS65_LH_OAI22X6 U2403 ( .A(n6471), .B(n385), .C(n6467), .D(n353), .Z(n990)
         );
  HS65_LH_NOR2X6 U2404 ( .A(n771), .B(\regfile_i[ADRREAD0][1] ), .Z(n2812) );
  HS65_LH_AOI212X4 U2405 ( .A(n6370), .B(n544), .C(n6367), .D(
        \registers[31][0] ), .E(n2821), .Z(n2816) );
  HS65_LH_OAI22X6 U2406 ( .A(n416), .B(n6364), .C(n352), .D(n6361), .Z(n2821)
         );
  HS65_LH_AOI212X4 U2407 ( .A(n6370), .B(n543), .C(n6367), .D(
        \registers[31][1] ), .E(n2656), .Z(n2653) );
  HS65_LH_OAI22X6 U2408 ( .A(n415), .B(n6364), .C(n351), .D(n6361), .Z(n2656)
         );
  HS65_LH_AOI212X4 U2409 ( .A(n6371), .B(n542), .C(n6368), .D(
        \registers[31][2] ), .E(n2502), .Z(n2499) );
  HS65_LH_OAI22X6 U2410 ( .A(n414), .B(n6365), .C(n350), .D(n6362), .Z(n2502)
         );
  HS65_LH_AOI212X4 U2411 ( .A(n6371), .B(n541), .C(n6368), .D(
        \registers[31][3] ), .E(n2460), .Z(n2457) );
  HS65_LH_OAI22X6 U2412 ( .A(n413), .B(n6366), .C(n349), .D(n6362), .Z(n2460)
         );
  HS65_LH_AOI212X4 U2413 ( .A(n6370), .B(n534), .C(n6367), .D(
        \registers[31][10] ), .E(n2796), .Z(n2793) );
  HS65_LH_OAI22X6 U2414 ( .A(n406), .B(n6364), .C(n342), .D(n6361), .Z(n2796)
         );
  HS65_LH_AOI212X4 U2415 ( .A(n6370), .B(n533), .C(n6367), .D(
        \registers[31][11] ), .E(n2782), .Z(n2779) );
  HS65_LH_OAI22X6 U2416 ( .A(n405), .B(n6364), .C(n341), .D(n6361), .Z(n2782)
         );
  HS65_LH_AOI212X4 U2417 ( .A(n6370), .B(n532), .C(n6367), .D(
        \registers[31][12] ), .E(n2768), .Z(n2765) );
  HS65_LH_OAI22X6 U2418 ( .A(n404), .B(n6364), .C(n340), .D(n6361), .Z(n2768)
         );
  HS65_LH_AOI212X4 U2419 ( .A(n6370), .B(n531), .C(n6367), .D(
        \registers[31][13] ), .E(n2754), .Z(n2751) );
  HS65_LH_OAI22X6 U2420 ( .A(n403), .B(n6364), .C(n339), .D(n6361), .Z(n2754)
         );
  HS65_LH_AOI212X4 U2421 ( .A(n6370), .B(n530), .C(n6367), .D(
        \registers[31][14] ), .E(n2740), .Z(n2737) );
  HS65_LH_OAI22X6 U2422 ( .A(n402), .B(n6364), .C(n338), .D(n6361), .Z(n2740)
         );
  HS65_LH_AOI212X4 U2423 ( .A(n6370), .B(n529), .C(n6367), .D(
        \registers[31][15] ), .E(n2726), .Z(n2723) );
  HS65_LH_OAI22X6 U2424 ( .A(n401), .B(n6364), .C(n337), .D(n6361), .Z(n2726)
         );
  HS65_LH_AOI212X4 U2425 ( .A(n6370), .B(n528), .C(n6367), .D(
        \registers[31][16] ), .E(n2712), .Z(n2709) );
  HS65_LH_OAI22X6 U2426 ( .A(n400), .B(n6364), .C(n336), .D(n6361), .Z(n2712)
         );
  HS65_LH_AOI212X4 U2427 ( .A(n6370), .B(n527), .C(n6367), .D(
        \registers[31][17] ), .E(n2698), .Z(n2695) );
  HS65_LH_OAI22X6 U2428 ( .A(n399), .B(n6364), .C(n335), .D(n6361), .Z(n2698)
         );
  HS65_LH_AOI212X4 U2429 ( .A(n6370), .B(n526), .C(n6367), .D(
        \registers[31][18] ), .E(n2684), .Z(n2681) );
  HS65_LH_OAI22X6 U2430 ( .A(n398), .B(n6364), .C(n334), .D(n6361), .Z(n2684)
         );
  HS65_LH_AOI212X4 U2431 ( .A(n6370), .B(n525), .C(n6367), .D(
        \registers[31][19] ), .E(n2670), .Z(n2667) );
  HS65_LH_OAI22X6 U2432 ( .A(n397), .B(n6364), .C(n333), .D(n6361), .Z(n2670)
         );
  HS65_LH_AOI212X4 U2433 ( .A(n6370), .B(n524), .C(n6367), .D(
        \registers[31][20] ), .E(n2642), .Z(n2639) );
  HS65_LH_OAI22X6 U2434 ( .A(n396), .B(n6365), .C(n332), .D(n6361), .Z(n2642)
         );
  HS65_LH_AOI212X4 U2435 ( .A(n6371), .B(n523), .C(n6368), .D(
        \registers[31][21] ), .E(n2628), .Z(n2625) );
  HS65_LH_OAI22X6 U2436 ( .A(n395), .B(n6365), .C(n331), .D(n6362), .Z(n2628)
         );
  HS65_LH_AOI212X4 U2437 ( .A(n6371), .B(n522), .C(n6368), .D(
        \registers[31][22] ), .E(n2614), .Z(n2611) );
  HS65_LH_OAI22X6 U2438 ( .A(n394), .B(n6365), .C(n330), .D(n6362), .Z(n2614)
         );
  HS65_LH_AOI212X4 U2439 ( .A(n6371), .B(n521), .C(n6368), .D(
        \registers[31][23] ), .E(n2600), .Z(n2597) );
  HS65_LH_OAI22X6 U2440 ( .A(n393), .B(n6365), .C(n329), .D(n6362), .Z(n2600)
         );
  HS65_LH_AOI212X4 U2441 ( .A(n6371), .B(n520), .C(n6368), .D(
        \registers[31][24] ), .E(n2586), .Z(n2583) );
  HS65_LH_OAI22X6 U2442 ( .A(n392), .B(n6365), .C(n328), .D(n6362), .Z(n2586)
         );
  HS65_LH_AOI212X4 U2443 ( .A(n6371), .B(n519), .C(n6368), .D(
        \registers[31][25] ), .E(n2572), .Z(n2569) );
  HS65_LH_OAI22X6 U2444 ( .A(n391), .B(n6365), .C(n327), .D(n6362), .Z(n2572)
         );
  HS65_LH_AOI212X4 U2445 ( .A(n6371), .B(n518), .C(n6368), .D(
        \registers[31][26] ), .E(n2558), .Z(n2555) );
  HS65_LH_OAI22X6 U2446 ( .A(n390), .B(n6365), .C(n326), .D(n6362), .Z(n2558)
         );
  HS65_LH_AOI212X4 U2447 ( .A(n6371), .B(n517), .C(n6368), .D(
        \registers[31][27] ), .E(n2544), .Z(n2541) );
  HS65_LH_OAI22X6 U2448 ( .A(n389), .B(n6365), .C(n325), .D(n6362), .Z(n2544)
         );
  HS65_LH_AOI212X4 U2449 ( .A(n6371), .B(n516), .C(n6368), .D(
        \registers[31][28] ), .E(n2530), .Z(n2527) );
  HS65_LH_OAI22X6 U2450 ( .A(n388), .B(n6365), .C(n324), .D(n6362), .Z(n2530)
         );
  HS65_LH_AOI212X4 U2451 ( .A(n6371), .B(n515), .C(n6368), .D(
        \registers[31][29] ), .E(n2516), .Z(n2513) );
  HS65_LH_OAI22X6 U2452 ( .A(n387), .B(n6365), .C(n323), .D(n6362), .Z(n2516)
         );
  HS65_LH_AOI212X4 U2453 ( .A(n6371), .B(n514), .C(n6368), .D(
        \registers[31][30] ), .E(n2488), .Z(n2485) );
  HS65_LH_OAI22X6 U2454 ( .A(n386), .B(n6365), .C(n322), .D(n6362), .Z(n2488)
         );
  HS65_LH_AOI212X4 U2455 ( .A(n6371), .B(n513), .C(n6368), .D(
        \registers[31][31] ), .E(n2474), .Z(n2471) );
  HS65_LH_OAI22X6 U2456 ( .A(n385), .B(n6366), .C(n321), .D(n6362), .Z(n2474)
         );
  HS65_LH_AOI212X4 U2457 ( .A(n6372), .B(n540), .C(n6369), .D(
        \registers[31][4] ), .E(n2446), .Z(n2443) );
  HS65_LH_OAI22X6 U2458 ( .A(n412), .B(n6366), .C(n348), .D(n6363), .Z(n2446)
         );
  HS65_LH_AOI212X4 U2459 ( .A(n6372), .B(n539), .C(n6369), .D(
        \registers[31][5] ), .E(n2432), .Z(n2429) );
  HS65_LH_OAI22X6 U2460 ( .A(n411), .B(n6366), .C(n347), .D(n6363), .Z(n2432)
         );
  HS65_LH_AOI212X4 U2461 ( .A(n6372), .B(n538), .C(n6369), .D(
        \registers[31][6] ), .E(n1426), .Z(n1423) );
  HS65_LH_OAI22X6 U2462 ( .A(n410), .B(n6366), .C(n346), .D(n6363), .Z(n1426)
         );
  HS65_LH_AOI212X4 U2463 ( .A(n6372), .B(n537), .C(n6369), .D(
        \registers[31][7] ), .E(n1412), .Z(n1409) );
  HS65_LH_OAI22X6 U2464 ( .A(n409), .B(n6366), .C(n345), .D(n6363), .Z(n1412)
         );
  HS65_LH_AOI212X4 U2465 ( .A(n6372), .B(n536), .C(n6369), .D(
        \registers[31][8] ), .E(n1398), .Z(n1395) );
  HS65_LH_OAI22X6 U2466 ( .A(n408), .B(n6366), .C(n344), .D(n6363), .Z(n1398)
         );
  HS65_LH_AOI212X4 U2467 ( .A(n6372), .B(n535), .C(n6369), .D(
        \registers[31][9] ), .E(n1374), .Z(n1365) );
  HS65_LH_OAI22X6 U2468 ( .A(n407), .B(n6366), .C(n343), .D(n6363), .Z(n1374)
         );
  HS65_LH_AOI212X4 U2469 ( .A(n6427), .B(n672), .C(n6424), .D(
        \registers[11][0] ), .E(n2804), .Z(n2803) );
  HS65_LH_OAI22X6 U2470 ( .A(n224), .B(n6421), .C(n160), .D(n6418), .Z(n2804)
         );
  HS65_LH_AOI212X4 U2471 ( .A(n6427), .B(n671), .C(n6424), .D(
        \registers[11][1] ), .E(n2650), .Z(n2649) );
  HS65_LH_OAI22X6 U2472 ( .A(n223), .B(n6421), .C(n159), .D(n6418), .Z(n2650)
         );
  HS65_LH_AOI212X4 U2473 ( .A(n6428), .B(n670), .C(n6425), .D(
        \registers[11][2] ), .E(n2496), .Z(n2495) );
  HS65_LH_OAI22X6 U2474 ( .A(n222), .B(n6422), .C(n158), .D(n6419), .Z(n2496)
         );
  HS65_LH_AOI212X4 U2475 ( .A(n6428), .B(n669), .C(n6425), .D(
        \registers[11][3] ), .E(n2454), .Z(n2453) );
  HS65_LH_OAI22X6 U2476 ( .A(n221), .B(n6423), .C(n157), .D(n6419), .Z(n2454)
         );
  HS65_LH_AOI212X4 U2477 ( .A(n6429), .B(n668), .C(n6426), .D(
        \registers[11][4] ), .E(n2440), .Z(n2439) );
  HS65_LH_OAI22X6 U2478 ( .A(n220), .B(n6423), .C(n156), .D(n6420), .Z(n2440)
         );
  HS65_LH_AOI212X4 U2479 ( .A(n6429), .B(n667), .C(n6426), .D(
        \registers[11][5] ), .E(n2426), .Z(n1433) );
  HS65_LH_OAI22X6 U2480 ( .A(n219), .B(n6423), .C(n155), .D(n6420), .Z(n2426)
         );
  HS65_LH_AOI212X4 U2481 ( .A(n6429), .B(n666), .C(n6426), .D(
        \registers[11][6] ), .E(n1420), .Z(n1419) );
  HS65_LH_OAI22X6 U2482 ( .A(n218), .B(n6423), .C(n154), .D(n6420), .Z(n1420)
         );
  HS65_LH_AOI212X4 U2483 ( .A(n6429), .B(n665), .C(n6426), .D(
        \registers[11][7] ), .E(n1406), .Z(n1405) );
  HS65_LH_OAI22X6 U2484 ( .A(n217), .B(n6423), .C(n153), .D(n6420), .Z(n1406)
         );
  HS65_LH_AOI212X4 U2485 ( .A(n6429), .B(n664), .C(n6426), .D(
        \registers[11][8] ), .E(n1392), .Z(n1391) );
  HS65_LH_OAI22X6 U2486 ( .A(n216), .B(n6423), .C(n152), .D(n6420), .Z(n1392)
         );
  HS65_LH_AOI212X4 U2487 ( .A(n6429), .B(n663), .C(n6426), .D(
        \registers[11][9] ), .E(n1349), .Z(n1346) );
  HS65_LH_OAI22X6 U2488 ( .A(n215), .B(n6423), .C(n151), .D(n6420), .Z(n1349)
         );
  HS65_LH_AOI212X4 U2489 ( .A(n6427), .B(n662), .C(n6424), .D(
        \registers[11][10] ), .E(n2790), .Z(n2789) );
  HS65_LH_OAI22X6 U2490 ( .A(n214), .B(n6421), .C(n150), .D(n6418), .Z(n2790)
         );
  HS65_LH_AOI212X4 U2491 ( .A(n6427), .B(n661), .C(n6424), .D(
        \registers[11][11] ), .E(n2776), .Z(n2775) );
  HS65_LH_OAI22X6 U2492 ( .A(n213), .B(n6421), .C(n149), .D(n6418), .Z(n2776)
         );
  HS65_LH_AOI212X4 U2493 ( .A(n6427), .B(n660), .C(n6424), .D(
        \registers[11][12] ), .E(n2762), .Z(n2761) );
  HS65_LH_OAI22X6 U2494 ( .A(n212), .B(n6421), .C(n148), .D(n6418), .Z(n2762)
         );
  HS65_LH_AOI212X4 U2495 ( .A(n6427), .B(n659), .C(n6424), .D(
        \registers[11][13] ), .E(n2748), .Z(n2747) );
  HS65_LH_OAI22X6 U2496 ( .A(n211), .B(n6421), .C(n147), .D(n6418), .Z(n2748)
         );
  HS65_LH_AOI212X4 U2497 ( .A(n6427), .B(n658), .C(n6424), .D(
        \registers[11][14] ), .E(n2734), .Z(n2733) );
  HS65_LH_OAI22X6 U2498 ( .A(n210), .B(n6421), .C(n146), .D(n6418), .Z(n2734)
         );
  HS65_LH_AOI212X4 U2499 ( .A(n6427), .B(n657), .C(n6424), .D(
        \registers[11][15] ), .E(n2720), .Z(n2719) );
  HS65_LH_OAI22X6 U2500 ( .A(n209), .B(n6421), .C(n145), .D(n6418), .Z(n2720)
         );
  HS65_LH_AOI212X4 U2501 ( .A(n6427), .B(n656), .C(n6424), .D(
        \registers[11][16] ), .E(n2706), .Z(n2705) );
  HS65_LH_OAI22X6 U2502 ( .A(n208), .B(n6421), .C(n144), .D(n6418), .Z(n2706)
         );
  HS65_LH_AOI212X4 U2503 ( .A(n6427), .B(n655), .C(n6424), .D(
        \registers[11][17] ), .E(n2692), .Z(n2691) );
  HS65_LH_OAI22X6 U2504 ( .A(n207), .B(n6421), .C(n143), .D(n6418), .Z(n2692)
         );
  HS65_LH_AOI212X4 U2505 ( .A(n6427), .B(n654), .C(n6424), .D(
        \registers[11][18] ), .E(n2678), .Z(n2677) );
  HS65_LH_OAI22X6 U2506 ( .A(n206), .B(n6421), .C(n142), .D(n6418), .Z(n2678)
         );
  HS65_LH_AOI212X4 U2507 ( .A(n6427), .B(n653), .C(n6424), .D(
        \registers[11][19] ), .E(n2664), .Z(n2663) );
  HS65_LH_OAI22X6 U2508 ( .A(n205), .B(n6421), .C(n141), .D(n6418), .Z(n2664)
         );
  HS65_LH_AOI212X4 U2509 ( .A(n6427), .B(n652), .C(n6424), .D(
        \registers[11][20] ), .E(n2636), .Z(n2635) );
  HS65_LH_OAI22X6 U2510 ( .A(n204), .B(n6422), .C(n140), .D(n6418), .Z(n2636)
         );
  HS65_LH_AOI212X4 U2511 ( .A(n6428), .B(n651), .C(n6425), .D(
        \registers[11][21] ), .E(n2622), .Z(n2621) );
  HS65_LH_OAI22X6 U2512 ( .A(n203), .B(n6422), .C(n139), .D(n6419), .Z(n2622)
         );
  HS65_LH_AOI212X4 U2513 ( .A(n6428), .B(n650), .C(n6425), .D(
        \registers[11][22] ), .E(n2608), .Z(n2607) );
  HS65_LH_OAI22X6 U2514 ( .A(n202), .B(n6422), .C(n138), .D(n6419), .Z(n2608)
         );
  HS65_LH_AOI212X4 U2515 ( .A(n6428), .B(n649), .C(n6425), .D(
        \registers[11][23] ), .E(n2594), .Z(n2593) );
  HS65_LH_OAI22X6 U2516 ( .A(n201), .B(n6422), .C(n137), .D(n6419), .Z(n2594)
         );
  HS65_LH_AOI212X4 U2517 ( .A(n6428), .B(n648), .C(n6425), .D(
        \registers[11][24] ), .E(n2580), .Z(n2579) );
  HS65_LH_OAI22X6 U2518 ( .A(n200), .B(n6422), .C(n136), .D(n6419), .Z(n2580)
         );
  HS65_LH_AOI212X4 U2519 ( .A(n6428), .B(n647), .C(n6425), .D(
        \registers[11][25] ), .E(n2566), .Z(n2565) );
  HS65_LH_OAI22X6 U2520 ( .A(n199), .B(n6422), .C(n135), .D(n6419), .Z(n2566)
         );
  HS65_LH_AOI212X4 U2521 ( .A(n6428), .B(n646), .C(n6425), .D(
        \registers[11][26] ), .E(n2552), .Z(n2551) );
  HS65_LH_OAI22X6 U2522 ( .A(n198), .B(n6422), .C(n134), .D(n6419), .Z(n2552)
         );
  HS65_LH_AOI212X4 U2523 ( .A(n6428), .B(n645), .C(n6425), .D(
        \registers[11][27] ), .E(n2538), .Z(n2537) );
  HS65_LH_OAI22X6 U2524 ( .A(n197), .B(n6422), .C(n133), .D(n6419), .Z(n2538)
         );
  HS65_LH_AOI212X4 U2525 ( .A(n6428), .B(n644), .C(n6425), .D(
        \registers[11][28] ), .E(n2524), .Z(n2523) );
  HS65_LH_OAI22X6 U2526 ( .A(n196), .B(n6422), .C(n132), .D(n6419), .Z(n2524)
         );
  HS65_LH_AOI212X4 U2527 ( .A(n6428), .B(n643), .C(n6425), .D(
        \registers[11][29] ), .E(n2510), .Z(n2509) );
  HS65_LH_OAI22X6 U2528 ( .A(n195), .B(n6422), .C(n131), .D(n6419), .Z(n2510)
         );
  HS65_LH_AOI212X4 U2529 ( .A(n6428), .B(n642), .C(n6425), .D(
        \registers[11][30] ), .E(n2482), .Z(n2481) );
  HS65_LH_OAI22X6 U2530 ( .A(n194), .B(n6422), .C(n130), .D(n6419), .Z(n2482)
         );
  HS65_LH_AOI212X4 U2531 ( .A(n6428), .B(n641), .C(n6425), .D(
        \registers[11][31] ), .E(n2468), .Z(n2467) );
  HS65_LH_OAI22X6 U2532 ( .A(n193), .B(n6423), .C(n129), .D(n6419), .Z(n2468)
         );
  HS65_LH_AOI212X4 U2533 ( .A(n6382), .B(\registers[17][0] ), .C(n6379), .D(
        \registers[19][0] ), .E(n2818), .Z(n2817) );
  HS65_LH_OAI22X6 U2534 ( .A(n288), .B(n6376), .C(n320), .D(n6373), .Z(n2818)
         );
  HS65_LH_AOI212X4 U2535 ( .A(n6382), .B(\registers[17][1] ), .C(n6379), .D(
        \registers[19][1] ), .E(n2655), .Z(n2654) );
  HS65_LH_OAI22X6 U2536 ( .A(n287), .B(n6376), .C(n319), .D(n6373), .Z(n2655)
         );
  HS65_LH_AOI212X4 U2537 ( .A(n6383), .B(\registers[17][2] ), .C(n6380), .D(
        \registers[19][2] ), .E(n2501), .Z(n2500) );
  HS65_LH_OAI22X6 U2538 ( .A(n286), .B(n6377), .C(n318), .D(n6374), .Z(n2501)
         );
  HS65_LH_AOI212X4 U2539 ( .A(n6383), .B(\registers[17][3] ), .C(n6380), .D(
        \registers[19][3] ), .E(n2459), .Z(n2458) );
  HS65_LH_OAI22X6 U2540 ( .A(n285), .B(n6378), .C(n317), .D(n6374), .Z(n2459)
         );
  HS65_LH_AOI212X4 U2541 ( .A(n6382), .B(\registers[17][10] ), .C(n6379), .D(
        \registers[19][10] ), .E(n2795), .Z(n2794) );
  HS65_LH_OAI22X6 U2542 ( .A(n278), .B(n6376), .C(n310), .D(n6373), .Z(n2795)
         );
  HS65_LH_AOI212X4 U2543 ( .A(n6382), .B(\registers[17][11] ), .C(n6379), .D(
        \registers[19][11] ), .E(n2781), .Z(n2780) );
  HS65_LH_OAI22X6 U2544 ( .A(n277), .B(n6376), .C(n309), .D(n6373), .Z(n2781)
         );
  HS65_LH_AOI212X4 U2545 ( .A(n6382), .B(\registers[17][12] ), .C(n6379), .D(
        \registers[19][12] ), .E(n2767), .Z(n2766) );
  HS65_LH_OAI22X6 U2546 ( .A(n276), .B(n6376), .C(n308), .D(n6373), .Z(n2767)
         );
  HS65_LH_AOI212X4 U2547 ( .A(n6382), .B(\registers[17][13] ), .C(n6379), .D(
        \registers[19][13] ), .E(n2753), .Z(n2752) );
  HS65_LH_OAI22X6 U2548 ( .A(n275), .B(n6376), .C(n307), .D(n6373), .Z(n2753)
         );
  HS65_LH_AOI212X4 U2549 ( .A(n6382), .B(\registers[17][14] ), .C(n6379), .D(
        \registers[19][14] ), .E(n2739), .Z(n2738) );
  HS65_LH_OAI22X6 U2550 ( .A(n274), .B(n6376), .C(n306), .D(n6373), .Z(n2739)
         );
  HS65_LH_AOI212X4 U2551 ( .A(n6382), .B(\registers[17][15] ), .C(n6379), .D(
        \registers[19][15] ), .E(n2725), .Z(n2724) );
  HS65_LH_OAI22X6 U2552 ( .A(n273), .B(n6376), .C(n305), .D(n6373), .Z(n2725)
         );
  HS65_LH_AOI212X4 U2553 ( .A(n6382), .B(\registers[17][16] ), .C(n6379), .D(
        \registers[19][16] ), .E(n2711), .Z(n2710) );
  HS65_LH_OAI22X6 U2554 ( .A(n272), .B(n6376), .C(n304), .D(n6373), .Z(n2711)
         );
  HS65_LH_AOI212X4 U2555 ( .A(n6382), .B(\registers[17][17] ), .C(n6379), .D(
        \registers[19][17] ), .E(n2697), .Z(n2696) );
  HS65_LH_OAI22X6 U2556 ( .A(n271), .B(n6376), .C(n303), .D(n6373), .Z(n2697)
         );
  HS65_LH_AOI212X4 U2557 ( .A(n6382), .B(\registers[17][18] ), .C(n6379), .D(
        \registers[19][18] ), .E(n2683), .Z(n2682) );
  HS65_LH_OAI22X6 U2558 ( .A(n270), .B(n6376), .C(n302), .D(n6373), .Z(n2683)
         );
  HS65_LH_AOI212X4 U2559 ( .A(n6382), .B(\registers[17][19] ), .C(n6379), .D(
        \registers[19][19] ), .E(n2669), .Z(n2668) );
  HS65_LH_OAI22X6 U2560 ( .A(n269), .B(n6376), .C(n301), .D(n6373), .Z(n2669)
         );
  HS65_LH_AOI212X4 U2561 ( .A(n6382), .B(\registers[17][20] ), .C(n6379), .D(
        \registers[19][20] ), .E(n2641), .Z(n2640) );
  HS65_LH_OAI22X6 U2562 ( .A(n268), .B(n6377), .C(n300), .D(n6373), .Z(n2641)
         );
  HS65_LH_AOI212X4 U2563 ( .A(n6383), .B(\registers[17][21] ), .C(n6380), .D(
        \registers[19][21] ), .E(n2627), .Z(n2626) );
  HS65_LH_OAI22X6 U2564 ( .A(n267), .B(n6377), .C(n299), .D(n6374), .Z(n2627)
         );
  HS65_LH_AOI212X4 U2565 ( .A(n6383), .B(\registers[17][22] ), .C(n6380), .D(
        \registers[19][22] ), .E(n2613), .Z(n2612) );
  HS65_LH_OAI22X6 U2566 ( .A(n266), .B(n6377), .C(n298), .D(n6374), .Z(n2613)
         );
  HS65_LH_AOI212X4 U2567 ( .A(n6383), .B(\registers[17][23] ), .C(n6380), .D(
        \registers[19][23] ), .E(n2599), .Z(n2598) );
  HS65_LH_OAI22X6 U2568 ( .A(n265), .B(n6377), .C(n297), .D(n6374), .Z(n2599)
         );
  HS65_LH_AOI212X4 U2569 ( .A(n6383), .B(\registers[17][24] ), .C(n6380), .D(
        \registers[19][24] ), .E(n2585), .Z(n2584) );
  HS65_LH_OAI22X6 U2570 ( .A(n264), .B(n6377), .C(n296), .D(n6374), .Z(n2585)
         );
  HS65_LH_AOI212X4 U2571 ( .A(n6383), .B(\registers[17][25] ), .C(n6380), .D(
        \registers[19][25] ), .E(n2571), .Z(n2570) );
  HS65_LH_OAI22X6 U2572 ( .A(n263), .B(n6377), .C(n295), .D(n6374), .Z(n2571)
         );
  HS65_LH_AOI212X4 U2573 ( .A(n6383), .B(\registers[17][26] ), .C(n6380), .D(
        \registers[19][26] ), .E(n2557), .Z(n2556) );
  HS65_LH_OAI22X6 U2574 ( .A(n262), .B(n6377), .C(n294), .D(n6374), .Z(n2557)
         );
  HS65_LH_AOI212X4 U2575 ( .A(n6383), .B(\registers[17][27] ), .C(n6380), .D(
        \registers[19][27] ), .E(n2543), .Z(n2542) );
  HS65_LH_OAI22X6 U2576 ( .A(n261), .B(n6377), .C(n293), .D(n6374), .Z(n2543)
         );
  HS65_LH_AOI212X4 U2577 ( .A(n6383), .B(\registers[17][28] ), .C(n6380), .D(
        \registers[19][28] ), .E(n2529), .Z(n2528) );
  HS65_LH_OAI22X6 U2578 ( .A(n260), .B(n6377), .C(n292), .D(n6374), .Z(n2529)
         );
  HS65_LH_AOI212X4 U2579 ( .A(n6383), .B(\registers[17][29] ), .C(n6380), .D(
        \registers[19][29] ), .E(n2515), .Z(n2514) );
  HS65_LH_OAI22X6 U2580 ( .A(n259), .B(n6377), .C(n291), .D(n6374), .Z(n2515)
         );
  HS65_LH_AOI212X4 U2581 ( .A(n6383), .B(\registers[17][30] ), .C(n6380), .D(
        \registers[19][30] ), .E(n2487), .Z(n2486) );
  HS65_LH_OAI22X6 U2582 ( .A(n258), .B(n6377), .C(n290), .D(n6374), .Z(n2487)
         );
  HS65_LH_AOI212X4 U2583 ( .A(n6383), .B(\registers[17][31] ), .C(n6380), .D(
        \registers[19][31] ), .E(n2473), .Z(n2472) );
  HS65_LH_OAI22X6 U2584 ( .A(n257), .B(n6378), .C(n289), .D(n6374), .Z(n2473)
         );
  HS65_LH_AOI212X4 U2585 ( .A(n6384), .B(\registers[17][4] ), .C(n6381), .D(
        \registers[19][4] ), .E(n2445), .Z(n2444) );
  HS65_LH_OAI22X6 U2586 ( .A(n284), .B(n6378), .C(n316), .D(n6375), .Z(n2445)
         );
  HS65_LH_AOI212X4 U2587 ( .A(n6384), .B(\registers[17][5] ), .C(n6381), .D(
        \registers[19][5] ), .E(n2431), .Z(n2430) );
  HS65_LH_OAI22X6 U2588 ( .A(n283), .B(n6378), .C(n315), .D(n6375), .Z(n2431)
         );
  HS65_LH_AOI212X4 U2589 ( .A(n6384), .B(\registers[17][6] ), .C(n6381), .D(
        \registers[19][6] ), .E(n1425), .Z(n1424) );
  HS65_LH_OAI22X6 U2590 ( .A(n282), .B(n6378), .C(n314), .D(n6375), .Z(n1425)
         );
  HS65_LH_AOI212X4 U2591 ( .A(n6384), .B(\registers[17][7] ), .C(n6381), .D(
        \registers[19][7] ), .E(n1411), .Z(n1410) );
  HS65_LH_OAI22X6 U2592 ( .A(n281), .B(n6378), .C(n313), .D(n6375), .Z(n1411)
         );
  HS65_LH_AOI212X4 U2593 ( .A(n6384), .B(\registers[17][8] ), .C(n6381), .D(
        \registers[19][8] ), .E(n1397), .Z(n1396) );
  HS65_LH_OAI22X6 U2594 ( .A(n280), .B(n6378), .C(n312), .D(n6375), .Z(n1397)
         );
  HS65_LH_AOI212X4 U2595 ( .A(n6384), .B(\registers[17][9] ), .C(n6381), .D(
        \registers[19][9] ), .E(n1369), .Z(n1366) );
  HS65_LH_OAI22X6 U2596 ( .A(n279), .B(n6378), .C(n311), .D(n6375), .Z(n1369)
         );
  HS65_LH_NOR3X4 U2597 ( .A(\regfile_i[ADRREAD0][3] ), .B(
        \regfile_i[ADRREAD0][4] ), .C(\regfile_i[ADRREAD0][0] ), .Z(n2810) );
  HS65_LH_NAND4ABX3 U2598 ( .A(n1308), .B(n1309), .C(n1310), .D(n1311), .Z(
        n1301) );
  HS65_LH_MX41X7 U2599 ( .D0(\registers[22][10] ), .S0(n6439), .D1(
        \registers[21][10] ), .S1(n6436), .D2(\registers[19][10] ), .S2(n6433), 
        .D3(n6430), .S3(n598), .Z(n1308) );
  HS65_LH_MX41X7 U2600 ( .D0(n6451), .S0(n758), .D1(\registers[30][10] ), .S1(
        n6448), .D2(n6445), .S2(n662), .D3(\registers[20][10] ), .S3(n6442), 
        .Z(n1309) );
  HS65_LH_AOI212X4 U2601 ( .A(\registers[18][10] ), .B(n6475), .C(
        \registers[24][10] ), .D(n6472), .E(n1312), .Z(n1311) );
  HS65_LH_IVX9 U2602 ( .A(\regfile_i[ADRREAD1][4] ), .Z(n774) );
  HS65_LH_IVX9 U2603 ( .A(\regfile_i[ADRREAD0][3] ), .Z(n770) );
  HS65_LH_IVX9 U2604 ( .A(\regfile_i[ADRWRITE][0] ), .Z(n814) );
  HS65_LH_IVX9 U2605 ( .A(\regfile_i[ADRREAD1][3] ), .Z(n775) );
  HS65_LH_IVX9 U2606 ( .A(\regfile_i[ADRREAD0][4] ), .Z(n769) );
  HS65_LH_IVX9 U2607 ( .A(\regfile_i[ADRWRITE][1] ), .Z(n813) );
  HS65_LH_MX41X7 U2608 ( .D0(\registers[5][0] ), .S0(n6487), .D1(
        \registers[11][0] ), .S1(n6484), .D2(\registers[7][0] ), .S2(n6481), 
        .D3(\registers[3][0] ), .S3(n6478), .Z(n1317) );
  HS65_LH_MX41X7 U2609 ( .D0(\registers[5][1] ), .S0(n6487), .D1(
        \registers[11][1] ), .S1(n6484), .D2(\registers[7][1] ), .S2(n6481), 
        .D3(\registers[3][1] ), .S3(n6478), .Z(n1163) );
  HS65_LH_MX41X7 U2610 ( .D0(\registers[5][2] ), .S0(n6488), .D1(
        \registers[11][2] ), .S1(n6485), .D2(\registers[7][2] ), .S2(n6482), 
        .D3(\registers[3][2] ), .S3(n6479), .Z(n1009) );
  HS65_LH_MX41X7 U2611 ( .D0(\registers[5][3] ), .S0(n6489), .D1(
        \registers[11][3] ), .S1(n6486), .D2(\registers[7][3] ), .S2(n6483), 
        .D3(\registers[3][3] ), .S3(n6480), .Z(n967) );
  HS65_LH_MX41X7 U2612 ( .D0(\registers[5][4] ), .S0(n6489), .D1(
        \registers[11][4] ), .S1(n6486), .D2(\registers[7][4] ), .S2(n6483), 
        .D3(\registers[3][4] ), .S3(n6480), .Z(n953) );
  HS65_LH_MX41X7 U2613 ( .D0(\registers[5][5] ), .S0(n6489), .D1(
        \registers[11][5] ), .S1(n6486), .D2(\registers[7][5] ), .S2(n6483), 
        .D3(\registers[3][5] ), .S3(n6480), .Z(n939) );
  HS65_LH_MX41X7 U2614 ( .D0(\registers[5][6] ), .S0(n6489), .D1(
        \registers[11][6] ), .S1(n6486), .D2(\registers[7][6] ), .S2(n6483), 
        .D3(\registers[3][6] ), .S3(n6480), .Z(n925) );
  HS65_LH_MX41X7 U2615 ( .D0(\registers[5][7] ), .S0(n6489), .D1(
        \registers[11][7] ), .S1(n6486), .D2(\registers[7][7] ), .S2(n6483), 
        .D3(\registers[3][7] ), .S3(n6480), .Z(n911) );
  HS65_LH_MX41X7 U2616 ( .D0(\registers[5][8] ), .S0(n6489), .D1(
        \registers[11][8] ), .S1(n6486), .D2(\registers[7][8] ), .S2(n6483), 
        .D3(\registers[3][8] ), .S3(n6480), .Z(n897) );
  HS65_LH_MX41X7 U2617 ( .D0(\registers[5][9] ), .S0(n6489), .D1(
        \registers[11][9] ), .S1(n6486), .D2(\registers[7][9] ), .S2(n6483), 
        .D3(\registers[3][9] ), .S3(n6480), .Z(n852) );
  HS65_LH_MX41X7 U2618 ( .D0(\registers[5][10] ), .S0(n6487), .D1(
        \registers[11][10] ), .S1(n6484), .D2(\registers[7][10] ), .S2(n6481), 
        .D3(\registers[3][10] ), .S3(n6478), .Z(n1303) );
  HS65_LH_MX41X7 U2619 ( .D0(\registers[5][11] ), .S0(n6487), .D1(
        \registers[11][11] ), .S1(n6484), .D2(\registers[7][11] ), .S2(n6481), 
        .D3(\registers[3][11] ), .S3(n6478), .Z(n1289) );
  HS65_LH_MX41X7 U2620 ( .D0(\registers[5][12] ), .S0(n6487), .D1(
        \registers[11][12] ), .S1(n6484), .D2(\registers[7][12] ), .S2(n6481), 
        .D3(\registers[3][12] ), .S3(n6478), .Z(n1275) );
  HS65_LH_MX41X7 U2621 ( .D0(\registers[5][13] ), .S0(n6487), .D1(
        \registers[11][13] ), .S1(n6484), .D2(\registers[7][13] ), .S2(n6481), 
        .D3(\registers[3][13] ), .S3(n6478), .Z(n1261) );
  HS65_LH_MX41X7 U2622 ( .D0(\registers[5][14] ), .S0(n6487), .D1(
        \registers[11][14] ), .S1(n6484), .D2(\registers[7][14] ), .S2(n6481), 
        .D3(\registers[3][14] ), .S3(n6478), .Z(n1247) );
  HS65_LH_MX41X7 U2623 ( .D0(\registers[5][15] ), .S0(n6487), .D1(
        \registers[11][15] ), .S1(n6484), .D2(\registers[7][15] ), .S2(n6481), 
        .D3(\registers[3][15] ), .S3(n6478), .Z(n1233) );
  HS65_LH_MX41X7 U2624 ( .D0(\registers[5][16] ), .S0(n6487), .D1(
        \registers[11][16] ), .S1(n6484), .D2(\registers[7][16] ), .S2(n6481), 
        .D3(\registers[3][16] ), .S3(n6478), .Z(n1219) );
  HS65_LH_MX41X7 U2625 ( .D0(\registers[5][17] ), .S0(n6487), .D1(
        \registers[11][17] ), .S1(n6484), .D2(\registers[7][17] ), .S2(n6481), 
        .D3(\registers[3][17] ), .S3(n6478), .Z(n1205) );
  HS65_LH_MX41X7 U2626 ( .D0(\registers[5][18] ), .S0(n6487), .D1(
        \registers[11][18] ), .S1(n6484), .D2(\registers[7][18] ), .S2(n6481), 
        .D3(\registers[3][18] ), .S3(n6478), .Z(n1191) );
  HS65_LH_MX41X7 U2627 ( .D0(\registers[5][19] ), .S0(n6487), .D1(
        \registers[11][19] ), .S1(n6484), .D2(\registers[7][19] ), .S2(n6481), 
        .D3(\registers[3][19] ), .S3(n6478), .Z(n1177) );
  HS65_LH_MX41X7 U2628 ( .D0(\registers[5][20] ), .S0(n6488), .D1(
        \registers[11][20] ), .S1(n6485), .D2(\registers[7][20] ), .S2(n6482), 
        .D3(\registers[3][20] ), .S3(n6479), .Z(n1149) );
  HS65_LH_MX41X7 U2629 ( .D0(\registers[5][21] ), .S0(n6488), .D1(
        \registers[11][21] ), .S1(n6485), .D2(\registers[7][21] ), .S2(n6482), 
        .D3(\registers[3][21] ), .S3(n6479), .Z(n1135) );
  HS65_LH_MX41X7 U2630 ( .D0(\registers[5][22] ), .S0(n6488), .D1(
        \registers[11][22] ), .S1(n6485), .D2(\registers[7][22] ), .S2(n6482), 
        .D3(\registers[3][22] ), .S3(n6479), .Z(n1121) );
  HS65_LH_MX41X7 U2631 ( .D0(\registers[5][23] ), .S0(n6488), .D1(
        \registers[11][23] ), .S1(n6485), .D2(\registers[7][23] ), .S2(n6482), 
        .D3(\registers[3][23] ), .S3(n6479), .Z(n1107) );
  HS65_LH_MX41X7 U2632 ( .D0(\registers[5][24] ), .S0(n6488), .D1(
        \registers[11][24] ), .S1(n6485), .D2(\registers[7][24] ), .S2(n6482), 
        .D3(\registers[3][24] ), .S3(n6479), .Z(n1093) );
  HS65_LH_MX41X7 U2633 ( .D0(\registers[5][25] ), .S0(n6488), .D1(
        \registers[11][25] ), .S1(n6485), .D2(\registers[7][25] ), .S2(n6482), 
        .D3(\registers[3][25] ), .S3(n6479), .Z(n1079) );
  HS65_LH_MX41X7 U2634 ( .D0(\registers[5][26] ), .S0(n6488), .D1(
        \registers[11][26] ), .S1(n6485), .D2(\registers[7][26] ), .S2(n6482), 
        .D3(\registers[3][26] ), .S3(n6479), .Z(n1065) );
  HS65_LH_MX41X7 U2635 ( .D0(\registers[5][27] ), .S0(n6488), .D1(
        \registers[11][27] ), .S1(n6485), .D2(\registers[7][27] ), .S2(n6482), 
        .D3(\registers[3][27] ), .S3(n6479), .Z(n1051) );
  HS65_LH_MX41X7 U2636 ( .D0(\registers[5][28] ), .S0(n6488), .D1(
        \registers[11][28] ), .S1(n6485), .D2(\registers[7][28] ), .S2(n6482), 
        .D3(\registers[3][28] ), .S3(n6479), .Z(n1037) );
  HS65_LH_MX41X7 U2637 ( .D0(\registers[5][29] ), .S0(n6488), .D1(
        \registers[11][29] ), .S1(n6485), .D2(\registers[7][29] ), .S2(n6482), 
        .D3(\registers[3][29] ), .S3(n6479), .Z(n1023) );
  HS65_LH_MX41X7 U2638 ( .D0(\registers[5][30] ), .S0(n6488), .D1(
        \registers[11][30] ), .S1(n6485), .D2(\registers[7][30] ), .S2(n6482), 
        .D3(\registers[3][30] ), .S3(n6479), .Z(n995) );
  HS65_LH_MX41X7 U2639 ( .D0(\registers[5][31] ), .S0(n6489), .D1(
        \registers[11][31] ), .S1(n6486), .D2(\registers[7][31] ), .S2(n6483), 
        .D3(\registers[3][31] ), .S3(n6480), .Z(n981) );
  HS65_LH_MX41X7 U2640 ( .D0(n6451), .S0(n768), .D1(\registers[30][0] ), .S1(
        n6448), .D2(n6445), .S2(n672), .D3(\registers[20][0] ), .S3(n6442), 
        .Z(n1333) );
  HS65_LH_MX41X7 U2641 ( .D0(n6451), .S0(n767), .D1(\registers[30][1] ), .S1(
        n6448), .D2(n6445), .S2(n671), .D3(\registers[20][1] ), .S3(n6442), 
        .Z(n1169) );
  HS65_LH_MX41X7 U2642 ( .D0(n6452), .S0(n766), .D1(\registers[30][2] ), .S1(
        n6449), .D2(n6446), .S2(n670), .D3(\registers[20][2] ), .S3(n6443), 
        .Z(n1015) );
  HS65_LH_MX41X7 U2643 ( .D0(n6452), .S0(n765), .D1(\registers[30][3] ), .S1(
        n6450), .D2(n6446), .S2(n669), .D3(\registers[20][3] ), .S3(n6444), 
        .Z(n973) );
  HS65_LH_MX41X7 U2644 ( .D0(n6453), .S0(n764), .D1(\registers[30][4] ), .S1(
        n6450), .D2(n6447), .S2(n668), .D3(\registers[20][4] ), .S3(n6444), 
        .Z(n959) );
  HS65_LH_MX41X7 U2645 ( .D0(n6453), .S0(n763), .D1(\registers[30][5] ), .S1(
        n6450), .D2(n6447), .S2(n667), .D3(\registers[20][5] ), .S3(n6444), 
        .Z(n945) );
  HS65_LH_MX41X7 U2646 ( .D0(n6453), .S0(n762), .D1(\registers[30][6] ), .S1(
        n6450), .D2(n6447), .S2(n666), .D3(\registers[20][6] ), .S3(n6444), 
        .Z(n931) );
  HS65_LH_MX41X7 U2647 ( .D0(n6453), .S0(n761), .D1(\registers[30][7] ), .S1(
        n6450), .D2(n6447), .S2(n665), .D3(\registers[20][7] ), .S3(n6444), 
        .Z(n917) );
  HS65_LH_MX41X7 U2648 ( .D0(n6453), .S0(n760), .D1(\registers[30][8] ), .S1(
        n6450), .D2(n6447), .S2(n664), .D3(\registers[20][8] ), .S3(n6444), 
        .Z(n903) );
  HS65_LH_MX41X7 U2649 ( .D0(n6453), .S0(n759), .D1(\registers[30][9] ), .S1(
        n6450), .D2(n6447), .S2(n663), .D3(\registers[20][9] ), .S3(n6444), 
        .Z(n873) );
  HS65_LH_MX41X7 U2650 ( .D0(n6451), .S0(n757), .D1(\registers[30][11] ), .S1(
        n6448), .D2(n6445), .S2(n661), .D3(\registers[20][11] ), .S3(n6442), 
        .Z(n1295) );
  HS65_LH_MX41X7 U2651 ( .D0(n6451), .S0(n756), .D1(\registers[30][12] ), .S1(
        n6448), .D2(n6445), .S2(n660), .D3(\registers[20][12] ), .S3(n6442), 
        .Z(n1281) );
  HS65_LH_MX41X7 U2652 ( .D0(n6451), .S0(n755), .D1(\registers[30][13] ), .S1(
        n6448), .D2(n6445), .S2(n659), .D3(\registers[20][13] ), .S3(n6442), 
        .Z(n1267) );
  HS65_LH_MX41X7 U2653 ( .D0(n6451), .S0(n754), .D1(\registers[30][14] ), .S1(
        n6448), .D2(n6445), .S2(n658), .D3(\registers[20][14] ), .S3(n6442), 
        .Z(n1253) );
  HS65_LH_MX41X7 U2654 ( .D0(n6451), .S0(n753), .D1(\registers[30][15] ), .S1(
        n6448), .D2(n6445), .S2(n657), .D3(\registers[20][15] ), .S3(n6442), 
        .Z(n1239) );
  HS65_LH_MX41X7 U2655 ( .D0(n6451), .S0(n752), .D1(\registers[30][16] ), .S1(
        n6448), .D2(n6445), .S2(n656), .D3(\registers[20][16] ), .S3(n6442), 
        .Z(n1225) );
  HS65_LH_MX41X7 U2656 ( .D0(n6451), .S0(n751), .D1(\registers[30][17] ), .S1(
        n6448), .D2(n6445), .S2(n655), .D3(\registers[20][17] ), .S3(n6442), 
        .Z(n1211) );
  HS65_LH_MX41X7 U2657 ( .D0(n6451), .S0(n750), .D1(\registers[30][18] ), .S1(
        n6448), .D2(n6445), .S2(n654), .D3(\registers[20][18] ), .S3(n6442), 
        .Z(n1197) );
  HS65_LH_MX41X7 U2658 ( .D0(n6451), .S0(n749), .D1(\registers[30][19] ), .S1(
        n6448), .D2(n6445), .S2(n653), .D3(\registers[20][19] ), .S3(n6442), 
        .Z(n1183) );
  HS65_LH_MX41X7 U2659 ( .D0(n6451), .S0(n748), .D1(\registers[30][20] ), .S1(
        n6449), .D2(n6445), .S2(n652), .D3(\registers[20][20] ), .S3(n6443), 
        .Z(n1155) );
  HS65_LH_MX41X7 U2660 ( .D0(n6452), .S0(n747), .D1(\registers[30][21] ), .S1(
        n6449), .D2(n6446), .S2(n651), .D3(\registers[20][21] ), .S3(n6443), 
        .Z(n1141) );
  HS65_LH_MX41X7 U2661 ( .D0(n6452), .S0(n746), .D1(\registers[30][22] ), .S1(
        n6449), .D2(n6446), .S2(n650), .D3(\registers[20][22] ), .S3(n6443), 
        .Z(n1127) );
  HS65_LH_MX41X7 U2662 ( .D0(n6452), .S0(n745), .D1(\registers[30][23] ), .S1(
        n6449), .D2(n6446), .S2(n649), .D3(\registers[20][23] ), .S3(n6443), 
        .Z(n1113) );
  HS65_LH_MX41X7 U2663 ( .D0(n6452), .S0(n744), .D1(\registers[30][24] ), .S1(
        n6449), .D2(n6446), .S2(n648), .D3(\registers[20][24] ), .S3(n6443), 
        .Z(n1099) );
  HS65_LH_MX41X7 U2664 ( .D0(n6452), .S0(n743), .D1(\registers[30][25] ), .S1(
        n6449), .D2(n6446), .S2(n647), .D3(\registers[20][25] ), .S3(n6443), 
        .Z(n1085) );
  HS65_LH_MX41X7 U2665 ( .D0(n6452), .S0(n742), .D1(\registers[30][26] ), .S1(
        n6449), .D2(n6446), .S2(n646), .D3(\registers[20][26] ), .S3(n6443), 
        .Z(n1071) );
  HS65_LH_MX41X7 U2666 ( .D0(n6452), .S0(n741), .D1(\registers[30][27] ), .S1(
        n6449), .D2(n6446), .S2(n645), .D3(\registers[20][27] ), .S3(n6443), 
        .Z(n1057) );
  HS65_LH_MX41X7 U2667 ( .D0(n6452), .S0(n740), .D1(\registers[30][28] ), .S1(
        n6449), .D2(n6446), .S2(n644), .D3(\registers[20][28] ), .S3(n6443), 
        .Z(n1043) );
  HS65_LH_MX41X7 U2668 ( .D0(n6452), .S0(n739), .D1(\registers[30][29] ), .S1(
        n6449), .D2(n6446), .S2(n643), .D3(\registers[20][29] ), .S3(n6443), 
        .Z(n1029) );
  HS65_LH_MX41X7 U2669 ( .D0(n6452), .S0(n738), .D1(\registers[30][30] ), .S1(
        n6449), .D2(n6446), .S2(n642), .D3(\registers[20][30] ), .S3(n6443), 
        .Z(n1001) );
  HS65_LH_MX41X7 U2670 ( .D0(n6452), .S0(n737), .D1(\registers[30][31] ), .S1(
        n6450), .D2(n6446), .S2(n641), .D3(\registers[20][31] ), .S3(n6444), 
        .Z(n987) );
  HS65_LH_MX41X7 U2671 ( .D0(\registers[2][0] ), .S0(n6499), .D1(n6496), .S1(
        n640), .D2(n6493), .S2(n576), .D3(\registers[23][0] ), .S3(n6490), .Z(
        n1318) );
  HS65_LH_IVX9 U2672 ( .A(n160), .Z(n576) );
  HS65_LH_MX41X7 U2673 ( .D0(\registers[2][1] ), .S0(n6499), .D1(n6496), .S1(
        n639), .D2(n6493), .S2(n575), .D3(\registers[23][1] ), .S3(n6490), .Z(
        n1164) );
  HS65_LH_IVX9 U2674 ( .A(n159), .Z(n575) );
  HS65_LH_MX41X7 U2675 ( .D0(\registers[2][2] ), .S0(n6500), .D1(n6497), .S1(
        n638), .D2(n6494), .S2(n574), .D3(\registers[23][2] ), .S3(n6491), .Z(
        n1010) );
  HS65_LH_IVX9 U2676 ( .A(n158), .Z(n574) );
  HS65_LH_MX41X7 U2677 ( .D0(\registers[2][3] ), .S0(n6501), .D1(n6498), .S1(
        n637), .D2(n6494), .S2(n573), .D3(\registers[23][3] ), .S3(n6492), .Z(
        n968) );
  HS65_LH_IVX9 U2678 ( .A(n157), .Z(n573) );
  HS65_LH_MX41X7 U2679 ( .D0(\registers[2][4] ), .S0(n6501), .D1(n6498), .S1(
        n636), .D2(n6495), .S2(n572), .D3(\registers[23][4] ), .S3(n6492), .Z(
        n954) );
  HS65_LH_IVX9 U2680 ( .A(n156), .Z(n572) );
  HS65_LH_MX41X7 U2681 ( .D0(\registers[2][5] ), .S0(n6501), .D1(n6498), .S1(
        n635), .D2(n6495), .S2(n571), .D3(\registers[23][5] ), .S3(n6492), .Z(
        n940) );
  HS65_LH_IVX9 U2682 ( .A(n155), .Z(n571) );
  HS65_LH_MX41X7 U2683 ( .D0(\registers[2][6] ), .S0(n6501), .D1(n6498), .S1(
        n634), .D2(n6495), .S2(n570), .D3(\registers[23][6] ), .S3(n6492), .Z(
        n926) );
  HS65_LH_IVX9 U2684 ( .A(n154), .Z(n570) );
  HS65_LH_MX41X7 U2685 ( .D0(\registers[2][7] ), .S0(n6501), .D1(n6498), .S1(
        n633), .D2(n6495), .S2(n569), .D3(\registers[23][7] ), .S3(n6492), .Z(
        n912) );
  HS65_LH_IVX9 U2686 ( .A(n153), .Z(n569) );
  HS65_LH_MX41X7 U2687 ( .D0(\registers[2][8] ), .S0(n6501), .D1(n6498), .S1(
        n632), .D2(n6495), .S2(n568), .D3(\registers[23][8] ), .S3(n6492), .Z(
        n898) );
  HS65_LH_IVX9 U2688 ( .A(n152), .Z(n568) );
  HS65_LH_MX41X7 U2689 ( .D0(\registers[2][9] ), .S0(n6501), .D1(n6498), .S1(
        n631), .D2(n6495), .S2(n567), .D3(\registers[23][9] ), .S3(n6492), .Z(
        n853) );
  HS65_LH_IVX9 U2690 ( .A(n151), .Z(n567) );
  HS65_LH_MX41X7 U2691 ( .D0(\registers[2][10] ), .S0(n6499), .D1(n6496), .S1(
        n630), .D2(n6493), .S2(n566), .D3(\registers[23][10] ), .S3(n6490), 
        .Z(n1304) );
  HS65_LH_IVX9 U2692 ( .A(n150), .Z(n566) );
  HS65_LH_MX41X7 U2693 ( .D0(\registers[2][11] ), .S0(n6499), .D1(n6496), .S1(
        n629), .D2(n6493), .S2(n565), .D3(\registers[23][11] ), .S3(n6490), 
        .Z(n1290) );
  HS65_LH_IVX9 U2694 ( .A(n149), .Z(n565) );
  HS65_LH_MX41X7 U2695 ( .D0(\registers[2][12] ), .S0(n6499), .D1(n6496), .S1(
        n628), .D2(n6493), .S2(n564), .D3(\registers[23][12] ), .S3(n6490), 
        .Z(n1276) );
  HS65_LH_IVX9 U2696 ( .A(n148), .Z(n564) );
  HS65_LH_MX41X7 U2697 ( .D0(\registers[2][13] ), .S0(n6499), .D1(n6496), .S1(
        n627), .D2(n6493), .S2(n563), .D3(\registers[23][13] ), .S3(n6490), 
        .Z(n1262) );
  HS65_LH_IVX9 U2698 ( .A(n147), .Z(n563) );
  HS65_LH_MX41X7 U2699 ( .D0(\registers[2][14] ), .S0(n6499), .D1(n6496), .S1(
        n626), .D2(n6493), .S2(n562), .D3(\registers[23][14] ), .S3(n6490), 
        .Z(n1248) );
  HS65_LH_IVX9 U2700 ( .A(n146), .Z(n562) );
  HS65_LH_MX41X7 U2701 ( .D0(\registers[2][15] ), .S0(n6499), .D1(n6496), .S1(
        n625), .D2(n6493), .S2(n561), .D3(\registers[23][15] ), .S3(n6490), 
        .Z(n1234) );
  HS65_LH_IVX9 U2702 ( .A(n145), .Z(n561) );
  HS65_LH_MX41X7 U2703 ( .D0(\registers[2][16] ), .S0(n6499), .D1(n6496), .S1(
        n624), .D2(n6493), .S2(n560), .D3(\registers[23][16] ), .S3(n6490), 
        .Z(n1220) );
  HS65_LH_IVX9 U2704 ( .A(n144), .Z(n560) );
  HS65_LH_MX41X7 U2705 ( .D0(\registers[2][17] ), .S0(n6499), .D1(n6496), .S1(
        n623), .D2(n6493), .S2(n559), .D3(\registers[23][17] ), .S3(n6490), 
        .Z(n1206) );
  HS65_LH_IVX9 U2706 ( .A(n143), .Z(n559) );
  HS65_LH_MX41X7 U2707 ( .D0(\registers[2][18] ), .S0(n6499), .D1(n6496), .S1(
        n622), .D2(n6493), .S2(n558), .D3(\registers[23][18] ), .S3(n6490), 
        .Z(n1192) );
  HS65_LH_IVX9 U2708 ( .A(n142), .Z(n558) );
  HS65_LH_MX41X7 U2709 ( .D0(\registers[2][19] ), .S0(n6499), .D1(n6496), .S1(
        n621), .D2(n6493), .S2(n557), .D3(\registers[23][19] ), .S3(n6490), 
        .Z(n1178) );
  HS65_LH_IVX9 U2710 ( .A(n141), .Z(n557) );
  HS65_LH_MX41X7 U2711 ( .D0(\registers[2][20] ), .S0(n6500), .D1(n6497), .S1(
        n620), .D2(n6493), .S2(n556), .D3(\registers[23][20] ), .S3(n6491), 
        .Z(n1150) );
  HS65_LH_IVX9 U2712 ( .A(n140), .Z(n556) );
  HS65_LH_MX41X7 U2713 ( .D0(\registers[2][21] ), .S0(n6500), .D1(n6497), .S1(
        n619), .D2(n6494), .S2(n555), .D3(\registers[23][21] ), .S3(n6491), 
        .Z(n1136) );
  HS65_LH_IVX9 U2714 ( .A(n139), .Z(n555) );
  HS65_LH_MX41X7 U2715 ( .D0(\registers[2][22] ), .S0(n6500), .D1(n6497), .S1(
        n618), .D2(n6494), .S2(n554), .D3(\registers[23][22] ), .S3(n6491), 
        .Z(n1122) );
  HS65_LH_IVX9 U2716 ( .A(n138), .Z(n554) );
  HS65_LH_MX41X7 U2717 ( .D0(\registers[2][23] ), .S0(n6500), .D1(n6497), .S1(
        n617), .D2(n6494), .S2(n553), .D3(\registers[23][23] ), .S3(n6491), 
        .Z(n1108) );
  HS65_LH_IVX9 U2718 ( .A(n137), .Z(n553) );
  HS65_LH_MX41X7 U2719 ( .D0(\registers[2][24] ), .S0(n6500), .D1(n6497), .S1(
        n616), .D2(n6494), .S2(n552), .D3(\registers[23][24] ), .S3(n6491), 
        .Z(n1094) );
  HS65_LH_IVX9 U2720 ( .A(n136), .Z(n552) );
  HS65_LH_MX41X7 U2721 ( .D0(\registers[2][25] ), .S0(n6500), .D1(n6497), .S1(
        n615), .D2(n6494), .S2(n551), .D3(\registers[23][25] ), .S3(n6491), 
        .Z(n1080) );
  HS65_LH_IVX9 U2722 ( .A(n135), .Z(n551) );
  HS65_LH_MX41X7 U2723 ( .D0(\registers[2][26] ), .S0(n6500), .D1(n6497), .S1(
        n614), .D2(n6494), .S2(n550), .D3(\registers[23][26] ), .S3(n6491), 
        .Z(n1066) );
  HS65_LH_IVX9 U2724 ( .A(n134), .Z(n550) );
  HS65_LH_MX41X7 U2725 ( .D0(\registers[2][27] ), .S0(n6500), .D1(n6497), .S1(
        n613), .D2(n6494), .S2(n549), .D3(\registers[23][27] ), .S3(n6491), 
        .Z(n1052) );
  HS65_LH_IVX9 U2726 ( .A(n133), .Z(n549) );
  HS65_LH_MX41X7 U2727 ( .D0(\registers[2][28] ), .S0(n6500), .D1(n6497), .S1(
        n612), .D2(n6494), .S2(n548), .D3(\registers[23][28] ), .S3(n6491), 
        .Z(n1038) );
  HS65_LH_IVX9 U2728 ( .A(n132), .Z(n548) );
  HS65_LH_MX41X7 U2729 ( .D0(\registers[2][29] ), .S0(n6500), .D1(n6497), .S1(
        n611), .D2(n6494), .S2(n547), .D3(\registers[23][29] ), .S3(n6491), 
        .Z(n1024) );
  HS65_LH_IVX9 U2730 ( .A(n131), .Z(n547) );
  HS65_LH_MX41X7 U2731 ( .D0(\registers[2][30] ), .S0(n6500), .D1(n6497), .S1(
        n610), .D2(n6494), .S2(n546), .D3(\registers[23][30] ), .S3(n6491), 
        .Z(n996) );
  HS65_LH_IVX9 U2732 ( .A(n130), .Z(n546) );
  HS65_LH_MX41X7 U2733 ( .D0(\registers[2][31] ), .S0(n6501), .D1(n6498), .S1(
        n609), .D2(n6494), .S2(n545), .D3(\registers[23][31] ), .S3(n6492), 
        .Z(n982) );
  HS65_LH_IVX9 U2734 ( .A(n129), .Z(n545) );
  HS65_LH_MX41X7 U2735 ( .D0(n6394), .S0(\registers[7][0] ), .D1(n6391), .S1(
        \registers[4][0] ), .D2(n6388), .S2(\registers[5][0] ), .D3(n6385), 
        .S3(\registers[1][0] ), .Z(n2800) );
  HS65_LH_MX41X7 U2736 ( .D0(n6394), .S0(\registers[7][1] ), .D1(n6391), .S1(
        \registers[4][1] ), .D2(n6388), .S2(\registers[5][1] ), .D3(n6385), 
        .S3(\registers[1][1] ), .Z(n2646) );
  HS65_LH_MX41X7 U2737 ( .D0(n6395), .S0(\registers[7][2] ), .D1(n6392), .S1(
        \registers[4][2] ), .D2(n6389), .S2(\registers[5][2] ), .D3(n6386), 
        .S3(\registers[1][2] ), .Z(n2492) );
  HS65_LH_MX41X7 U2738 ( .D0(n6395), .S0(\registers[7][3] ), .D1(n6393), .S1(
        \registers[4][3] ), .D2(n6389), .S2(\registers[5][3] ), .D3(n6387), 
        .S3(\registers[1][3] ), .Z(n2450) );
  HS65_LH_MX41X7 U2739 ( .D0(n6396), .S0(\registers[7][4] ), .D1(n6393), .S1(
        \registers[4][4] ), .D2(n6390), .S2(\registers[5][4] ), .D3(n6387), 
        .S3(\registers[1][4] ), .Z(n2436) );
  HS65_LH_MX41X7 U2740 ( .D0(n6396), .S0(\registers[7][5] ), .D1(n6393), .S1(
        \registers[4][5] ), .D2(n6390), .S2(\registers[5][5] ), .D3(n6387), 
        .S3(\registers[1][5] ), .Z(n1430) );
  HS65_LH_MX41X7 U2741 ( .D0(n6396), .S0(\registers[7][6] ), .D1(n6393), .S1(
        \registers[4][6] ), .D2(n6390), .S2(\registers[5][6] ), .D3(n6387), 
        .S3(\registers[1][6] ), .Z(n1416) );
  HS65_LH_MX41X7 U2742 ( .D0(n6396), .S0(\registers[7][7] ), .D1(n6393), .S1(
        \registers[4][7] ), .D2(n6390), .S2(\registers[5][7] ), .D3(n6387), 
        .S3(\registers[1][7] ), .Z(n1402) );
  HS65_LH_MX41X7 U2743 ( .D0(n6396), .S0(\registers[7][8] ), .D1(n6393), .S1(
        \registers[4][8] ), .D2(n6390), .S2(\registers[5][8] ), .D3(n6387), 
        .S3(\registers[1][8] ), .Z(n1388) );
  HS65_LH_MX41X7 U2744 ( .D0(n6396), .S0(\registers[7][9] ), .D1(n6393), .S1(
        \registers[4][9] ), .D2(n6390), .S2(\registers[5][9] ), .D3(n6387), 
        .S3(\registers[1][9] ), .Z(n1343) );
  HS65_LH_MX41X7 U2745 ( .D0(n6394), .S0(\registers[7][10] ), .D1(n6391), .S1(
        \registers[4][10] ), .D2(n6388), .S2(\registers[5][10] ), .D3(n6385), 
        .S3(\registers[1][10] ), .Z(n2786) );
  HS65_LH_MX41X7 U2746 ( .D0(n6394), .S0(\registers[7][11] ), .D1(n6391), .S1(
        \registers[4][11] ), .D2(n6388), .S2(\registers[5][11] ), .D3(n6385), 
        .S3(\registers[1][11] ), .Z(n2772) );
  HS65_LH_MX41X7 U2747 ( .D0(n6394), .S0(\registers[7][12] ), .D1(n6391), .S1(
        \registers[4][12] ), .D2(n6388), .S2(\registers[5][12] ), .D3(n6385), 
        .S3(\registers[1][12] ), .Z(n2758) );
  HS65_LH_MX41X7 U2748 ( .D0(n6394), .S0(\registers[7][13] ), .D1(n6391), .S1(
        \registers[4][13] ), .D2(n6388), .S2(\registers[5][13] ), .D3(n6385), 
        .S3(\registers[1][13] ), .Z(n2744) );
  HS65_LH_MX41X7 U2749 ( .D0(n6394), .S0(\registers[7][14] ), .D1(n6391), .S1(
        \registers[4][14] ), .D2(n6388), .S2(\registers[5][14] ), .D3(n6385), 
        .S3(\registers[1][14] ), .Z(n2730) );
  HS65_LH_MX41X7 U2750 ( .D0(n6394), .S0(\registers[7][15] ), .D1(n6391), .S1(
        \registers[4][15] ), .D2(n6388), .S2(\registers[5][15] ), .D3(n6385), 
        .S3(\registers[1][15] ), .Z(n2716) );
  HS65_LH_MX41X7 U2751 ( .D0(n6394), .S0(\registers[7][16] ), .D1(n6391), .S1(
        \registers[4][16] ), .D2(n6388), .S2(\registers[5][16] ), .D3(n6385), 
        .S3(\registers[1][16] ), .Z(n2702) );
  HS65_LH_MX41X7 U2752 ( .D0(n6394), .S0(\registers[7][17] ), .D1(n6391), .S1(
        \registers[4][17] ), .D2(n6388), .S2(\registers[5][17] ), .D3(n6385), 
        .S3(\registers[1][17] ), .Z(n2688) );
  HS65_LH_MX41X7 U2753 ( .D0(n6394), .S0(\registers[7][18] ), .D1(n6391), .S1(
        \registers[4][18] ), .D2(n6388), .S2(\registers[5][18] ), .D3(n6385), 
        .S3(\registers[1][18] ), .Z(n2674) );
  HS65_LH_MX41X7 U2754 ( .D0(n6394), .S0(\registers[7][19] ), .D1(n6391), .S1(
        \registers[4][19] ), .D2(n6388), .S2(\registers[5][19] ), .D3(n6385), 
        .S3(\registers[1][19] ), .Z(n2660) );
  HS65_LH_MX41X7 U2755 ( .D0(n6394), .S0(\registers[7][20] ), .D1(n6392), .S1(
        \registers[4][20] ), .D2(n6388), .S2(\registers[5][20] ), .D3(n6386), 
        .S3(\registers[1][20] ), .Z(n2632) );
  HS65_LH_MX41X7 U2756 ( .D0(n6395), .S0(\registers[7][21] ), .D1(n6392), .S1(
        \registers[4][21] ), .D2(n6389), .S2(\registers[5][21] ), .D3(n6386), 
        .S3(\registers[1][21] ), .Z(n2618) );
  HS65_LH_MX41X7 U2757 ( .D0(n6395), .S0(\registers[7][22] ), .D1(n6392), .S1(
        \registers[4][22] ), .D2(n6389), .S2(\registers[5][22] ), .D3(n6386), 
        .S3(\registers[1][22] ), .Z(n2604) );
  HS65_LH_MX41X7 U2758 ( .D0(n6395), .S0(\registers[7][23] ), .D1(n6392), .S1(
        \registers[4][23] ), .D2(n6389), .S2(\registers[5][23] ), .D3(n6386), 
        .S3(\registers[1][23] ), .Z(n2590) );
  HS65_LH_MX41X7 U2759 ( .D0(n6395), .S0(\registers[7][24] ), .D1(n6392), .S1(
        \registers[4][24] ), .D2(n6389), .S2(\registers[5][24] ), .D3(n6386), 
        .S3(\registers[1][24] ), .Z(n2576) );
  HS65_LH_MX41X7 U2760 ( .D0(n6395), .S0(\registers[7][25] ), .D1(n6392), .S1(
        \registers[4][25] ), .D2(n6389), .S2(\registers[5][25] ), .D3(n6386), 
        .S3(\registers[1][25] ), .Z(n2562) );
  HS65_LH_MX41X7 U2761 ( .D0(n6395), .S0(\registers[7][26] ), .D1(n6392), .S1(
        \registers[4][26] ), .D2(n6389), .S2(\registers[5][26] ), .D3(n6386), 
        .S3(\registers[1][26] ), .Z(n2548) );
  HS65_LH_MX41X7 U2762 ( .D0(n6395), .S0(\registers[7][27] ), .D1(n6392), .S1(
        \registers[4][27] ), .D2(n6389), .S2(\registers[5][27] ), .D3(n6386), 
        .S3(\registers[1][27] ), .Z(n2534) );
  HS65_LH_MX41X7 U2763 ( .D0(n6395), .S0(\registers[7][28] ), .D1(n6392), .S1(
        \registers[4][28] ), .D2(n6389), .S2(\registers[5][28] ), .D3(n6386), 
        .S3(\registers[1][28] ), .Z(n2520) );
  HS65_LH_MX41X7 U2764 ( .D0(n6395), .S0(\registers[7][29] ), .D1(n6392), .S1(
        \registers[4][29] ), .D2(n6389), .S2(\registers[5][29] ), .D3(n6386), 
        .S3(\registers[1][29] ), .Z(n2506) );
  HS65_LH_MX41X7 U2765 ( .D0(n6395), .S0(\registers[7][30] ), .D1(n6392), .S1(
        \registers[4][30] ), .D2(n6389), .S2(\registers[5][30] ), .D3(n6386), 
        .S3(\registers[1][30] ), .Z(n2478) );
  HS65_LH_MX41X7 U2766 ( .D0(n6395), .S0(\registers[7][31] ), .D1(n6393), .S1(
        \registers[4][31] ), .D2(n6389), .S2(\registers[5][31] ), .D3(n6387), 
        .S3(\registers[1][31] ), .Z(n2464) );
  HS65_LH_MX41X7 U2767 ( .D0(\registers[22][0] ), .S0(n6439), .D1(
        \registers[21][0] ), .S1(n6436), .D2(\registers[19][0] ), .S2(n6433), 
        .D3(n6430), .S3(n608), .Z(n1332) );
  HS65_LH_MX41X7 U2768 ( .D0(\registers[22][1] ), .S0(n6439), .D1(
        \registers[21][1] ), .S1(n6436), .D2(\registers[19][1] ), .S2(n6433), 
        .D3(n6430), .S3(n607), .Z(n1168) );
  HS65_LH_MX41X7 U2769 ( .D0(\registers[22][2] ), .S0(n6440), .D1(
        \registers[21][2] ), .S1(n6437), .D2(\registers[19][2] ), .S2(n6434), 
        .D3(n6431), .S3(n606), .Z(n1014) );
  HS65_LH_MX41X7 U2770 ( .D0(\registers[22][3] ), .S0(n6441), .D1(
        \registers[21][3] ), .S1(n6438), .D2(\registers[19][3] ), .S2(n6435), 
        .D3(n6432), .S3(n605), .Z(n972) );
  HS65_LH_MX41X7 U2771 ( .D0(\registers[22][4] ), .S0(n6441), .D1(
        \registers[21][4] ), .S1(n6438), .D2(\registers[19][4] ), .S2(n6435), 
        .D3(n6432), .S3(n604), .Z(n958) );
  HS65_LH_MX41X7 U2772 ( .D0(\registers[22][5] ), .S0(n6441), .D1(
        \registers[21][5] ), .S1(n6438), .D2(\registers[19][5] ), .S2(n6435), 
        .D3(n6432), .S3(n603), .Z(n944) );
  HS65_LH_MX41X7 U2773 ( .D0(\registers[22][6] ), .S0(n6441), .D1(
        \registers[21][6] ), .S1(n6438), .D2(\registers[19][6] ), .S2(n6435), 
        .D3(n6432), .S3(n602), .Z(n930) );
  HS65_LH_MX41X7 U2774 ( .D0(\registers[22][7] ), .S0(n6441), .D1(
        \registers[21][7] ), .S1(n6438), .D2(\registers[19][7] ), .S2(n6435), 
        .D3(n6432), .S3(n601), .Z(n916) );
  HS65_LH_MX41X7 U2775 ( .D0(\registers[22][8] ), .S0(n6441), .D1(
        \registers[21][8] ), .S1(n6438), .D2(\registers[19][8] ), .S2(n6435), 
        .D3(n6432), .S3(n600), .Z(n902) );
  HS65_LH_MX41X7 U2776 ( .D0(\registers[22][9] ), .S0(n6441), .D1(
        \registers[21][9] ), .S1(n6438), .D2(\registers[19][9] ), .S2(n6435), 
        .D3(n6432), .S3(n599), .Z(n872) );
  HS65_LH_MX41X7 U2777 ( .D0(\registers[22][11] ), .S0(n6439), .D1(
        \registers[21][11] ), .S1(n6436), .D2(\registers[19][11] ), .S2(n6433), 
        .D3(n6430), .S3(n597), .Z(n1294) );
  HS65_LH_MX41X7 U2778 ( .D0(\registers[22][12] ), .S0(n6439), .D1(
        \registers[21][12] ), .S1(n6436), .D2(\registers[19][12] ), .S2(n6433), 
        .D3(n6430), .S3(n596), .Z(n1280) );
  HS65_LH_MX41X7 U2779 ( .D0(\registers[22][13] ), .S0(n6439), .D1(
        \registers[21][13] ), .S1(n6436), .D2(\registers[19][13] ), .S2(n6433), 
        .D3(n6430), .S3(n595), .Z(n1266) );
  HS65_LH_MX41X7 U2780 ( .D0(\registers[22][14] ), .S0(n6439), .D1(
        \registers[21][14] ), .S1(n6436), .D2(\registers[19][14] ), .S2(n6433), 
        .D3(n6430), .S3(n594), .Z(n1252) );
  HS65_LH_MX41X7 U2781 ( .D0(\registers[22][15] ), .S0(n6439), .D1(
        \registers[21][15] ), .S1(n6436), .D2(\registers[19][15] ), .S2(n6433), 
        .D3(n6430), .S3(n593), .Z(n1238) );
  HS65_LH_MX41X7 U2782 ( .D0(\registers[22][16] ), .S0(n6439), .D1(
        \registers[21][16] ), .S1(n6436), .D2(\registers[19][16] ), .S2(n6433), 
        .D3(n6430), .S3(n592), .Z(n1224) );
  HS65_LH_MX41X7 U2783 ( .D0(\registers[22][17] ), .S0(n6439), .D1(
        \registers[21][17] ), .S1(n6436), .D2(\registers[19][17] ), .S2(n6433), 
        .D3(n6430), .S3(n591), .Z(n1210) );
  HS65_LH_MX41X7 U2784 ( .D0(\registers[22][18] ), .S0(n6439), .D1(
        \registers[21][18] ), .S1(n6436), .D2(\registers[19][18] ), .S2(n6433), 
        .D3(n6430), .S3(n590), .Z(n1196) );
  HS65_LH_MX41X7 U2785 ( .D0(\registers[22][19] ), .S0(n6439), .D1(
        \registers[21][19] ), .S1(n6436), .D2(\registers[19][19] ), .S2(n6433), 
        .D3(n6430), .S3(n589), .Z(n1182) );
  HS65_LH_MX41X7 U2786 ( .D0(\registers[22][20] ), .S0(n6440), .D1(
        \registers[21][20] ), .S1(n6437), .D2(\registers[19][20] ), .S2(n6434), 
        .D3(n6431), .S3(n588), .Z(n1154) );
  HS65_LH_MX41X7 U2787 ( .D0(\registers[22][21] ), .S0(n6440), .D1(
        \registers[21][21] ), .S1(n6437), .D2(\registers[19][21] ), .S2(n6434), 
        .D3(n6431), .S3(n587), .Z(n1140) );
  HS65_LH_MX41X7 U2788 ( .D0(\registers[22][22] ), .S0(n6440), .D1(
        \registers[21][22] ), .S1(n6437), .D2(\registers[19][22] ), .S2(n6434), 
        .D3(n6431), .S3(n586), .Z(n1126) );
  HS65_LH_MX41X7 U2789 ( .D0(\registers[22][23] ), .S0(n6440), .D1(
        \registers[21][23] ), .S1(n6437), .D2(\registers[19][23] ), .S2(n6434), 
        .D3(n6431), .S3(n585), .Z(n1112) );
  HS65_LH_MX41X7 U2790 ( .D0(\registers[22][24] ), .S0(n6440), .D1(
        \registers[21][24] ), .S1(n6437), .D2(\registers[19][24] ), .S2(n6434), 
        .D3(n6431), .S3(n584), .Z(n1098) );
  HS65_LH_MX41X7 U2791 ( .D0(\registers[22][25] ), .S0(n6440), .D1(
        \registers[21][25] ), .S1(n6437), .D2(\registers[19][25] ), .S2(n6434), 
        .D3(n6431), .S3(n583), .Z(n1084) );
  HS65_LH_MX41X7 U2792 ( .D0(\registers[22][26] ), .S0(n6440), .D1(
        \registers[21][26] ), .S1(n6437), .D2(\registers[19][26] ), .S2(n6434), 
        .D3(n6431), .S3(n582), .Z(n1070) );
  HS65_LH_MX41X7 U2793 ( .D0(\registers[22][27] ), .S0(n6440), .D1(
        \registers[21][27] ), .S1(n6437), .D2(\registers[19][27] ), .S2(n6434), 
        .D3(n6431), .S3(n581), .Z(n1056) );
  HS65_LH_MX41X7 U2794 ( .D0(\registers[22][28] ), .S0(n6440), .D1(
        \registers[21][28] ), .S1(n6437), .D2(\registers[19][28] ), .S2(n6434), 
        .D3(n6431), .S3(n580), .Z(n1042) );
  HS65_LH_MX41X7 U2795 ( .D0(\registers[22][29] ), .S0(n6440), .D1(
        \registers[21][29] ), .S1(n6437), .D2(\registers[19][29] ), .S2(n6434), 
        .D3(n6431), .S3(n579), .Z(n1028) );
  HS65_LH_MX41X7 U2796 ( .D0(\registers[22][30] ), .S0(n6440), .D1(
        \registers[21][30] ), .S1(n6437), .D2(\registers[19][30] ), .S2(n6434), 
        .D3(n6431), .S3(n578), .Z(n1000) );
  HS65_LH_MX41X7 U2797 ( .D0(\registers[22][31] ), .S0(n6441), .D1(
        \registers[21][31] ), .S1(n6438), .D2(\registers[19][31] ), .S2(n6435), 
        .D3(n6432), .S3(n577), .Z(n986) );
  HS65_LH_MX41X7 U2798 ( .D0(n6358), .S0(n704), .D1(n6355), .S1(
        \registers[30][0] ), .D2(n6352), .S2(n608), .D3(n6349), .S3(
        \registers[20][0] ), .Z(n2815) );
  HS65_LH_MX41X7 U2799 ( .D0(n6358), .S0(n703), .D1(n6355), .S1(
        \registers[30][1] ), .D2(n6352), .S2(n607), .D3(n6349), .S3(
        \registers[20][1] ), .Z(n2652) );
  HS65_LH_MX41X7 U2800 ( .D0(n6359), .S0(n702), .D1(n6356), .S1(
        \registers[30][2] ), .D2(n6353), .S2(n606), .D3(n6350), .S3(
        \registers[20][2] ), .Z(n2498) );
  HS65_LH_MX41X7 U2801 ( .D0(n6359), .S0(n701), .D1(n6357), .S1(
        \registers[30][3] ), .D2(n6353), .S2(n605), .D3(n6351), .S3(
        \registers[20][3] ), .Z(n2456) );
  HS65_LH_MX41X7 U2802 ( .D0(n6360), .S0(n700), .D1(n6357), .S1(
        \registers[30][4] ), .D2(n6354), .S2(n604), .D3(n6351), .S3(
        \registers[20][4] ), .Z(n2442) );
  HS65_LH_MX41X7 U2803 ( .D0(n6360), .S0(n699), .D1(n6357), .S1(
        \registers[30][5] ), .D2(n6354), .S2(n603), .D3(n6351), .S3(
        \registers[20][5] ), .Z(n2428) );
  HS65_LH_MX41X7 U2804 ( .D0(n6360), .S0(n698), .D1(n6357), .S1(
        \registers[30][6] ), .D2(n6354), .S2(n602), .D3(n6351), .S3(
        \registers[20][6] ), .Z(n1422) );
  HS65_LH_MX41X7 U2805 ( .D0(n6360), .S0(n697), .D1(n6357), .S1(
        \registers[30][7] ), .D2(n6354), .S2(n601), .D3(n6351), .S3(
        \registers[20][7] ), .Z(n1408) );
  HS65_LH_MX41X7 U2806 ( .D0(n6360), .S0(n696), .D1(n6357), .S1(
        \registers[30][8] ), .D2(n6354), .S2(n600), .D3(n6351), .S3(
        \registers[20][8] ), .Z(n1394) );
  HS65_LH_MX41X7 U2807 ( .D0(n6360), .S0(n695), .D1(n6357), .S1(
        \registers[30][9] ), .D2(n6354), .S2(n599), .D3(n6351), .S3(
        \registers[20][9] ), .Z(n1364) );
  HS65_LH_MX41X7 U2808 ( .D0(n6358), .S0(n694), .D1(n6355), .S1(
        \registers[30][10] ), .D2(n6352), .S2(n598), .D3(n6349), .S3(
        \registers[20][10] ), .Z(n2792) );
  HS65_LH_MX41X7 U2809 ( .D0(n6358), .S0(n693), .D1(n6355), .S1(
        \registers[30][11] ), .D2(n6352), .S2(n597), .D3(n6349), .S3(
        \registers[20][11] ), .Z(n2778) );
  HS65_LH_MX41X7 U2810 ( .D0(n6358), .S0(n692), .D1(n6355), .S1(
        \registers[30][12] ), .D2(n6352), .S2(n596), .D3(n6349), .S3(
        \registers[20][12] ), .Z(n2764) );
  HS65_LH_MX41X7 U2811 ( .D0(n6358), .S0(n691), .D1(n6355), .S1(
        \registers[30][13] ), .D2(n6352), .S2(n595), .D3(n6349), .S3(
        \registers[20][13] ), .Z(n2750) );
  HS65_LH_MX41X7 U2812 ( .D0(n6358), .S0(n690), .D1(n6355), .S1(
        \registers[30][14] ), .D2(n6352), .S2(n594), .D3(n6349), .S3(
        \registers[20][14] ), .Z(n2736) );
  HS65_LH_MX41X7 U2813 ( .D0(n6358), .S0(n689), .D1(n6355), .S1(
        \registers[30][15] ), .D2(n6352), .S2(n593), .D3(n6349), .S3(
        \registers[20][15] ), .Z(n2722) );
  HS65_LH_MX41X7 U2814 ( .D0(n6358), .S0(n688), .D1(n6355), .S1(
        \registers[30][16] ), .D2(n6352), .S2(n592), .D3(n6349), .S3(
        \registers[20][16] ), .Z(n2708) );
  HS65_LH_MX41X7 U2815 ( .D0(n6358), .S0(n687), .D1(n6355), .S1(
        \registers[30][17] ), .D2(n6352), .S2(n591), .D3(n6349), .S3(
        \registers[20][17] ), .Z(n2694) );
  HS65_LH_MX41X7 U2816 ( .D0(n6358), .S0(n686), .D1(n6355), .S1(
        \registers[30][18] ), .D2(n6352), .S2(n590), .D3(n6349), .S3(
        \registers[20][18] ), .Z(n2680) );
  HS65_LH_MX41X7 U2817 ( .D0(n6358), .S0(n685), .D1(n6355), .S1(
        \registers[30][19] ), .D2(n6352), .S2(n589), .D3(n6349), .S3(
        \registers[20][19] ), .Z(n2666) );
  HS65_LH_MX41X7 U2818 ( .D0(n6358), .S0(n684), .D1(n6356), .S1(
        \registers[30][20] ), .D2(n6352), .S2(n588), .D3(n6350), .S3(
        \registers[20][20] ), .Z(n2638) );
  HS65_LH_MX41X7 U2819 ( .D0(n6359), .S0(n683), .D1(n6356), .S1(
        \registers[30][21] ), .D2(n6353), .S2(n587), .D3(n6350), .S3(
        \registers[20][21] ), .Z(n2624) );
  HS65_LH_MX41X7 U2820 ( .D0(n6359), .S0(n682), .D1(n6356), .S1(
        \registers[30][22] ), .D2(n6353), .S2(n586), .D3(n6350), .S3(
        \registers[20][22] ), .Z(n2610) );
  HS65_LH_MX41X7 U2821 ( .D0(n6359), .S0(n681), .D1(n6356), .S1(
        \registers[30][23] ), .D2(n6353), .S2(n585), .D3(n6350), .S3(
        \registers[20][23] ), .Z(n2596) );
  HS65_LH_MX41X7 U2822 ( .D0(n6359), .S0(n680), .D1(n6356), .S1(
        \registers[30][24] ), .D2(n6353), .S2(n584), .D3(n6350), .S3(
        \registers[20][24] ), .Z(n2582) );
  HS65_LH_MX41X7 U2823 ( .D0(n6359), .S0(n679), .D1(n6356), .S1(
        \registers[30][25] ), .D2(n6353), .S2(n583), .D3(n6350), .S3(
        \registers[20][25] ), .Z(n2568) );
  HS65_LH_MX41X7 U2824 ( .D0(n6359), .S0(n678), .D1(n6356), .S1(
        \registers[30][26] ), .D2(n6353), .S2(n582), .D3(n6350), .S3(
        \registers[20][26] ), .Z(n2554) );
  HS65_LH_MX41X7 U2825 ( .D0(n6359), .S0(n677), .D1(n6356), .S1(
        \registers[30][27] ), .D2(n6353), .S2(n581), .D3(n6350), .S3(
        \registers[20][27] ), .Z(n2540) );
  HS65_LH_MX41X7 U2826 ( .D0(n6359), .S0(n676), .D1(n6356), .S1(
        \registers[30][28] ), .D2(n6353), .S2(n580), .D3(n6350), .S3(
        \registers[20][28] ), .Z(n2526) );
  HS65_LH_MX41X7 U2827 ( .D0(n6359), .S0(n675), .D1(n6356), .S1(
        \registers[30][29] ), .D2(n6353), .S2(n579), .D3(n6350), .S3(
        \registers[20][29] ), .Z(n2512) );
  HS65_LH_MX41X7 U2828 ( .D0(n6359), .S0(n674), .D1(n6356), .S1(
        \registers[30][30] ), .D2(n6353), .S2(n578), .D3(n6350), .S3(
        \registers[20][30] ), .Z(n2484) );
  HS65_LH_MX41X7 U2829 ( .D0(n6359), .S0(n673), .D1(n6357), .S1(
        \registers[30][31] ), .D2(n6353), .S2(n577), .D3(n6351), .S3(
        \registers[20][31] ), .Z(n2470) );
  HS65_LH_MX41X7 U2830 ( .D0(n6346), .S0(\registers[22][0] ), .D1(n6343), .S1(
        \registers[21][0] ), .D2(n6340), .S2(\registers[23][0] ), .D3(n6337), 
        .S3(\registers[12][0] ), .Z(n2814) );
  HS65_LH_MX41X7 U2831 ( .D0(n6346), .S0(\registers[22][1] ), .D1(n6343), .S1(
        \registers[21][1] ), .D2(n6340), .S2(\registers[23][1] ), .D3(n6337), 
        .S3(\registers[12][1] ), .Z(n2651) );
  HS65_LH_MX41X7 U2832 ( .D0(n6347), .S0(\registers[22][2] ), .D1(n6344), .S1(
        \registers[21][2] ), .D2(n6341), .S2(\registers[23][2] ), .D3(n6338), 
        .S3(\registers[12][2] ), .Z(n2497) );
  HS65_LH_MX41X7 U2833 ( .D0(n6347), .S0(\registers[22][3] ), .D1(n6345), .S1(
        \registers[21][3] ), .D2(n6341), .S2(\registers[23][3] ), .D3(n6339), 
        .S3(\registers[12][3] ), .Z(n2455) );
  HS65_LH_MX41X7 U2834 ( .D0(n6348), .S0(\registers[22][4] ), .D1(n6345), .S1(
        \registers[21][4] ), .D2(n6342), .S2(\registers[23][4] ), .D3(n6339), 
        .S3(\registers[12][4] ), .Z(n2441) );
  HS65_LH_MX41X7 U2835 ( .D0(n6348), .S0(\registers[22][5] ), .D1(n6345), .S1(
        \registers[21][5] ), .D2(n6342), .S2(\registers[23][5] ), .D3(n6339), 
        .S3(\registers[12][5] ), .Z(n2427) );
  HS65_LH_MX41X7 U2836 ( .D0(n6348), .S0(\registers[22][6] ), .D1(n6345), .S1(
        \registers[21][6] ), .D2(n6342), .S2(\registers[23][6] ), .D3(n6339), 
        .S3(\registers[12][6] ), .Z(n1421) );
  HS65_LH_MX41X7 U2837 ( .D0(n6348), .S0(\registers[22][7] ), .D1(n6345), .S1(
        \registers[21][7] ), .D2(n6342), .S2(\registers[23][7] ), .D3(n6339), 
        .S3(\registers[12][7] ), .Z(n1407) );
  HS65_LH_MX41X7 U2838 ( .D0(n6348), .S0(\registers[22][8] ), .D1(n6345), .S1(
        \registers[21][8] ), .D2(n6342), .S2(\registers[23][8] ), .D3(n6339), 
        .S3(\registers[12][8] ), .Z(n1393) );
  HS65_LH_MX41X7 U2839 ( .D0(n6348), .S0(\registers[22][9] ), .D1(n6345), .S1(
        \registers[21][9] ), .D2(n6342), .S2(\registers[23][9] ), .D3(n6339), 
        .S3(\registers[12][9] ), .Z(n1363) );
  HS65_LH_MX41X7 U2840 ( .D0(n6346), .S0(\registers[22][10] ), .D1(n6343), 
        .S1(\registers[21][10] ), .D2(n6340), .S2(\registers[23][10] ), .D3(
        n6337), .S3(\registers[12][10] ), .Z(n2791) );
  HS65_LH_MX41X7 U2841 ( .D0(n6346), .S0(\registers[22][11] ), .D1(n6343), 
        .S1(\registers[21][11] ), .D2(n6340), .S2(\registers[23][11] ), .D3(
        n6337), .S3(\registers[12][11] ), .Z(n2777) );
  HS65_LH_MX41X7 U2842 ( .D0(n6346), .S0(\registers[22][12] ), .D1(n6343), 
        .S1(\registers[21][12] ), .D2(n6340), .S2(\registers[23][12] ), .D3(
        n6337), .S3(\registers[12][12] ), .Z(n2763) );
  HS65_LH_MX41X7 U2843 ( .D0(n6346), .S0(\registers[22][13] ), .D1(n6343), 
        .S1(\registers[21][13] ), .D2(n6340), .S2(\registers[23][13] ), .D3(
        n6337), .S3(\registers[12][13] ), .Z(n2749) );
  HS65_LH_MX41X7 U2844 ( .D0(n6346), .S0(\registers[22][14] ), .D1(n6343), 
        .S1(\registers[21][14] ), .D2(n6340), .S2(\registers[23][14] ), .D3(
        n6337), .S3(\registers[12][14] ), .Z(n2735) );
  HS65_LH_MX41X7 U2845 ( .D0(n6346), .S0(\registers[22][15] ), .D1(n6343), 
        .S1(\registers[21][15] ), .D2(n6340), .S2(\registers[23][15] ), .D3(
        n6337), .S3(\registers[12][15] ), .Z(n2721) );
  HS65_LH_MX41X7 U2846 ( .D0(n6346), .S0(\registers[22][16] ), .D1(n6343), 
        .S1(\registers[21][16] ), .D2(n6340), .S2(\registers[23][16] ), .D3(
        n6337), .S3(\registers[12][16] ), .Z(n2707) );
  HS65_LH_MX41X7 U2847 ( .D0(n6346), .S0(\registers[22][17] ), .D1(n6343), 
        .S1(\registers[21][17] ), .D2(n6340), .S2(\registers[23][17] ), .D3(
        n6337), .S3(\registers[12][17] ), .Z(n2693) );
  HS65_LH_MX41X7 U2848 ( .D0(n6346), .S0(\registers[22][18] ), .D1(n6343), 
        .S1(\registers[21][18] ), .D2(n6340), .S2(\registers[23][18] ), .D3(
        n6337), .S3(\registers[12][18] ), .Z(n2679) );
  HS65_LH_MX41X7 U2849 ( .D0(n6346), .S0(\registers[22][19] ), .D1(n6343), 
        .S1(\registers[21][19] ), .D2(n6340), .S2(\registers[23][19] ), .D3(
        n6337), .S3(\registers[12][19] ), .Z(n2665) );
  HS65_LH_MX41X7 U2850 ( .D0(n6346), .S0(\registers[22][20] ), .D1(n6344), 
        .S1(\registers[21][20] ), .D2(n6340), .S2(\registers[23][20] ), .D3(
        n6338), .S3(\registers[12][20] ), .Z(n2637) );
  HS65_LH_MX41X7 U2851 ( .D0(n6347), .S0(\registers[22][21] ), .D1(n6344), 
        .S1(\registers[21][21] ), .D2(n6341), .S2(\registers[23][21] ), .D3(
        n6338), .S3(\registers[12][21] ), .Z(n2623) );
  HS65_LH_MX41X7 U2852 ( .D0(n6347), .S0(\registers[22][22] ), .D1(n6344), 
        .S1(\registers[21][22] ), .D2(n6341), .S2(\registers[23][22] ), .D3(
        n6338), .S3(\registers[12][22] ), .Z(n2609) );
  HS65_LH_MX41X7 U2853 ( .D0(n6347), .S0(\registers[22][23] ), .D1(n6344), 
        .S1(\registers[21][23] ), .D2(n6341), .S2(\registers[23][23] ), .D3(
        n6338), .S3(\registers[12][23] ), .Z(n2595) );
  HS65_LH_MX41X7 U2854 ( .D0(n6347), .S0(\registers[22][24] ), .D1(n6344), 
        .S1(\registers[21][24] ), .D2(n6341), .S2(\registers[23][24] ), .D3(
        n6338), .S3(\registers[12][24] ), .Z(n2581) );
  HS65_LH_MX41X7 U2855 ( .D0(n6347), .S0(\registers[22][25] ), .D1(n6344), 
        .S1(\registers[21][25] ), .D2(n6341), .S2(\registers[23][25] ), .D3(
        n6338), .S3(\registers[12][25] ), .Z(n2567) );
  HS65_LH_MX41X7 U2856 ( .D0(n6347), .S0(\registers[22][26] ), .D1(n6344), 
        .S1(\registers[21][26] ), .D2(n6341), .S2(\registers[23][26] ), .D3(
        n6338), .S3(\registers[12][26] ), .Z(n2553) );
  HS65_LH_MX41X7 U2857 ( .D0(n6347), .S0(\registers[22][27] ), .D1(n6344), 
        .S1(\registers[21][27] ), .D2(n6341), .S2(\registers[23][27] ), .D3(
        n6338), .S3(\registers[12][27] ), .Z(n2539) );
  HS65_LH_MX41X7 U2858 ( .D0(n6347), .S0(\registers[22][28] ), .D1(n6344), 
        .S1(\registers[21][28] ), .D2(n6341), .S2(\registers[23][28] ), .D3(
        n6338), .S3(\registers[12][28] ), .Z(n2525) );
  HS65_LH_MX41X7 U2859 ( .D0(n6347), .S0(\registers[22][29] ), .D1(n6344), 
        .S1(\registers[21][29] ), .D2(n6341), .S2(\registers[23][29] ), .D3(
        n6338), .S3(\registers[12][29] ), .Z(n2511) );
  HS65_LH_MX41X7 U2860 ( .D0(n6347), .S0(\registers[22][30] ), .D1(n6344), 
        .S1(\registers[21][30] ), .D2(n6341), .S2(\registers[23][30] ), .D3(
        n6338), .S3(\registers[12][30] ), .Z(n2483) );
  HS65_LH_MX41X7 U2861 ( .D0(n6347), .S0(\registers[22][31] ), .D1(n6345), 
        .S1(\registers[21][31] ), .D2(n6341), .S2(\registers[23][31] ), .D3(
        n6339), .S3(\registers[12][31] ), .Z(n2469) );
  HS65_LH_IVX9 U2862 ( .A(\regfile_i[ADRREAD1][0] ), .Z(n778) );
  HS65_LH_IVX9 U2863 ( .A(\regfile_i[ADRREAD0][0] ), .Z(n773) );
  HS65_LH_IVX9 U2864 ( .A(\regfile_i[ADRWRITE][2] ), .Z(n812) );
  HS65_LH_MX41X7 U2865 ( .D0(n6406), .S0(n640), .D1(n6403), .S1(
        \registers[2][0] ), .D2(n6400), .S2(\registers[3][0] ), .D3(n6397), 
        .S3(n768), .Z(n2801) );
  HS65_LH_MX41X7 U2866 ( .D0(n6406), .S0(n639), .D1(n6403), .S1(
        \registers[2][1] ), .D2(n6400), .S2(\registers[3][1] ), .D3(n6397), 
        .S3(n767), .Z(n2647) );
  HS65_LH_MX41X7 U2867 ( .D0(n6407), .S0(n638), .D1(n6404), .S1(
        \registers[2][2] ), .D2(n6401), .S2(\registers[3][2] ), .D3(n6398), 
        .S3(n766), .Z(n2493) );
  HS65_LH_MX41X7 U2868 ( .D0(n6406), .S0(n630), .D1(n6403), .S1(
        \registers[2][10] ), .D2(n6400), .S2(\registers[3][10] ), .D3(n6397), 
        .S3(n758), .Z(n2787) );
  HS65_LH_MX41X7 U2869 ( .D0(n6406), .S0(n629), .D1(n6403), .S1(
        \registers[2][11] ), .D2(n6400), .S2(\registers[3][11] ), .D3(n6397), 
        .S3(n757), .Z(n2773) );
  HS65_LH_MX41X7 U2870 ( .D0(n6406), .S0(n628), .D1(n6403), .S1(
        \registers[2][12] ), .D2(n6400), .S2(\registers[3][12] ), .D3(n6397), 
        .S3(n756), .Z(n2759) );
  HS65_LH_MX41X7 U2871 ( .D0(n6406), .S0(n627), .D1(n6403), .S1(
        \registers[2][13] ), .D2(n6400), .S2(\registers[3][13] ), .D3(n6397), 
        .S3(n755), .Z(n2745) );
  HS65_LH_MX41X7 U2872 ( .D0(n6406), .S0(n626), .D1(n6403), .S1(
        \registers[2][14] ), .D2(n6400), .S2(\registers[3][14] ), .D3(n6397), 
        .S3(n754), .Z(n2731) );
  HS65_LH_MX41X7 U2873 ( .D0(n6406), .S0(n625), .D1(n6403), .S1(
        \registers[2][15] ), .D2(n6400), .S2(\registers[3][15] ), .D3(n6397), 
        .S3(n753), .Z(n2717) );
  HS65_LH_MX41X7 U2874 ( .D0(n6406), .S0(n624), .D1(n6403), .S1(
        \registers[2][16] ), .D2(n6400), .S2(\registers[3][16] ), .D3(n6397), 
        .S3(n752), .Z(n2703) );
  HS65_LH_MX41X7 U2875 ( .D0(n6406), .S0(n623), .D1(n6403), .S1(
        \registers[2][17] ), .D2(n6400), .S2(\registers[3][17] ), .D3(n6397), 
        .S3(n751), .Z(n2689) );
  HS65_LH_MX41X7 U2876 ( .D0(n6406), .S0(n622), .D1(n6403), .S1(
        \registers[2][18] ), .D2(n6400), .S2(\registers[3][18] ), .D3(n6397), 
        .S3(n750), .Z(n2675) );
  HS65_LH_MX41X7 U2877 ( .D0(n6406), .S0(n621), .D1(n6403), .S1(
        \registers[2][19] ), .D2(n6400), .S2(\registers[3][19] ), .D3(n6397), 
        .S3(n749), .Z(n2661) );
  HS65_LH_MX41X7 U2878 ( .D0(n6406), .S0(n620), .D1(n6404), .S1(
        \registers[2][20] ), .D2(n6400), .S2(\registers[3][20] ), .D3(n6398), 
        .S3(n748), .Z(n2633) );
  HS65_LH_MX41X7 U2879 ( .D0(n6407), .S0(n619), .D1(n6404), .S1(
        \registers[2][21] ), .D2(n6401), .S2(\registers[3][21] ), .D3(n6398), 
        .S3(n747), .Z(n2619) );
  HS65_LH_MX41X7 U2880 ( .D0(n6407), .S0(n618), .D1(n6404), .S1(
        \registers[2][22] ), .D2(n6401), .S2(\registers[3][22] ), .D3(n6398), 
        .S3(n746), .Z(n2605) );
  HS65_LH_MX41X7 U2881 ( .D0(n6407), .S0(n617), .D1(n6404), .S1(
        \registers[2][23] ), .D2(n6401), .S2(\registers[3][23] ), .D3(n6398), 
        .S3(n745), .Z(n2591) );
  HS65_LH_MX41X7 U2882 ( .D0(n6407), .S0(n616), .D1(n6404), .S1(
        \registers[2][24] ), .D2(n6401), .S2(\registers[3][24] ), .D3(n6398), 
        .S3(n744), .Z(n2577) );
  HS65_LH_MX41X7 U2883 ( .D0(n6407), .S0(n615), .D1(n6404), .S1(
        \registers[2][25] ), .D2(n6401), .S2(\registers[3][25] ), .D3(n6398), 
        .S3(n743), .Z(n2563) );
  HS65_LH_MX41X7 U2884 ( .D0(n6407), .S0(n614), .D1(n6404), .S1(
        \registers[2][26] ), .D2(n6401), .S2(\registers[3][26] ), .D3(n6398), 
        .S3(n742), .Z(n2549) );
  HS65_LH_MX41X7 U2885 ( .D0(n6407), .S0(n613), .D1(n6404), .S1(
        \registers[2][27] ), .D2(n6401), .S2(\registers[3][27] ), .D3(n6398), 
        .S3(n741), .Z(n2535) );
  HS65_LH_MX41X7 U2886 ( .D0(n6407), .S0(n612), .D1(n6404), .S1(
        \registers[2][28] ), .D2(n6401), .S2(\registers[3][28] ), .D3(n6398), 
        .S3(n740), .Z(n2521) );
  HS65_LH_MX41X7 U2887 ( .D0(n6407), .S0(n611), .D1(n6404), .S1(
        \registers[2][29] ), .D2(n6401), .S2(\registers[3][29] ), .D3(n6398), 
        .S3(n739), .Z(n2507) );
  HS65_LH_MX41X7 U2888 ( .D0(n6407), .S0(n610), .D1(n6404), .S1(
        \registers[2][30] ), .D2(n6401), .S2(\registers[3][30] ), .D3(n6398), 
        .S3(n738), .Z(n2479) );
  HS65_LH_IVX9 U2889 ( .A(\regfile_i[WRITE_DATA][0] ), .Z(n846) );
  HS65_LH_IVX9 U2890 ( .A(\regfile_i[WRITE_DATA][1] ), .Z(n845) );
  HS65_LH_IVX9 U2891 ( .A(\regfile_i[WRITE_DATA][2] ), .Z(n844) );
  HS65_LH_IVX9 U2892 ( .A(\regfile_i[WRITE_DATA][3] ), .Z(n843) );
  HS65_LH_IVX9 U2893 ( .A(\regfile_i[WRITE_DATA][4] ), .Z(n842) );
  HS65_LH_IVX9 U2894 ( .A(\regfile_i[WRITE_DATA][5] ), .Z(n841) );
  HS65_LH_IVX9 U2895 ( .A(\regfile_i[WRITE_DATA][6] ), .Z(n840) );
  HS65_LH_IVX9 U2896 ( .A(\regfile_i[WRITE_DATA][7] ), .Z(n839) );
  HS65_LH_IVX9 U2897 ( .A(\regfile_i[WRITE_DATA][8] ), .Z(n838) );
  HS65_LH_IVX9 U2898 ( .A(\regfile_i[WRITE_DATA][9] ), .Z(n837) );
  HS65_LH_IVX9 U2899 ( .A(\regfile_i[WRITE_DATA][10] ), .Z(n836) );
  HS65_LH_IVX9 U2900 ( .A(\regfile_i[WRITE_DATA][11] ), .Z(n835) );
  HS65_LH_IVX9 U2901 ( .A(\regfile_i[WRITE_DATA][12] ), .Z(n834) );
  HS65_LH_IVX9 U2902 ( .A(\regfile_i[WRITE_DATA][13] ), .Z(n833) );
  HS65_LH_IVX9 U2903 ( .A(\regfile_i[WRITE_DATA][14] ), .Z(n832) );
  HS65_LH_IVX9 U2904 ( .A(\regfile_i[WRITE_DATA][15] ), .Z(n831) );
  HS65_LH_IVX9 U2905 ( .A(\regfile_i[WRITE_DATA][16] ), .Z(n830) );
  HS65_LH_IVX9 U2906 ( .A(\regfile_i[WRITE_DATA][17] ), .Z(n829) );
  HS65_LH_IVX9 U2907 ( .A(\regfile_i[WRITE_DATA][18] ), .Z(n828) );
  HS65_LH_IVX9 U2908 ( .A(\regfile_i[WRITE_DATA][19] ), .Z(n827) );
  HS65_LH_IVX9 U2909 ( .A(\regfile_i[WRITE_DATA][20] ), .Z(n826) );
  HS65_LH_IVX9 U2910 ( .A(\regfile_i[WRITE_DATA][21] ), .Z(n825) );
  HS65_LH_IVX9 U2911 ( .A(\regfile_i[WRITE_DATA][22] ), .Z(n824) );
  HS65_LH_IVX9 U2912 ( .A(\regfile_i[WRITE_DATA][23] ), .Z(n823) );
  HS65_LH_IVX9 U2913 ( .A(\regfile_i[WRITE_DATA][24] ), .Z(n822) );
  HS65_LH_IVX9 U2914 ( .A(\regfile_i[WRITE_DATA][25] ), .Z(n821) );
  HS65_LH_IVX9 U2915 ( .A(\regfile_i[WRITE_DATA][26] ), .Z(n820) );
  HS65_LH_IVX9 U2916 ( .A(\regfile_i[WRITE_DATA][27] ), .Z(n819) );
  HS65_LH_IVX9 U2917 ( .A(\regfile_i[WRITE_DATA][28] ), .Z(n818) );
  HS65_LH_IVX9 U2918 ( .A(\regfile_i[WRITE_DATA][29] ), .Z(n817) );
  HS65_LH_IVX9 U2919 ( .A(\regfile_i[WRITE_DATA][30] ), .Z(n816) );
  HS65_LH_IVX9 U2920 ( .A(\regfile_i[WRITE_DATA][31] ), .Z(n815) );
  HS65_LH_MX41X7 U2921 ( .D0(n6407), .S0(n637), .D1(n6405), .S1(
        \registers[2][3] ), .D2(n6401), .S2(\registers[3][3] ), .D3(n6399), 
        .S3(n765), .Z(n2451) );
  HS65_LH_MX41X7 U2922 ( .D0(n6408), .S0(n636), .D1(n6405), .S1(
        \registers[2][4] ), .D2(n6402), .S2(\registers[3][4] ), .D3(n6399), 
        .S3(n764), .Z(n2437) );
  HS65_LH_MX41X7 U2923 ( .D0(n6408), .S0(n635), .D1(n6405), .S1(
        \registers[2][5] ), .D2(n6402), .S2(\registers[3][5] ), .D3(n6399), 
        .S3(n763), .Z(n1431) );
  HS65_LH_MX41X7 U2924 ( .D0(n6408), .S0(n634), .D1(n6405), .S1(
        \registers[2][6] ), .D2(n6402), .S2(\registers[3][6] ), .D3(n6399), 
        .S3(n762), .Z(n1417) );
  HS65_LH_MX41X7 U2925 ( .D0(n6408), .S0(n633), .D1(n6405), .S1(
        \registers[2][7] ), .D2(n6402), .S2(\registers[3][7] ), .D3(n6399), 
        .S3(n761), .Z(n1403) );
  HS65_LH_MX41X7 U2926 ( .D0(n6408), .S0(n632), .D1(n6405), .S1(
        \registers[2][8] ), .D2(n6402), .S2(\registers[3][8] ), .D3(n6399), 
        .S3(n760), .Z(n1389) );
  HS65_LH_MX41X7 U2927 ( .D0(n6408), .S0(n631), .D1(n6405), .S1(
        \registers[2][9] ), .D2(n6402), .S2(\registers[3][9] ), .D3(n6399), 
        .S3(n759), .Z(n1344) );
  HS65_LH_MX41X7 U2928 ( .D0(n6407), .S0(n609), .D1(n6405), .S1(
        \registers[2][31] ), .D2(n6401), .S2(\registers[3][31] ), .D3(n6399), 
        .S3(n737), .Z(n2465) );
  HS65_LH_BFX9 U2929 ( .A(rst_n), .Z(n6536) );
  HS65_LH_IVX9 U2930 ( .A(n96), .Z(n544) );
  HS65_LH_IVX9 U2931 ( .A(n95), .Z(n543) );
  HS65_LH_IVX9 U2932 ( .A(n94), .Z(n542) );
  HS65_LH_IVX9 U2933 ( .A(n93), .Z(n541) );
  HS65_LH_IVX9 U2934 ( .A(n92), .Z(n540) );
  HS65_LH_IVX9 U2935 ( .A(n91), .Z(n539) );
  HS65_LH_IVX9 U2936 ( .A(n90), .Z(n538) );
  HS65_LH_IVX9 U2937 ( .A(n89), .Z(n537) );
  HS65_LH_IVX9 U2938 ( .A(n88), .Z(n536) );
  HS65_LH_IVX9 U2939 ( .A(n87), .Z(n535) );
  HS65_LH_IVX9 U2940 ( .A(n86), .Z(n534) );
  HS65_LH_IVX9 U2941 ( .A(n85), .Z(n533) );
  HS65_LH_IVX9 U2942 ( .A(n84), .Z(n532) );
  HS65_LH_IVX9 U2943 ( .A(n83), .Z(n531) );
  HS65_LH_IVX9 U2944 ( .A(n82), .Z(n530) );
  HS65_LH_IVX9 U2945 ( .A(n81), .Z(n529) );
  HS65_LH_IVX9 U2946 ( .A(n80), .Z(n528) );
  HS65_LH_IVX9 U2947 ( .A(n79), .Z(n527) );
  HS65_LH_IVX9 U2948 ( .A(n78), .Z(n526) );
  HS65_LH_IVX9 U2949 ( .A(n77), .Z(n525) );
  HS65_LH_IVX9 U2950 ( .A(n76), .Z(n524) );
  HS65_LH_IVX9 U2951 ( .A(n75), .Z(n523) );
  HS65_LH_IVX9 U2952 ( .A(n74), .Z(n522) );
  HS65_LH_IVX9 U2953 ( .A(n73), .Z(n521) );
  HS65_LH_IVX9 U2954 ( .A(n72), .Z(n520) );
  HS65_LH_IVX9 U2955 ( .A(n71), .Z(n519) );
  HS65_LH_IVX9 U2956 ( .A(n70), .Z(n518) );
  HS65_LH_IVX9 U2957 ( .A(n69), .Z(n517) );
  HS65_LH_IVX9 U2958 ( .A(n68), .Z(n516) );
  HS65_LH_IVX9 U2959 ( .A(n67), .Z(n515) );
  HS65_LH_IVX9 U2960 ( .A(n66), .Z(n514) );
  HS65_LH_IVX9 U2961 ( .A(n65), .Z(n513) );
  HS65_LH_IVX9 U2962 ( .A(n32), .Z(n704) );
  HS65_LH_IVX9 U2963 ( .A(n31), .Z(n703) );
  HS65_LH_IVX9 U2964 ( .A(n30), .Z(n702) );
  HS65_LH_IVX9 U2965 ( .A(n29), .Z(n701) );
  HS65_LH_IVX9 U2966 ( .A(n28), .Z(n700) );
  HS65_LH_IVX9 U2967 ( .A(n27), .Z(n699) );
  HS65_LH_IVX9 U2968 ( .A(n26), .Z(n698) );
  HS65_LH_IVX9 U2969 ( .A(n25), .Z(n697) );
  HS65_LH_IVX9 U2970 ( .A(n24), .Z(n696) );
  HS65_LH_IVX9 U2971 ( .A(n23), .Z(n695) );
  HS65_LH_IVX9 U2972 ( .A(n22), .Z(n694) );
  HS65_LH_IVX9 U2973 ( .A(n21), .Z(n693) );
  HS65_LH_IVX9 U2974 ( .A(n20), .Z(n692) );
  HS65_LH_IVX9 U2975 ( .A(n19), .Z(n691) );
  HS65_LH_IVX9 U2976 ( .A(n18), .Z(n690) );
  HS65_LH_IVX9 U2977 ( .A(n17), .Z(n689) );
  HS65_LH_IVX9 U2978 ( .A(n16), .Z(n688) );
  HS65_LH_IVX9 U2979 ( .A(n15), .Z(n687) );
  HS65_LH_IVX9 U2980 ( .A(n14), .Z(n686) );
  HS65_LH_IVX9 U2981 ( .A(n13), .Z(n685) );
  HS65_LH_IVX9 U2982 ( .A(n12), .Z(n684) );
  HS65_LH_IVX9 U2983 ( .A(n11), .Z(n683) );
  HS65_LH_IVX9 U2984 ( .A(n10), .Z(n682) );
  HS65_LH_IVX9 U2985 ( .A(n9), .Z(n681) );
  HS65_LH_IVX9 U2986 ( .A(n8), .Z(n680) );
  HS65_LH_IVX9 U2987 ( .A(n7), .Z(n679) );
  HS65_LH_IVX9 U2988 ( .A(n6), .Z(n678) );
  HS65_LH_IVX9 U2989 ( .A(n5), .Z(n677) );
  HS65_LH_IVX9 U2990 ( .A(n4), .Z(n676) );
  HS65_LH_IVX9 U2991 ( .A(n3), .Z(n675) );
  HS65_LH_IVX9 U2992 ( .A(n2), .Z(n674) );
  HS65_LH_IVX9 U2993 ( .A(n1), .Z(n673) );
  HS65_LH_IVX9 U2994 ( .A(\regfile_i[ADRREAD1][2] ), .Z(n776) );
  HS65_LH_IVX9 U2995 ( .A(\regfile_i[ADRREAD0][2] ), .Z(n771) );
  HS65_LH_IVX9 U2996 ( .A(n128), .Z(n672) );
  HS65_LH_IVX9 U2997 ( .A(n127), .Z(n671) );
  HS65_LH_IVX9 U2998 ( .A(n126), .Z(n670) );
  HS65_LH_IVX9 U2999 ( .A(n125), .Z(n669) );
  HS65_LH_IVX9 U3000 ( .A(n124), .Z(n668) );
  HS65_LH_IVX9 U3001 ( .A(n123), .Z(n667) );
  HS65_LH_IVX9 U3002 ( .A(n122), .Z(n666) );
  HS65_LH_IVX9 U3003 ( .A(n121), .Z(n665) );
  HS65_LH_IVX9 U3004 ( .A(n120), .Z(n664) );
  HS65_LH_IVX9 U3005 ( .A(n119), .Z(n663) );
  HS65_LH_IVX9 U3006 ( .A(n118), .Z(n662) );
  HS65_LH_IVX9 U3007 ( .A(n117), .Z(n661) );
  HS65_LH_IVX9 U3008 ( .A(n116), .Z(n660) );
  HS65_LH_IVX9 U3009 ( .A(n115), .Z(n659) );
  HS65_LH_IVX9 U3010 ( .A(n114), .Z(n658) );
  HS65_LH_IVX9 U3011 ( .A(n113), .Z(n657) );
  HS65_LH_IVX9 U3012 ( .A(n112), .Z(n656) );
  HS65_LH_IVX9 U3013 ( .A(n111), .Z(n655) );
  HS65_LH_IVX9 U3014 ( .A(n110), .Z(n654) );
  HS65_LH_IVX9 U3015 ( .A(n109), .Z(n653) );
  HS65_LH_IVX9 U3016 ( .A(n108), .Z(n652) );
  HS65_LH_IVX9 U3017 ( .A(n107), .Z(n651) );
  HS65_LH_IVX9 U3018 ( .A(n106), .Z(n650) );
  HS65_LH_IVX9 U3019 ( .A(n105), .Z(n649) );
  HS65_LH_IVX9 U3020 ( .A(n104), .Z(n648) );
  HS65_LH_IVX9 U3021 ( .A(n103), .Z(n647) );
  HS65_LH_IVX9 U3022 ( .A(n102), .Z(n646) );
  HS65_LH_IVX9 U3023 ( .A(n101), .Z(n645) );
  HS65_LH_IVX9 U3024 ( .A(n100), .Z(n644) );
  HS65_LH_IVX9 U3025 ( .A(n99), .Z(n643) );
  HS65_LH_IVX9 U3026 ( .A(n98), .Z(n642) );
  HS65_LH_IVX9 U3027 ( .A(n97), .Z(n641) );
  HS65_LH_IVX9 U3028 ( .A(\regfile_i[ADRREAD1][1] ), .Z(n777) );
  HS65_LH_IVX9 U3029 ( .A(\regfile_i[ADRREAD0][1] ), .Z(n772) );
  HS65_LH_IVX9 U3030 ( .A(n256), .Z(n768) );
  HS65_LH_IVX9 U3031 ( .A(n255), .Z(n767) );
  HS65_LH_IVX9 U3032 ( .A(n254), .Z(n766) );
  HS65_LH_IVX9 U3033 ( .A(n253), .Z(n765) );
  HS65_LH_IVX9 U3034 ( .A(n252), .Z(n764) );
  HS65_LH_IVX9 U3035 ( .A(n251), .Z(n763) );
  HS65_LH_IVX9 U3036 ( .A(n250), .Z(n762) );
  HS65_LH_IVX9 U3037 ( .A(n249), .Z(n761) );
  HS65_LH_IVX9 U3038 ( .A(n248), .Z(n760) );
  HS65_LH_IVX9 U3039 ( .A(n247), .Z(n759) );
  HS65_LH_IVX9 U3040 ( .A(n246), .Z(n758) );
  HS65_LH_IVX9 U3041 ( .A(n245), .Z(n757) );
  HS65_LH_IVX9 U3042 ( .A(n244), .Z(n756) );
  HS65_LH_IVX9 U3043 ( .A(n243), .Z(n755) );
  HS65_LH_IVX9 U3044 ( .A(n242), .Z(n754) );
  HS65_LH_IVX9 U3045 ( .A(n241), .Z(n753) );
  HS65_LH_IVX9 U3046 ( .A(n240), .Z(n752) );
  HS65_LH_IVX9 U3047 ( .A(n239), .Z(n751) );
  HS65_LH_IVX9 U3048 ( .A(n238), .Z(n750) );
  HS65_LH_IVX9 U3049 ( .A(n237), .Z(n749) );
  HS65_LH_IVX9 U3050 ( .A(n236), .Z(n748) );
  HS65_LH_IVX9 U3051 ( .A(n235), .Z(n747) );
  HS65_LH_IVX9 U3052 ( .A(n234), .Z(n746) );
  HS65_LH_IVX9 U3053 ( .A(n233), .Z(n745) );
  HS65_LH_IVX9 U3054 ( .A(n232), .Z(n744) );
  HS65_LH_IVX9 U3055 ( .A(n231), .Z(n743) );
  HS65_LH_IVX9 U3056 ( .A(n230), .Z(n742) );
  HS65_LH_IVX9 U3057 ( .A(n229), .Z(n741) );
  HS65_LH_IVX9 U3058 ( .A(n228), .Z(n740) );
  HS65_LH_IVX9 U3059 ( .A(n227), .Z(n739) );
  HS65_LH_IVX9 U3060 ( .A(n226), .Z(n738) );
  HS65_LH_IVX9 U3061 ( .A(n225), .Z(n737) );
  HS65_LH_IVX9 U3062 ( .A(n64), .Z(n608) );
  HS65_LH_IVX9 U3063 ( .A(n63), .Z(n607) );
  HS65_LH_IVX9 U3064 ( .A(n62), .Z(n606) );
  HS65_LH_IVX9 U3065 ( .A(n61), .Z(n605) );
  HS65_LH_IVX9 U3066 ( .A(n60), .Z(n604) );
  HS65_LH_IVX9 U3067 ( .A(n59), .Z(n603) );
  HS65_LH_IVX9 U3068 ( .A(n58), .Z(n602) );
  HS65_LH_IVX9 U3069 ( .A(n57), .Z(n601) );
  HS65_LH_IVX9 U3070 ( .A(n56), .Z(n600) );
  HS65_LH_IVX9 U3071 ( .A(n55), .Z(n599) );
  HS65_LH_IVX9 U3072 ( .A(n54), .Z(n598) );
  HS65_LH_IVX9 U3073 ( .A(n53), .Z(n597) );
  HS65_LH_IVX9 U3074 ( .A(n52), .Z(n596) );
  HS65_LH_IVX9 U3075 ( .A(n51), .Z(n595) );
  HS65_LH_IVX9 U3076 ( .A(n50), .Z(n594) );
  HS65_LH_IVX9 U3077 ( .A(n49), .Z(n593) );
  HS65_LH_IVX9 U3078 ( .A(n48), .Z(n592) );
  HS65_LH_IVX9 U3079 ( .A(n47), .Z(n591) );
  HS65_LH_IVX9 U3080 ( .A(n46), .Z(n590) );
  HS65_LH_IVX9 U3081 ( .A(n45), .Z(n589) );
  HS65_LH_IVX9 U3082 ( .A(n44), .Z(n588) );
  HS65_LH_IVX9 U3083 ( .A(n43), .Z(n587) );
  HS65_LH_IVX9 U3084 ( .A(n42), .Z(n586) );
  HS65_LH_IVX9 U3085 ( .A(n41), .Z(n585) );
  HS65_LH_IVX9 U3086 ( .A(n40), .Z(n584) );
  HS65_LH_IVX9 U3087 ( .A(n39), .Z(n583) );
  HS65_LH_IVX9 U3088 ( .A(n38), .Z(n582) );
  HS65_LH_IVX9 U3089 ( .A(n37), .Z(n581) );
  HS65_LH_IVX9 U3090 ( .A(n36), .Z(n580) );
  HS65_LH_IVX9 U3091 ( .A(n35), .Z(n579) );
  HS65_LH_IVX9 U3092 ( .A(n34), .Z(n578) );
  HS65_LH_IVX9 U3093 ( .A(n33), .Z(n577) );
  HS65_LH_IVX9 U3094 ( .A(n192), .Z(n640) );
  HS65_LH_IVX9 U3095 ( .A(n191), .Z(n639) );
  HS65_LH_IVX9 U3096 ( .A(n190), .Z(n638) );
  HS65_LH_IVX9 U3097 ( .A(n189), .Z(n637) );
  HS65_LH_IVX9 U3098 ( .A(n188), .Z(n636) );
  HS65_LH_IVX9 U3099 ( .A(n187), .Z(n635) );
  HS65_LH_IVX9 U3100 ( .A(n186), .Z(n634) );
  HS65_LH_IVX9 U3101 ( .A(n185), .Z(n633) );
  HS65_LH_IVX9 U3102 ( .A(n184), .Z(n632) );
  HS65_LH_IVX9 U3103 ( .A(n183), .Z(n631) );
  HS65_LH_IVX9 U3104 ( .A(n182), .Z(n630) );
  HS65_LH_IVX9 U3105 ( .A(n181), .Z(n629) );
  HS65_LH_IVX9 U3106 ( .A(n180), .Z(n628) );
  HS65_LH_IVX9 U3107 ( .A(n179), .Z(n627) );
  HS65_LH_IVX9 U3108 ( .A(n178), .Z(n626) );
  HS65_LH_IVX9 U3109 ( .A(n177), .Z(n625) );
  HS65_LH_IVX9 U3110 ( .A(n176), .Z(n624) );
  HS65_LH_IVX9 U3111 ( .A(n175), .Z(n623) );
  HS65_LH_IVX9 U3112 ( .A(n174), .Z(n622) );
  HS65_LH_IVX9 U3113 ( .A(n173), .Z(n621) );
  HS65_LH_IVX9 U3114 ( .A(n172), .Z(n620) );
  HS65_LH_IVX9 U3115 ( .A(n171), .Z(n619) );
  HS65_LH_IVX9 U3116 ( .A(n170), .Z(n618) );
  HS65_LH_IVX9 U3117 ( .A(n169), .Z(n617) );
  HS65_LH_IVX9 U3118 ( .A(n168), .Z(n616) );
  HS65_LH_IVX9 U3119 ( .A(n167), .Z(n615) );
  HS65_LH_IVX9 U3120 ( .A(n166), .Z(n614) );
  HS65_LH_IVX9 U3121 ( .A(n165), .Z(n613) );
  HS65_LH_IVX9 U3122 ( .A(n164), .Z(n612) );
  HS65_LH_IVX9 U3123 ( .A(n163), .Z(n611) );
  HS65_LH_IVX9 U3124 ( .A(n162), .Z(n610) );
  HS65_LH_IVX9 U3125 ( .A(n161), .Z(n609) );
  HS65_LH_IVX9 U3126 ( .A(\regfile_i[ADRWRITE][4] ), .Z(n795) );
  HS65_LH_IVX9 U3127 ( .A(\regfile_i[ADRWRITE][3] ), .Z(n811) );
endmodule


module id_top ( clk, rst_n, .id_top_i({\id_top_i[INSTRUCTION][31] , 
        \id_top_i[INSTRUCTION][30] , \id_top_i[INSTRUCTION][29] , 
        \id_top_i[INSTRUCTION][28] , \id_top_i[INSTRUCTION][27] , 
        \id_top_i[INSTRUCTION][26] , \id_top_i[INSTRUCTION][25] , 
        \id_top_i[INSTRUCTION][24] , \id_top_i[INSTRUCTION][23] , 
        \id_top_i[INSTRUCTION][22] , \id_top_i[INSTRUCTION][21] , 
        \id_top_i[INSTRUCTION][20] , \id_top_i[INSTRUCTION][19] , 
        \id_top_i[INSTRUCTION][18] , \id_top_i[INSTRUCTION][17] , 
        \id_top_i[INSTRUCTION][16] , \id_top_i[INSTRUCTION][15] , 
        \id_top_i[INSTRUCTION][14] , \id_top_i[INSTRUCTION][13] , 
        \id_top_i[INSTRUCTION][12] , \id_top_i[INSTRUCTION][11] , 
        \id_top_i[INSTRUCTION][10] , \id_top_i[INSTRUCTION][9] , 
        \id_top_i[INSTRUCTION][8] , \id_top_i[INSTRUCTION][7] , 
        \id_top_i[INSTRUCTION][6] , \id_top_i[INSTRUCTION][5] , 
        \id_top_i[INSTRUCTION][4] , \id_top_i[INSTRUCTION][3] , 
        \id_top_i[INSTRUCTION][2] , \id_top_i[INSTRUCTION][1] , 
        \id_top_i[INSTRUCTION][0] , \id_top_i[WRITEBACK_DATA][31] , 
        \id_top_i[WRITEBACK_DATA][30] , \id_top_i[WRITEBACK_DATA][29] , 
        \id_top_i[WRITEBACK_DATA][28] , \id_top_i[WRITEBACK_DATA][27] , 
        \id_top_i[WRITEBACK_DATA][26] , \id_top_i[WRITEBACK_DATA][25] , 
        \id_top_i[WRITEBACK_DATA][24] , \id_top_i[WRITEBACK_DATA][23] , 
        \id_top_i[WRITEBACK_DATA][22] , \id_top_i[WRITEBACK_DATA][21] , 
        \id_top_i[WRITEBACK_DATA][20] , \id_top_i[WRITEBACK_DATA][19] , 
        \id_top_i[WRITEBACK_DATA][18] , \id_top_i[WRITEBACK_DATA][17] , 
        \id_top_i[WRITEBACK_DATA][16] , \id_top_i[WRITEBACK_DATA][15] , 
        \id_top_i[WRITEBACK_DATA][14] , \id_top_i[WRITEBACK_DATA][13] , 
        \id_top_i[WRITEBACK_DATA][12] , \id_top_i[WRITEBACK_DATA][11] , 
        \id_top_i[WRITEBACK_DATA][10] , \id_top_i[WRITEBACK_DATA][9] , 
        \id_top_i[WRITEBACK_DATA][8] , \id_top_i[WRITEBACK_DATA][7] , 
        \id_top_i[WRITEBACK_DATA][6] , \id_top_i[WRITEBACK_DATA][5] , 
        \id_top_i[WRITEBACK_DATA][4] , \id_top_i[WRITEBACK_DATA][3] , 
        \id_top_i[WRITEBACK_DATA][2] , \id_top_i[WRITEBACK_DATA][1] , 
        \id_top_i[WRITEBACK_DATA][0] , \id_top_i[FORWARD_A] , 
        \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] , \id_top_i[WRITE_REG][4] , 
        \id_top_i[WRITE_REG][3] , \id_top_i[WRITE_REG][2] , 
        \id_top_i[WRITE_REG][1] , \id_top_i[WRITE_REG][0] }), .id_top_o({
        \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] , 
        \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] , 
        \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] , 
        \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] , 
        \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] , 
        \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] , 
        \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] , 
        \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] , 
        \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] , 
        \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] , 
        \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] , 
        \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] , 
        \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] , 
        \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] , 
        \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] , 
        \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] , 
        \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] , 
        \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] , 
        \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] , 
        \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] , 
        \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] , 
        \id_top_o[REG_B][0] , \id_top_o[INSTR_31_26][5] , 
        \id_top_o[INSTR_31_26][4] , \id_top_o[INSTR_31_26][3] , 
        \id_top_o[INSTR_31_26][2] , \id_top_o[INSTR_31_26][1] , 
        \id_top_o[INSTR_31_26][0] , \id_top_o[RS][4] , \id_top_o[RS][3] , 
        \id_top_o[RS][2] , \id_top_o[RS][1] , \id_top_o[RS][0] , 
        \id_top_o[RT][4] , \id_top_o[RT][3] , \id_top_o[RT][2] , 
        \id_top_o[RT][1] , \id_top_o[RT][0] , \id_top_o[RD][4] , 
        \id_top_o[RD][3] , \id_top_o[RD][2] , \id_top_o[RD][1] , 
        \id_top_o[RD][0] , \id_top_o[INSTR_10_6][4] , 
        \id_top_o[INSTR_10_6][3] , \id_top_o[INSTR_10_6][2] , 
        \id_top_o[INSTR_10_6][1] , \id_top_o[INSTR_10_6][0] , 
        \id_top_o[INSTR_5_0][5] , \id_top_o[INSTR_5_0][4] , 
        \id_top_o[INSTR_5_0][3] , \id_top_o[INSTR_5_0][2] , 
        \id_top_o[INSTR_5_0][1] , \id_top_o[INSTR_5_0][0] , 
        \id_top_o[SIGN_EXTEND][31] , \id_top_o[SIGN_EXTEND][30] , 
        \id_top_o[SIGN_EXTEND][29] , \id_top_o[SIGN_EXTEND][28] , 
        \id_top_o[SIGN_EXTEND][27] , \id_top_o[SIGN_EXTEND][26] , 
        \id_top_o[SIGN_EXTEND][25] , \id_top_o[SIGN_EXTEND][24] , 
        \id_top_o[SIGN_EXTEND][23] , \id_top_o[SIGN_EXTEND][22] , 
        \id_top_o[SIGN_EXTEND][21] , \id_top_o[SIGN_EXTEND][20] , 
        \id_top_o[SIGN_EXTEND][19] , \id_top_o[SIGN_EXTEND][18] , 
        \id_top_o[SIGN_EXTEND][17] , \id_top_o[SIGN_EXTEND][16] , 
        \id_top_o[SIGN_EXTEND][15] , \id_top_o[SIGN_EXTEND][14] , 
        \id_top_o[SIGN_EXTEND][13] , \id_top_o[SIGN_EXTEND][12] , 
        \id_top_o[SIGN_EXTEND][11] , \id_top_o[SIGN_EXTEND][10] , 
        \id_top_o[SIGN_EXTEND][9] , \id_top_o[SIGN_EXTEND][8] , 
        \id_top_o[SIGN_EXTEND][7] , \id_top_o[SIGN_EXTEND][6] , 
        \id_top_o[SIGN_EXTEND][5] , \id_top_o[SIGN_EXTEND][4] , 
        \id_top_o[SIGN_EXTEND][3] , \id_top_o[SIGN_EXTEND][2] , 
        \id_top_o[SIGN_EXTEND][1] , \id_top_o[SIGN_EXTEND][0] }) );
  input clk, rst_n, \id_top_i[INSTRUCTION][31] , \id_top_i[INSTRUCTION][30] ,
         \id_top_i[INSTRUCTION][29] , \id_top_i[INSTRUCTION][28] ,
         \id_top_i[INSTRUCTION][27] , \id_top_i[INSTRUCTION][26] ,
         \id_top_i[INSTRUCTION][25] , \id_top_i[INSTRUCTION][24] ,
         \id_top_i[INSTRUCTION][23] , \id_top_i[INSTRUCTION][22] ,
         \id_top_i[INSTRUCTION][21] , \id_top_i[INSTRUCTION][20] ,
         \id_top_i[INSTRUCTION][19] , \id_top_i[INSTRUCTION][18] ,
         \id_top_i[INSTRUCTION][17] , \id_top_i[INSTRUCTION][16] ,
         \id_top_i[INSTRUCTION][15] , \id_top_i[INSTRUCTION][14] ,
         \id_top_i[INSTRUCTION][13] , \id_top_i[INSTRUCTION][12] ,
         \id_top_i[INSTRUCTION][11] , \id_top_i[INSTRUCTION][10] ,
         \id_top_i[INSTRUCTION][9] , \id_top_i[INSTRUCTION][8] ,
         \id_top_i[INSTRUCTION][7] , \id_top_i[INSTRUCTION][6] ,
         \id_top_i[INSTRUCTION][5] , \id_top_i[INSTRUCTION][4] ,
         \id_top_i[INSTRUCTION][3] , \id_top_i[INSTRUCTION][2] ,
         \id_top_i[INSTRUCTION][1] , \id_top_i[INSTRUCTION][0] ,
         \id_top_i[WRITEBACK_DATA][31] , \id_top_i[WRITEBACK_DATA][30] ,
         \id_top_i[WRITEBACK_DATA][29] , \id_top_i[WRITEBACK_DATA][28] ,
         \id_top_i[WRITEBACK_DATA][27] , \id_top_i[WRITEBACK_DATA][26] ,
         \id_top_i[WRITEBACK_DATA][25] , \id_top_i[WRITEBACK_DATA][24] ,
         \id_top_i[WRITEBACK_DATA][23] , \id_top_i[WRITEBACK_DATA][22] ,
         \id_top_i[WRITEBACK_DATA][21] , \id_top_i[WRITEBACK_DATA][20] ,
         \id_top_i[WRITEBACK_DATA][19] , \id_top_i[WRITEBACK_DATA][18] ,
         \id_top_i[WRITEBACK_DATA][17] , \id_top_i[WRITEBACK_DATA][16] ,
         \id_top_i[WRITEBACK_DATA][15] , \id_top_i[WRITEBACK_DATA][14] ,
         \id_top_i[WRITEBACK_DATA][13] , \id_top_i[WRITEBACK_DATA][12] ,
         \id_top_i[WRITEBACK_DATA][11] , \id_top_i[WRITEBACK_DATA][10] ,
         \id_top_i[WRITEBACK_DATA][9] , \id_top_i[WRITEBACK_DATA][8] ,
         \id_top_i[WRITEBACK_DATA][7] , \id_top_i[WRITEBACK_DATA][6] ,
         \id_top_i[WRITEBACK_DATA][5] , \id_top_i[WRITEBACK_DATA][4] ,
         \id_top_i[WRITEBACK_DATA][3] , \id_top_i[WRITEBACK_DATA][2] ,
         \id_top_i[WRITEBACK_DATA][1] , \id_top_i[WRITEBACK_DATA][0] ,
         \id_top_i[FORWARD_A] , \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] ,
         \id_top_i[WRITE_REG][4] , \id_top_i[WRITE_REG][3] ,
         \id_top_i[WRITE_REG][2] , \id_top_i[WRITE_REG][1] ,
         \id_top_i[WRITE_REG][0] ;
  output \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] ,
         \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] ,
         \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] ,
         \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] ,
         \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] ,
         \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] ,
         \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] ,
         \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] ,
         \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] ,
         \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] ,
         \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] ,
         \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] ,
         \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] ,
         \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] ,
         \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] ,
         \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] ,
         \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] ,
         \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] ,
         \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] ,
         \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] ,
         \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] ,
         \id_top_o[REG_B][0] , \id_top_o[INSTR_31_26][5] ,
         \id_top_o[INSTR_31_26][4] , \id_top_o[INSTR_31_26][3] ,
         \id_top_o[INSTR_31_26][2] , \id_top_o[INSTR_31_26][1] ,
         \id_top_o[INSTR_31_26][0] , \id_top_o[RS][4] , \id_top_o[RS][3] ,
         \id_top_o[RS][2] , \id_top_o[RS][1] , \id_top_o[RS][0] ,
         \id_top_o[RT][4] , \id_top_o[RT][3] , \id_top_o[RT][2] ,
         \id_top_o[RT][1] , \id_top_o[RT][0] , \id_top_o[RD][4] ,
         \id_top_o[RD][3] , \id_top_o[RD][2] , \id_top_o[RD][1] ,
         \id_top_o[RD][0] , \id_top_o[INSTR_10_6][4] ,
         \id_top_o[INSTR_10_6][3] , \id_top_o[INSTR_10_6][2] ,
         \id_top_o[INSTR_10_6][1] , \id_top_o[INSTR_10_6][0] ,
         \id_top_o[INSTR_5_0][5] , \id_top_o[INSTR_5_0][4] ,
         \id_top_o[INSTR_5_0][3] , \id_top_o[INSTR_5_0][2] ,
         \id_top_o[INSTR_5_0][1] , \id_top_o[INSTR_5_0][0] ,
         \id_top_o[SIGN_EXTEND][31] , \id_top_o[SIGN_EXTEND][30] ,
         \id_top_o[SIGN_EXTEND][29] , \id_top_o[SIGN_EXTEND][28] ,
         \id_top_o[SIGN_EXTEND][27] , \id_top_o[SIGN_EXTEND][26] ,
         \id_top_o[SIGN_EXTEND][25] , \id_top_o[SIGN_EXTEND][24] ,
         \id_top_o[SIGN_EXTEND][23] , \id_top_o[SIGN_EXTEND][22] ,
         \id_top_o[SIGN_EXTEND][21] , \id_top_o[SIGN_EXTEND][20] ,
         \id_top_o[SIGN_EXTEND][19] , \id_top_o[SIGN_EXTEND][18] ,
         \id_top_o[SIGN_EXTEND][17] , \id_top_o[SIGN_EXTEND][16] ,
         \id_top_o[SIGN_EXTEND][15] , \id_top_o[SIGN_EXTEND][14] ,
         \id_top_o[SIGN_EXTEND][13] , \id_top_o[SIGN_EXTEND][12] ,
         \id_top_o[SIGN_EXTEND][11] , \id_top_o[SIGN_EXTEND][10] ,
         \id_top_o[SIGN_EXTEND][9] , \id_top_o[SIGN_EXTEND][8] ,
         \id_top_o[SIGN_EXTEND][7] , \id_top_o[SIGN_EXTEND][6] ,
         \id_top_o[SIGN_EXTEND][5] , \id_top_o[SIGN_EXTEND][4] ,
         \id_top_o[SIGN_EXTEND][3] , \id_top_o[SIGN_EXTEND][2] ,
         \id_top_o[SIGN_EXTEND][1] , \id_top_o[SIGN_EXTEND][0] ;
  wire   \id_top_o[INSTR_31_26][5] , \id_top_o[INSTR_31_26][4] ,
         \id_top_o[INSTR_31_26][3] , \id_top_o[INSTR_31_26][2] ,
         \id_top_o[INSTR_31_26][1] , \id_top_o[INSTR_31_26][0] ,
         \id_top_o[RS][4] , \id_top_o[RS][3] , \id_top_o[RS][2] ,
         \id_top_o[RS][1] , \id_top_o[RS][0] , \id_top_o[RT][4] ,
         \id_top_o[RT][3] , \id_top_o[RT][2] , \id_top_o[RT][1] ,
         \id_top_o[RT][0] , \id_top_o[RD][4] , \id_top_o[RD][3] ,
         \id_top_o[RD][2] , \id_top_o[RD][1] , \id_top_o[RD][0] ,
         \id_top_o[INSTR_10_6][4] , \id_top_o[INSTR_10_6][3] ,
         \id_top_o[INSTR_10_6][2] , \id_top_o[INSTR_10_6][1] ,
         \id_top_o[INSTR_10_6][0] , \id_top_o[INSTR_5_0][5] ,
         \id_top_o[INSTR_5_0][4] , \id_top_o[INSTR_5_0][3] ,
         \id_top_o[INSTR_5_0][2] , \id_top_o[INSTR_5_0][1] ,
         \id_top_o[INSTR_5_0][0] ;
  assign \id_top_o[INSTR_31_26][5]  = \id_top_i[INSTRUCTION][31] ;
  assign \id_top_o[INSTR_31_26][4]  = \id_top_i[INSTRUCTION][30] ;
  assign \id_top_o[INSTR_31_26][3]  = \id_top_i[INSTRUCTION][29] ;
  assign \id_top_o[INSTR_31_26][2]  = \id_top_i[INSTRUCTION][28] ;
  assign \id_top_o[INSTR_31_26][1]  = \id_top_i[INSTRUCTION][27] ;
  assign \id_top_o[INSTR_31_26][0]  = \id_top_i[INSTRUCTION][26] ;
  assign \id_top_o[RS][4]  = \id_top_i[INSTRUCTION][25] ;
  assign \id_top_o[RS][3]  = \id_top_i[INSTRUCTION][24] ;
  assign \id_top_o[RS][2]  = \id_top_i[INSTRUCTION][23] ;
  assign \id_top_o[RS][1]  = \id_top_i[INSTRUCTION][22] ;
  assign \id_top_o[RS][0]  = \id_top_i[INSTRUCTION][21] ;
  assign \id_top_o[RT][4]  = \id_top_i[INSTRUCTION][20] ;
  assign \id_top_o[RT][3]  = \id_top_i[INSTRUCTION][19] ;
  assign \id_top_o[RT][2]  = \id_top_i[INSTRUCTION][18] ;
  assign \id_top_o[RT][1]  = \id_top_i[INSTRUCTION][17] ;
  assign \id_top_o[RT][0]  = \id_top_i[INSTRUCTION][16] ;
  assign \id_top_o[SIGN_EXTEND][15]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][16]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][17]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][18]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][19]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][20]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][21]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][22]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][23]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][24]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][25]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][26]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][27]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][28]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][29]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][30]  = \id_top_o[RD][4] ;
  assign \id_top_o[SIGN_EXTEND][31]  = \id_top_o[RD][4] ;
  assign \id_top_o[RD][4]  = \id_top_i[INSTRUCTION][15] ;
  assign \id_top_o[SIGN_EXTEND][14]  = \id_top_o[RD][3] ;
  assign \id_top_o[RD][3]  = \id_top_i[INSTRUCTION][14] ;
  assign \id_top_o[SIGN_EXTEND][13]  = \id_top_o[RD][2] ;
  assign \id_top_o[RD][2]  = \id_top_i[INSTRUCTION][13] ;
  assign \id_top_o[SIGN_EXTEND][12]  = \id_top_o[RD][1] ;
  assign \id_top_o[RD][1]  = \id_top_i[INSTRUCTION][12] ;
  assign \id_top_o[SIGN_EXTEND][11]  = \id_top_o[RD][0] ;
  assign \id_top_o[RD][0]  = \id_top_i[INSTRUCTION][11] ;
  assign \id_top_o[SIGN_EXTEND][10]  = \id_top_o[INSTR_10_6][4] ;
  assign \id_top_o[INSTR_10_6][4]  = \id_top_i[INSTRUCTION][10] ;
  assign \id_top_o[SIGN_EXTEND][9]  = \id_top_o[INSTR_10_6][3] ;
  assign \id_top_o[INSTR_10_6][3]  = \id_top_i[INSTRUCTION][9] ;
  assign \id_top_o[SIGN_EXTEND][8]  = \id_top_o[INSTR_10_6][2] ;
  assign \id_top_o[INSTR_10_6][2]  = \id_top_i[INSTRUCTION][8] ;
  assign \id_top_o[SIGN_EXTEND][7]  = \id_top_o[INSTR_10_6][1] ;
  assign \id_top_o[INSTR_10_6][1]  = \id_top_i[INSTRUCTION][7] ;
  assign \id_top_o[SIGN_EXTEND][6]  = \id_top_o[INSTR_10_6][0] ;
  assign \id_top_o[INSTR_10_6][0]  = \id_top_i[INSTRUCTION][6] ;
  assign \id_top_o[SIGN_EXTEND][5]  = \id_top_o[INSTR_5_0][5] ;
  assign \id_top_o[INSTR_5_0][5]  = \id_top_i[INSTRUCTION][5] ;
  assign \id_top_o[SIGN_EXTEND][4]  = \id_top_o[INSTR_5_0][4] ;
  assign \id_top_o[INSTR_5_0][4]  = \id_top_i[INSTRUCTION][4] ;
  assign \id_top_o[SIGN_EXTEND][3]  = \id_top_o[INSTR_5_0][3] ;
  assign \id_top_o[INSTR_5_0][3]  = \id_top_i[INSTRUCTION][3] ;
  assign \id_top_o[SIGN_EXTEND][2]  = \id_top_o[INSTR_5_0][2] ;
  assign \id_top_o[INSTR_5_0][2]  = \id_top_i[INSTRUCTION][2] ;
  assign \id_top_o[SIGN_EXTEND][1]  = \id_top_o[INSTR_5_0][1] ;
  assign \id_top_o[INSTR_5_0][1]  = \id_top_i[INSTRUCTION][1] ;
  assign \id_top_o[SIGN_EXTEND][0]  = \id_top_o[INSTR_5_0][0] ;
  assign \id_top_o[INSTR_5_0][0]  = \id_top_i[INSTRUCTION][0] ;

  regfile regfile_inst ( .clk(clk), .rst_n(rst_n), .regfile_i({
        \id_top_o[RS][4] , \id_top_o[RS][3] , \id_top_o[RS][2] , 
        \id_top_o[RS][1] , \id_top_o[RS][0] , \id_top_o[RT][4] , 
        \id_top_o[RT][3] , \id_top_o[RT][2] , \id_top_o[RT][1] , 
        \id_top_o[RT][0] , \id_top_i[WRITE_REG][4] , \id_top_i[WRITE_REG][3] , 
        \id_top_i[WRITE_REG][2] , \id_top_i[WRITE_REG][1] , 
        \id_top_i[WRITE_REG][0] , \id_top_i[WRITEBACK_DATA][31] , 
        \id_top_i[WRITEBACK_DATA][30] , \id_top_i[WRITEBACK_DATA][29] , 
        \id_top_i[WRITEBACK_DATA][28] , \id_top_i[WRITEBACK_DATA][27] , 
        \id_top_i[WRITEBACK_DATA][26] , \id_top_i[WRITEBACK_DATA][25] , 
        \id_top_i[WRITEBACK_DATA][24] , \id_top_i[WRITEBACK_DATA][23] , 
        \id_top_i[WRITEBACK_DATA][22] , \id_top_i[WRITEBACK_DATA][21] , 
        \id_top_i[WRITEBACK_DATA][20] , \id_top_i[WRITEBACK_DATA][19] , 
        \id_top_i[WRITEBACK_DATA][18] , \id_top_i[WRITEBACK_DATA][17] , 
        \id_top_i[WRITEBACK_DATA][16] , \id_top_i[WRITEBACK_DATA][15] , 
        \id_top_i[WRITEBACK_DATA][14] , \id_top_i[WRITEBACK_DATA][13] , 
        \id_top_i[WRITEBACK_DATA][12] , \id_top_i[WRITEBACK_DATA][11] , 
        \id_top_i[WRITEBACK_DATA][10] , \id_top_i[WRITEBACK_DATA][9] , 
        \id_top_i[WRITEBACK_DATA][8] , \id_top_i[WRITEBACK_DATA][7] , 
        \id_top_i[WRITEBACK_DATA][6] , \id_top_i[WRITEBACK_DATA][5] , 
        \id_top_i[WRITEBACK_DATA][4] , \id_top_i[WRITEBACK_DATA][3] , 
        \id_top_i[WRITEBACK_DATA][2] , \id_top_i[WRITEBACK_DATA][1] , 
        \id_top_i[WRITEBACK_DATA][0] , \id_top_i[FORWARD_A] , 
        \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] }), .regfile_o({
        \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] , 
        \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] , 
        \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] , 
        \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] , 
        \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] , 
        \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] , 
        \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] , 
        \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] , 
        \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] , 
        \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] , 
        \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] , 
        \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] , 
        \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] , 
        \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] , 
        \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] , 
        \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] , 
        \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] , 
        \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] , 
        \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] , 
        \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] , 
        \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] , 
        \id_top_o[REG_B][0] }) );
endmodule

