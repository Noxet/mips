
library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity exe_top_DW01_add_0 is

   port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (11 downto 0);  CO : out std_logic);

end exe_top_DW01_add_0;

architecture SYN_rpl of exe_top_DW01_add_0 is

   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1 : std_logic;

begin
   
   U1_11 : HS65_LHS_XOR3X2 port map( A => A(11), B => B(11), C => carry_11_port
                           , Z => SUM(11));
   U1_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => B(10), CI => 
                           carry_10_port, CO => carry_11_port, S0 => SUM(10));
   U1_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => B(9), CI => carry_9_port, 
                           CO => carry_10_port, S0 => SUM(9));
   U1_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => B(8), CI => carry_8_port, 
                           CO => carry_9_port, S0 => SUM(8));
   U1_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => B(7), CI => carry_7_port, 
                           CO => carry_8_port, S0 => SUM(7));
   U1_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => B(6), CI => carry_6_port, 
                           CO => carry_7_port, S0 => SUM(6));
   U1_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => B(5), CI => carry_5_port, 
                           CO => carry_6_port, S0 => SUM(5));
   U1_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => B(4), CI => carry_4_port, 
                           CO => carry_5_port, S0 => SUM(4));
   U1_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => B(3), CI => carry_3_port, 
                           CO => carry_4_port, S0 => SUM(3));
   U1_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => B(2), CI => carry_2_port, 
                           CO => carry_3_port, S0 => SUM(2));
   U1_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => B(1), CI => n1, CO => 
                           carry_2_port, S0 => SUM(1));
   U1 : HS65_LH_AND2X4 port map( A => A(0), B => B(0), Z => n1);
   U2 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => SUM(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_mult_uns_0 is

   port( a, b : in std_logic_vector (31 downto 0);  product : out 
         std_logic_vector (63 downto 0));

end alu_DW_mult_uns_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_mult_uns_0 is

   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_HA1X4
      port( A0, B0 : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n292, n293, n294, n295, n296, n297, n299, n300, 
      n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n330, n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n354, 
      n355, n356, n357, n358, n359, n360, n361, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n2417, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, 
      n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
      n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
      n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, 
      n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
      n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
      n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, 
      n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
      n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
      n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, 
      n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, 
      n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, 
      n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
      n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
      n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, 
      n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, 
      n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, 
      n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, 
      n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, 
      n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, 
      n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, 
      n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
      n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
      n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
      n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
      n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, 
      n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, 
      n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, 
      n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, 
      n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
      n3098, n3099, n3100, n3101, n3102, n3103, n3104, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719 : std_logic;

begin
   
   U1941 : HS65_LH_NOR3AX2 port map( A => n2758, B => n2754, C => n2753, Z => 
                           n2723);
   U1942 : HS65_LH_NOR3AX2 port map( A => n3058, B => n3054, C => n3053, Z => 
                           n3023);
   U1943 : HS65_LH_NOR3AX2 port map( A => n3101, B => n3097, C => n3096, Z => 
                           n3066);
   U1944 : HS65_LH_NOR3AX2 port map( A => n2929, B => n2925, C => n2924, Z => 
                           n2894);
   U1945 : HS65_LH_NOR3AX2 port map( A => n2801, B => n2797, C => n2796, Z => 
                           n2766);
   U1946 : HS65_LH_NOR3AX2 port map( A => n2843, B => n2839, C => n2838, Z => 
                           n2808);
   U1947 : HS65_LH_NOR3AX2 port map( A => n2886, B => n2882, C => n2881, Z => 
                           n2851);
   U1948 : HS65_LH_NOR3AX2 port map( A => n2972, B => n2968, C => n2967, Z => 
                           n2937);
   U1949 : HS65_LH_NOR3AX2 port map( A => n3015, B => n3011, C => n3010, Z => 
                           n2980);
   U1950 : HS65_LH_AND2X4 port map( A => n2753, B => n2754, Z => n2718);
   U1951 : HS65_LH_AND2X4 port map( A => n3010, B => n3011, Z => n2975);
   U1952 : HS65_LH_AND2X4 port map( A => n2796, B => n2797, Z => n2761);
   U1953 : HS65_LH_AND2X4 port map( A => n2838, B => n2839, Z => n2417);
   U1954 : HS65_LH_AND2X4 port map( A => n2881, B => n2882, Z => n2846);
   U1955 : HS65_LH_AND2X4 port map( A => n2924, B => n2925, Z => n2889);
   U1956 : HS65_LH_AND2X4 port map( A => n2967, B => n2968, Z => n2932);
   U1957 : HS65_LH_AND2X4 port map( A => n3053, B => n3054, Z => n3018);
   U1958 : HS65_LH_AND2X4 port map( A => n3096, B => n3097, Z => n3061);
   U1959 : HS65_LH_NOR3AX2 port map( A => a(31), B => n3104, C => n3103, Z => 
                           n2670);
   U1960 : HS65_LH_NOR3AX2 port map( A => n2711, B => a(0), C => a(1), Z => 
                           n2681);
   U1961 : HS65_LH_IVX9 port map( A => n1007, Z => n4719);
   U1962 : HS65_LH_FA1X4 port map( A0 => n530, B0 => n546, CI => n253, CO => 
                           n252, S0 => product(37));
   U1963 : HS65_LH_FA1X4 port map( A0 => n480, B0 => n494, CI => n250, CO => 
                           n249, S0 => product(40));
   U1964 : HS65_LH_FA1X4 port map( A0 => n435, B0 => n448, CI => n247, CO => 
                           n246, S0 => product(43));
   U1965 : HS65_LH_FA1X4 port map( A0 => n397, B0 => n407, CI => n244, CO => 
                           n243, S0 => product(46));
   U1966 : HS65_LH_FA1X4 port map( A0 => n364, B0 => n373, CI => n241, CO => 
                           n240, S0 => product(49));
   U1967 : HS65_LH_FA1X4 port map( A0 => n338, B0 => n344, CI => n238, CO => 
                           n237, S0 => product(52));
   U1968 : HS65_LH_FA1X4 port map( A0 => n317, B0 => n322, CI => n235, CO => 
                           n234, S0 => product(55));
   U1969 : HS65_LH_FA1X4 port map( A0 => n303, B0 => n305, CI => n232, CO => 
                           n231, S0 => product(58));
   U1970 : HS65_LH_HA1X4 port map( A0 => n4678, B0 => n975, CO => n1006, S0 => 
                           n1007);
   U1971 : HS65_LH_OAI22X6 port map( A => n4676, B => n2757, C => n4580, D => 
                           n2757, Z => n2756);
   U1972 : HS65_LH_AND2X4 port map( A => n4585, B => n4679, Z => n2757);
   U1973 : HS65_LH_OAI22X6 port map( A => n4676, B => n3100, C => n4495, D => 
                           n3100, Z => n3099);
   U1974 : HS65_LH_AND2X4 port map( A => n4500, B => n4679, Z => n3100);
   U1975 : HS65_LH_FA1X4 port map( A0 => n1351, B0 => n1319, CI => n549, CO => 
                           n546, S0 => n547);
   U1976 : HS65_LHS_XOR2X6 port map( A => n4684, B => n2759, Z => n1351);
   U1977 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2794, Z => n1319);
   U1978 : HS65_LH_AOI22X6 port map( A => n4586, B => n1006, C => n4580, D => 
                           n4678, Z => n2759);
   U1979 : HS65_LH_FA1X4 port map( A0 => n1281, B0 => n1249, CI => n451, CO => 
                           n448, S0 => n449);
   U1980 : HS65_LHS_XOR2X6 port map( A => n4690, B => n2844, Z => n1281);
   U1981 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2879, Z => n1249);
   U1982 : HS65_LH_AOI22X6 port map( A => n4567, B => n1006, C => n4561, D => 
                           n4678, Z => n2844);
   U1983 : HS65_LH_FA1X4 port map( A0 => n1141, B0 => n1109, CI => n325, CO => 
                           n322, S0 => n323);
   U1984 : HS65_LHS_XOR2X6 port map( A => n4702, B => n3016, Z => n1141);
   U1985 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3051, Z => n1109);
   U1986 : HS65_LH_AOI22X6 port map( A => n4523, B => n1006, C => n4517, D => 
                           n4678, Z => n3016);
   U1987 : HS65_LH_FA1X4 port map( A0 => n1106, B0 => n1074, CI => n308, CO => 
                           n305, S0 => n306);
   U1988 : HS65_LHS_XOR2X6 port map( A => n4705, B => n3059, Z => n1106);
   U1989 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3094, Z => n1074);
   U1990 : HS65_LH_AOI22X6 port map( A => n4512, B => n1006, C => n4506, D => 
                           n4678, Z => n3059);
   U1991 : HS65_LH_FA1X4 port map( A0 => n1318, B0 => n532, CI => n548, CO => 
                           n529, S0 => n530);
   U1992 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2795, Z => n1318);
   U1993 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1008, D1 => n4570, S1 
                           => n4675, D2 => n4574, S2 => n4677, D3 => n4579, S3 
                           => n4678, Z => n2795);
   U1994 : HS65_LH_FA1X4 port map( A0 => n1316, B0 => n1284, CI => n497, CO => 
                           n494, S0 => n495);
   U1995 : HS65_LHS_XOR2X6 port map( A => n4687, B => n2802, Z => n1316);
   U1996 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2836, Z => n1284);
   U1997 : HS65_LH_AOI22X6 port map( A => n4575, B => n1006, C => n4569, D => 
                           n4678, Z => n2802);
   U1998 : HS65_LH_FA1X4 port map( A0 => n1283, B0 => n482, CI => n496, CO => 
                           n479, S0 => n480);
   U1999 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2837, Z => n1283);
   U2000 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1008, D1 => n4566, S1 
                           => n4677, D2 => n4611, S2 => n4679, D3 => n4562, S3 
                           => n4674, Z => n2837);
   U2001 : HS65_LH_FA1X4 port map( A0 => n1248, B0 => n437, CI => n450, CO => 
                           n434, S0 => n435);
   U2002 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2880, Z => n1248);
   U2003 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1008, D1 => n4551, S1 
                           => n4675, D2 => n4555, S2 => n4677, D3 => n4560, S3 
                           => n4678, Z => n2880);
   U2004 : HS65_LH_FA1X4 port map( A0 => n1246, B0 => n1214, CI => n410, CO => 
                           n407, S0 => n408);
   U2005 : HS65_LHS_XOR2X6 port map( A => n4693, B => n2887, Z => n1246);
   U2006 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2922, Z => n1214);
   U2007 : HS65_LH_AOI22X6 port map( A => n4556, B => n1006, C => n4550, D => 
                           n4678, Z => n2887);
   U2008 : HS65_LH_FA1X4 port map( A0 => n1213, B0 => n399, CI => n409, CO => 
                           n396, S0 => n397);
   U2009 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2923, Z => n1213);
   U2010 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1008, D1 => n4540, S1 
                           => n4675, D2 => n4544, S2 => n4677, D3 => n4549, S3 
                           => n4678, Z => n2923);
   U2011 : HS65_LH_FA1X4 port map( A0 => n1211, B0 => n1179, CI => n376, CO => 
                           n373, S0 => n374);
   U2012 : HS65_LHS_XOR2X6 port map( A => n4696, B => n2930, Z => n1211);
   U2013 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2965, Z => n1179);
   U2014 : HS65_LH_AOI22X6 port map( A => n4545, B => n1006, C => n4539, D => 
                           n4678, Z => n2930);
   U2015 : HS65_LH_FA1X4 port map( A0 => n1178, B0 => n366, CI => n375, CO => 
                           n363, S0 => n364);
   U2016 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2966, Z => n1178);
   U2017 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1008, D1 => n4529, S1 
                           => n4675, D2 => n4533, S2 => n4677, D3 => n4538, S3 
                           => n4678, Z => n2966);
   U2018 : HS65_LH_FA1X4 port map( A0 => n1176, B0 => n1144, CI => n347, CO => 
                           n344, S0 => n345);
   U2019 : HS65_LHS_XOR2X6 port map( A => n4699, B => n2973, Z => n1176);
   U2020 : HS65_LHS_XOR2X6 port map( A => n4701, B => n3008, Z => n1144);
   U2021 : HS65_LH_AOI22X6 port map( A => n4534, B => n1006, C => n4528, D => 
                           n4678, Z => n2973);
   U2022 : HS65_LH_FA1X4 port map( A0 => n1143, B0 => n340, CI => n346, CO => 
                           n337, S0 => n338);
   U2023 : HS65_LHS_XOR2X6 port map( A => a(23), B => n3009, Z => n1143);
   U2024 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1008, D1 => n4527, S1 
                           => n4679, D2 => n4518, S2 => n4675, D3 => n4522, S3 
                           => n4677, Z => n3009);
   U2025 : HS65_LH_FA1X4 port map( A0 => n1108, B0 => n319, CI => n324, CO => 
                           n316, S0 => n317);
   U2026 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3052, Z => n1108);
   U2027 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1008, D1 => n4507, S1 
                           => n4674, D2 => n4511, S2 => n4677, D3 => n4516, S3 
                           => n4679, Z => n3052);
   U2028 : HS65_LH_FA1X4 port map( A0 => n1073, B0 => n304, CI => n307, CO => 
                           n302, S0 => n303);
   U2029 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3095, Z => n1073);
   U2030 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1008, D1 => n4495, S1 
                           => n4674, D2 => n4500, S2 => n4677, D3 => n4505, S3 
                           => n4679, Z => n3095);
   U2031 : HS65_LH_FA1X4 port map( A0 => n585, B0 => n602, CI => n1353, CO => 
                           n582, S0 => n583);
   U2032 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2752, Z => n1353);
   U2033 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1008, D1 => n4581, S1 
                           => n4675, D2 => n4585, S2 => n4677, D3 => n4590, S3 
                           => n4678, Z => n2752);
   U2034 : HS65_LH_HA1X4 port map( A0 => a(8), B0 => n1349, CO => n934, S0 => 
                           n935);
   U2035 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2760, Z => n1349);
   U2036 : HS65_LH_AO22X9 port map( A => n4616, B => n4579, C => n4615, D => 
                           n2762, Z => n2760);
   U2037 : HS65_LH_HA1X4 port map( A0 => a(5), B0 => n1384, CO => n940, S0 => 
                           n941);
   U2038 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2717, Z => n1384);
   U2039 : HS65_LH_AO22X9 port map( A => n4616, B => n4590, C => n4615, D => 
                           n2719, Z => n2717);
   U2040 : HS65_LH_HA1X4 port map( A0 => a(11), B0 => n1314, CO => n922, S0 => 
                           n923);
   U2041 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2803, Z => n1314);
   U2042 : HS65_LH_AO22X9 port map( A => n4616, B => n4613, C => n4615, D => 
                           n2804, Z => n2803);
   U2043 : HS65_LH_HA1X4 port map( A0 => a(14), B0 => n1279, CO => n904, S0 => 
                           n905);
   U2044 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2845, Z => n1279);
   U2045 : HS65_LH_AO22X9 port map( A => n4615, B => n4560, C => n4615, D => 
                           n2847, Z => n2845);
   U2046 : HS65_LH_HA1X4 port map( A0 => a(17), B0 => n1244, CO => n880, S0 => 
                           n881);
   U2047 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2888, Z => n1244);
   U2048 : HS65_LH_AO22X9 port map( A => n4616, B => n4549, C => n4615, D => 
                           n2890, Z => n2888);
   U2049 : HS65_LH_HA1X4 port map( A0 => a(20), B0 => n1209, CO => n850, S0 => 
                           n851);
   U2050 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2931, Z => n1209);
   U2051 : HS65_LH_AO22X9 port map( A => n4616, B => n4538, C => n4615, D => 
                           n2933, Z => n2931);
   U2052 : HS65_LH_HA1X4 port map( A0 => n4700, B0 => n1174, CO => n814, S0 => 
                           n815);
   U2053 : HS65_LHS_XOR2X6 port map( A => a(23), B => n2974, Z => n1174);
   U2054 : HS65_LH_AO22X9 port map( A => n4616, B => n4527, C => n4615, D => 
                           n2976, Z => n2974);
   U2055 : HS65_LH_HA1X4 port map( A0 => n4703, B0 => n1139, CO => n772, S0 => 
                           n773);
   U2056 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3017, Z => n1139);
   U2057 : HS65_LH_AO22X9 port map( A => n4616, B => n4516, C => n4615, D => 
                           n3019, Z => n3017);
   U2058 : HS65_LH_HA1X4 port map( A0 => a(29), B0 => n1104, CO => n724, S0 => 
                           n725);
   U2059 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3060, Z => n1104);
   U2060 : HS65_LH_AO22X9 port map( A => n4616, B => n4505, C => n4615, D => 
                           n3062, Z => n3060);
   U2061 : HS65_LH_HA1X4 port map( A0 => n1383, B0 => n940, CO => n938, S0 => 
                           n939);
   U2062 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2720, Z => n1383);
   U2063 : HS65_LH_AO222X4 port map( A => n4619, B => n4590, C => n4615, D => 
                           n4585, E => n1038, F => n2719, Z => n2720);
   U2064 : HS65_LH_HA1X4 port map( A0 => n1348, B0 => n934, CO => n930, S0 => 
                           n931);
   U2065 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2763, Z => n1348);
   U2066 : HS65_LH_AO222X4 port map( A => n4619, B => n4579, C => n4615, D => 
                           n4574, E => n1038, F => n2762, Z => n2763);
   U2067 : HS65_LH_HA1X4 port map( A0 => n1313, B0 => n922, CO => n916, S0 => 
                           n917);
   U2068 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2805, Z => n1313);
   U2069 : HS65_LH_AO222X4 port map( A => n4619, B => n4613, C => n4615, D => 
                           n4566, E => n1038, F => n2804, Z => n2805);
   U2070 : HS65_LH_HA1X4 port map( A0 => n1278, B0 => n904, CO => n896, S0 => 
                           n897);
   U2071 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2848, Z => n1278);
   U2072 : HS65_LH_AO222X4 port map( A => n4619, B => n4560, C => n4615, D => 
                           n4555, E => n1038, F => n2847, Z => n2848);
   U2073 : HS65_LH_HA1X4 port map( A0 => n1243, B0 => n880, CO => n870, S0 => 
                           n871);
   U2074 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2891, Z => n1243);
   U2075 : HS65_LH_AO222X4 port map( A => n4619, B => n4549, C => n4615, D => 
                           n4544, E => n1038, F => n2890, Z => n2891);
   U2076 : HS65_LH_HA1X4 port map( A0 => n1208, B0 => n850, CO => n838, S0 => 
                           n839);
   U2077 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2934, Z => n1208);
   U2078 : HS65_LH_AO222X4 port map( A => n4619, B => n4538, C => n4615, D => 
                           n4533, E => n1038, F => n2933, Z => n2934);
   U2079 : HS65_LH_HA1X4 port map( A0 => n1173, B0 => n814, CO => n800, S0 => 
                           n801);
   U2080 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2977, Z => n1173);
   U2081 : HS65_LH_AO222X4 port map( A => n4619, B => n4527, C => n4615, D => 
                           n4522, E => n1038, F => n2976, Z => n2977);
   U2082 : HS65_LH_HA1X4 port map( A0 => n1138, B0 => n772, CO => n756, S0 => 
                           n757);
   U2083 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3020, Z => n1138);
   U2084 : HS65_LH_AO222X4 port map( A => n4619, B => n4516, C => n4615, D => 
                           n4511, E => n1038, F => n3019, Z => n3020);
   U2085 : HS65_LH_HA1X4 port map( A0 => n1103, B0 => n724, CO => n706, S0 => 
                           n707);
   U2086 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3063, Z => n1103);
   U2087 : HS65_LH_AO222X4 port map( A => n4619, B => n4505, C => n4615, D => 
                           n4500, E => n1038, F => n3062, Z => n3063);
   U2088 : HS65_LH_HA1X4 port map( A0 => n1382, B0 => n938, CO => n936, S0 => 
                           n937);
   U2089 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2722, Z => n1382);
   U2090 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1037, D1 => n4581, S1 
                           => n4616, D2 => n4585, S2 => n4618, D3 => n4590, S3 
                           => n4620, Z => n2722);
   U2091 : HS65_LH_HA1X4 port map( A0 => n1347, B0 => n930, CO => n926, S0 => 
                           n927);
   U2092 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2765, Z => n1347);
   U2093 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1037, D1 => n4570, S1 
                           => n4616, D2 => n4574, S2 => n4618, D3 => n4579, S3 
                           => n4620, Z => n2765);
   U2094 : HS65_LH_HA1X4 port map( A0 => n1312, B0 => n916, CO => n910, S0 => 
                           n911);
   U2095 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2807, Z => n1312);
   U2096 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1037, D1 => n4613, S1 
                           => n4620, D2 => n4565, S2 => n4618, D3 => n4562, S3 
                           => n4616, Z => n2807);
   U2097 : HS65_LH_HA1X4 port map( A0 => n1277, B0 => n896, CO => n888, S0 => 
                           n889);
   U2098 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2850, Z => n1277);
   U2099 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1037, D1 => n4551, S1 
                           => n4616, D2 => n4555, S2 => n4618, D3 => n4560, S3 
                           => n4620, Z => n2850);
   U2100 : HS65_LH_HA1X4 port map( A0 => n1242, B0 => n870, CO => n860, S0 => 
                           n861);
   U2101 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2893, Z => n1242);
   U2102 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1037, D1 => n4540, S1 
                           => n4616, D2 => n4544, S2 => n4618, D3 => n4549, S3 
                           => n4620, Z => n2893);
   U2103 : HS65_LH_HA1X4 port map( A0 => n1207, B0 => n838, CO => n826, S0 => 
                           n827);
   U2104 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2936, Z => n1207);
   U2105 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1037, D1 => n4529, S1 
                           => n4616, D2 => n4533, S2 => n4619, D3 => n4538, S3 
                           => n4620, Z => n2936);
   U2106 : HS65_LH_HA1X4 port map( A0 => n1172, B0 => n800, CO => n786, S0 => 
                           n787);
   U2107 : HS65_LHS_XOR2X6 port map( A => a(23), B => n2979, Z => n1172);
   U2108 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1037, D1 => n4527, S1 
                           => n4620, D2 => n4518, S2 => n4617, D3 => n4522, S3 
                           => n4618, Z => n2979);
   U2109 : HS65_LH_HA1X4 port map( A0 => n1137, B0 => n756, CO => n740, S0 => 
                           n741);
   U2110 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3022, Z => n1137);
   U2111 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1037, D1 => n4507, S1 
                           => n4616, D2 => n4511, S2 => n4619, D3 => n4516, S3 
                           => n4620, Z => n3022);
   U2112 : HS65_LH_HA1X4 port map( A0 => n1102, B0 => n706, CO => n688, S0 => 
                           n689);
   U2113 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3065, Z => n1102);
   U2114 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1037, D1 => n4496, S1 
                           => n4616, D2 => n4500, S2 => n4618, D3 => n4505, S3 
                           => n4620, Z => n3065);
   U2115 : HS65_LH_FA1X4 port map( A0 => n1381, B0 => n935, CI => n936, CO => 
                           n932, S0 => n933);
   U2116 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2724, Z => n1381);
   U2117 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1036, D1 => n4581, S1 
                           => n4618, D2 => n4585, S2 => n4621, D3 => n4590, S3 
                           => n4622, Z => n2724);
   U2118 : HS65_LH_FA1X4 port map( A0 => n1346, B0 => n923, CI => n926, CO => 
                           n920, S0 => n921);
   U2119 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2767, Z => n1346);
   U2120 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1036, D1 => n4570, S1 
                           => n4618, D2 => n4574, S2 => n4621, D3 => n4579, S3 
                           => n4622, Z => n2767);
   U2121 : HS65_LH_FA1X4 port map( A0 => n1276, B0 => n881, CI => n888, CO => 
                           n878, S0 => n879);
   U2122 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2852, Z => n1276);
   U2123 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1036, D1 => n4551, S1 
                           => n4618, D2 => n4555, S2 => n4621, D3 => n4560, S3 
                           => n4622, Z => n2852);
   U2124 : HS65_LH_FA1X4 port map( A0 => n1241, B0 => n851, CI => n860, CO => 
                           n848, S0 => n849);
   U2125 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2895, Z => n1241);
   U2126 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1036, D1 => n4540, S1 
                           => n4618, D2 => n4544, S2 => n4621, D3 => n4549, S3 
                           => n4622, Z => n2895);
   U2127 : HS65_LH_FA1X4 port map( A0 => n1206, B0 => n815, CI => n826, CO => 
                           n812, S0 => n813);
   U2128 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2938, Z => n1206);
   U2129 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1036, D1 => n4529, S1 
                           => n4618, D2 => n4532, S2 => n4621, D3 => n4538, S3 
                           => n4622, Z => n2938);
   U2130 : HS65_LH_FA1X4 port map( A0 => n1171, B0 => n773, CI => n786, CO => 
                           n770, S0 => n771);
   U2131 : HS65_LHS_XOR2X6 port map( A => a(23), B => n2981, Z => n1171);
   U2132 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1036, D1 => n4527, S1 
                           => n4622, D2 => n4518, S2 => n4619, D3 => n4522, S3 
                           => n4620, Z => n2981);
   U2133 : HS65_LH_FA1X4 port map( A0 => n1136, B0 => n725, CI => n740, CO => 
                           n722, S0 => n723);
   U2134 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3024, Z => n1136);
   U2135 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1036, D1 => n4507, S1 
                           => n4618, D2 => n4510, S2 => n4621, D3 => n4516, S3 
                           => n4622, Z => n3024);
   U2136 : HS65_LH_FA1X4 port map( A0 => n1311, B0 => n905, CI => n910, CO => 
                           n902, S0 => n903);
   U2137 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2809, Z => n1311);
   U2138 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1036, D1 => n4613, S1 
                           => n4623, D2 => n4565, S2 => n4621, D3 => n4562, S3 
                           => n4618, Z => n2809);
   U2139 : HS65_LH_FA1X4 port map( A0 => n507, B0 => n524, CI => n522, CO => 
                           n504, S0 => n505);
   U2140 : HS65_LH_FA1X4 port map( A0 => n583, B0 => n600, CI => n256, CO => 
                           n255, S0 => product(34));
   U2141 : HS65_LH_FA1X4 port map( A0 => n565, B0 => n582, CI => n255, CO => 
                           n254, S0 => product(35));
   U2142 : HS65_LH_FA1X4 port map( A0 => n503, B0 => n520, CI => n518, CO => 
                           n500, S0 => n501);
   U2143 : HS65_LH_FA1X4 port map( A0 => n513, B0 => n529, CI => n252, CO => 
                           n251, S0 => product(38));
   U2144 : HS65_LH_FA1X4 port map( A0 => n457, B0 => n472, CI => n470, CO => 
                           n454, S0 => n455);
   U2145 : HS65_LH_FA1X4 port map( A0 => n465, B0 => n479, CI => n249, CO => 
                           n248, S0 => product(41));
   U2146 : HS65_LH_FA1X4 port map( A0 => n416, B0 => n429, CI => n427, CO => 
                           n413, S0 => n414);
   U2147 : HS65_LH_FA1X4 port map( A0 => n577, B0 => n594, CI => n592, CO => 
                           n574, S0 => n575);
   U2148 : HS65_LH_FA1X4 port map( A0 => n559, B0 => n576, CI => n574, CO => 
                           n556, S0 => n557);
   U2149 : HS65_LH_FA1X4 port map( A0 => n573, B0 => n590, CI => n588, CO => 
                           n570, S0 => n571);
   U2150 : HS65_LH_FA1X4 port map( A0 => n547, B0 => n564, CI => n254, CO => 
                           n253, S0 => product(36));
   U2151 : HS65_LH_FA1X4 port map( A0 => n461, B0 => n476, CI => n474, CO => 
                           n458, S0 => n459);
   U2152 : HS65_LH_FA1X4 port map( A0 => n499, B0 => n516, CI => n514, CO => 
                           n496, S0 => n497);
   U2153 : HS65_LH_FA1X4 port map( A0 => n495, B0 => n512, CI => n251, CO => 
                           n250, S0 => product(39));
   U2154 : HS65_LH_FA1X4 port map( A0 => n453, B0 => n468, CI => n466, CO => 
                           n450, S0 => n451);
   U2155 : HS65_LH_FA1X4 port map( A0 => n449, B0 => n464, CI => n248, CO => 
                           n247, S0 => product(42));
   U2156 : HS65_LH_FA1X4 port map( A0 => n412, B0 => n425, CI => n423, CO => 
                           n409, S0 => n410);
   U2157 : HS65_LH_FA1X4 port map( A0 => n422, B0 => n434, CI => n246, CO => 
                           n245, S0 => product(44));
   U2158 : HS65_LH_FA1X4 port map( A0 => n382, B0 => n393, CI => n391, CO => 
                           n379, S0 => n380);
   U2159 : HS65_LH_FA1X4 port map( A0 => n408, B0 => n421, CI => n245, CO => 
                           n244, S0 => product(45));
   U2160 : HS65_LH_FA1X4 port map( A0 => n378, B0 => n389, CI => n387, CO => 
                           n375, S0 => n376);
   U2161 : HS65_LH_FA1X4 port map( A0 => n386, B0 => n396, CI => n243, CO => 
                           n242, S0 => product(47));
   U2162 : HS65_LH_FA1X4 port map( A0 => n374, B0 => n385, CI => n242, CO => 
                           n241, S0 => product(48));
   U2163 : HS65_LH_FA1X4 port map( A0 => n349, B0 => n358, CI => n356, CO => 
                           n346, S0 => n347);
   U2164 : HS65_LH_FA1X4 port map( A0 => n355, B0 => n363, CI => n240, CO => 
                           n239, S0 => product(50));
   U2165 : HS65_LH_FA1X4 port map( A0 => n345, B0 => n354, CI => n239, CO => 
                           n238, S0 => product(51));
   U2166 : HS65_LH_FA1X4 port map( A0 => n327, B0 => n334, CI => n332, CO => 
                           n324, S0 => n325);
   U2167 : HS65_LH_FA1X4 port map( A0 => n331, B0 => n337, CI => n237, CO => 
                           n236, S0 => product(53));
   U2168 : HS65_LH_FA1X4 port map( A0 => n312, B0 => n316, CI => n234, CO => 
                           n233, S0 => product(56));
   U2169 : HS65_LH_FA1X4 port map( A0 => n296, B0 => n299, CI => n230, CO => 
                           n229, S0 => product(60));
   U2170 : HS65_LH_FA1X4 port map( A0 => n555, B0 => n572, CI => n570, CO => 
                           n552, S0 => n553);
   U2171 : HS65_LH_FA1X4 port map( A0 => n323, B0 => n330, CI => n236, CO => 
                           n235, S0 => product(54));
   U2172 : HS65_LH_FA1X4 port map( A0 => n306, B0 => n311, CI => n233, CO => 
                           n232, S0 => product(57));
   U2173 : HS65_LH_FA1X4 port map( A0 => n300, B0 => n302, CI => n231, CO => 
                           n230, S0 => product(59));
   U2174 : HS65_LH_FA1X4 port map( A0 => n295, B0 => n294, CI => n229, CO => 
                           n228, S0 => product(61));
   U2175 : HS65_LH_FA1X4 port map( A0 => n4618, B0 => n4620, CI => n1005, CO =>
                           n1004, S0 => n1037);
   U2176 : HS65_LH_FA1X4 port map( A0 => n4620, B0 => n4622, CI => n1004, CO =>
                           n1003, S0 => n1036);
   U2177 : HS65_LH_FA1X4 port map( A0 => n4660, B0 => n4662, CI => n984, CO => 
                           n983, S0 => n1016);
   U2178 : HS65_LH_FA1X4 port map( A0 => n4674, B0 => n4676, CI => n977, CO => 
                           n976, S0 => n1009);
   U2179 : HS65_LH_IVX9 port map( A => n462, Z => n4710);
   U2180 : HS65_LH_IVX9 port map( A => n383, Z => n4711);
   U2181 : HS65_LH_IVX9 port map( A => n328, Z => n4712);
   U2182 : HS65_LH_IVX9 port map( A => n297, Z => n4716);
   U2183 : HS65_LH_IVX9 port map( A => n510, Z => n4709);
   U2184 : HS65_LH_IVX9 port map( A => n419, Z => n4713);
   U2185 : HS65_LH_IVX9 port map( A => n352, Z => n4714);
   U2186 : HS65_LH_IVX9 port map( A => n309, Z => n4715);
   U2187 : HS65_LH_FA1X4 port map( A0 => n4676, B0 => n4678, CI => n976, CO => 
                           n975, S0 => n1008);
   U2188 : HS65_LH_AND2X4 port map( A => n4574, B => n4679, Z => n2800);
   U2189 : HS65_LH_AND2X4 port map( A => n4566, B => n4679, Z => n2842);
   U2190 : HS65_LH_AND2X4 port map( A => n4555, B => n4679, Z => n2885);
   U2191 : HS65_LH_AND2X4 port map( A => n4544, B => n4679, Z => n2928);
   U2192 : HS65_LH_AND2X4 port map( A => n4533, B => n4679, Z => n2971);
   U2193 : HS65_LH_AND2X4 port map( A => n4520, B => n4679, Z => n3014);
   U2194 : HS65_LH_AND2X4 port map( A => n4511, B => n4679, Z => n3057);
   U2195 : HS65_LH_BFX9 port map( A => n4614, Z => n4615);
   U2196 : HS65_LH_BFX9 port map( A => n4614, Z => n4616);
   U2197 : HS65_LH_HA1X4 port map( A0 => n4618, B0 => n4615, CO => n1005, S0 =>
                           n1038);
   U2198 : HS65_LH_BFX9 port map( A => n4614, Z => n4617);
   U2199 : HS65_LH_FA1X4 port map( A0 => n510, B0 => n4687, CI => n1059, CO => 
                           n462, S0 => n493);
   U2200 : HS65_LH_MX41X7 port map( D0 => n1029, S0 => n4491, D1 => n4636, S1 
                           => n4607, D2 => n4634, S2 => n4603, D3 => n4632, S3 
                           => n4609, Z => n1059);
   U2201 : HS65_LH_FA1X4 port map( A0 => n4684, B0 => n4682, CI => n1062, CO =>
                           n510, S0 => n545);
   U2202 : HS65_LH_MX41X7 port map( D0 => n1032, S0 => n4492, D1 => n4630, S1 
                           => n4607, D2 => n4628, S2 => n4603, D3 => n4626, S3 
                           => n4609, Z => n1062);
   U2203 : HS65_LH_FA1X4 port map( A0 => n419, B0 => n4693, CI => n1054, CO => 
                           n383, S0 => n406);
   U2204 : HS65_LH_MX41X7 port map( D0 => n1023, S0 => n4491, D1 => n4644, S1 
                           => n4610, D2 => n4646, S2 => n4603, D3 => n4648, S3 
                           => n4607, Z => n1054);
   U2205 : HS65_LH_FA1X4 port map( A0 => n352, B0 => n4699, CI => n1049, CO => 
                           n328, S0 => n343);
   U2206 : HS65_LH_MX41X7 port map( D0 => n1017, S0 => n4491, D1 => n4656, S1 
                           => n4610, D2 => n4658, S2 => n4603, D3 => n4660, S3 
                           => n4607, Z => n1049);
   U2207 : HS65_LH_FA1X4 port map( A0 => n309, B0 => n4705, CI => n1044, CO => 
                           n297, S0 => n304);
   U2208 : HS65_LH_MX41X7 port map( D0 => n1011, S0 => n4490, D1 => n4668, S1 
                           => n4609, D2 => n4670, S2 => n4603, D3 => n4672, S3 
                           => n4607, Z => n1044);
   U2209 : HS65_LH_FA1X4 port map( A0 => n462, B0 => n4690, CI => n1056, CO => 
                           n446, S0 => n447);
   U2210 : HS65_LH_MX41X7 port map( D0 => n1026, S0 => n4490, D1 => n4606, S1 
                           => n4642, D2 => n4640, S2 => n4602, D3 => n4638, S3 
                           => n4609, Z => n1056);
   U2211 : HS65_LH_FA1X4 port map( A0 => n383, B0 => n4696, CI => n1051, CO => 
                           n371, S0 => n372);
   U2212 : HS65_LH_MX41X7 port map( D0 => n1020, S0 => n4491, D1 => n4650, S1 
                           => n4610, D2 => n4652, S2 => n4603, D3 => n4654, S3 
                           => n4607, Z => n1051);
   U2213 : HS65_LH_FA1X4 port map( A0 => n328, B0 => n4702, CI => n1046, CO => 
                           n320, S0 => n321);
   U2214 : HS65_LH_MX41X7 port map( D0 => n1014, S0 => n4490, D1 => n4662, S1 
                           => n4609, D2 => n4664, S2 => n4602, D3 => n4666, S3 
                           => n4606, Z => n1046);
   U2215 : HS65_LH_FA1X4 port map( A0 => n1194, B0 => n613, CI => n628, CO => 
                           n610, S0 => n611);
   U2216 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2950, Z => n1194);
   U2217 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1024, D1 => n4528, S1 
                           => n4642, D2 => n4531, S2 => n4645, D3 => n4536, S3 
                           => n4646, Z => n2950);
   U2218 : HS65_LH_FA1X4 port map( A0 => n1226, B0 => n611, CI => n626, CO => 
                           n608, S0 => n609);
   U2219 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2910, Z => n1226);
   U2220 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1021, D1 => n4540, S1 
                           => n4649, D2 => n4543, S2 => n4651, D3 => n4548, S3 
                           => n4652, Z => n2910);
   U2221 : HS65_LH_FA1X4 port map( A0 => n1258, B0 => n609, CI => n624, CO => 
                           n606, S0 => n607);
   U2222 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2870, Z => n1258);
   U2223 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1018, D1 => n4550, S1 
                           => n4654, D2 => n4553, S2 => n4657, D3 => n4558, S3 
                           => n4658, Z => n2870);
   U2224 : HS65_LH_FA1X4 port map( A0 => n1290, B0 => n607, CI => n622, CO => 
                           n604, S0 => n605);
   U2225 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2830, Z => n1290);
   U2226 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1015, D1 => n4612, S1 
                           => n4665, D2 => n4564, S2 => n4663, D3 => n4561, S3 
                           => n4660, Z => n2830);
   U2227 : HS65_LH_FA1X4 port map( A0 => n1126, B0 => n544, CI => n560, CO => 
                           n541, S0 => n542);
   U2228 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3034, Z => n1126);
   U2229 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1026, D1 => n4507, S1 
                           => n4639, D2 => n4510, S2 => n4641, D3 => n4515, S3 
                           => n4642, Z => n3034);
   U2230 : HS65_LH_FA1X4 port map( A0 => n1322, B0 => n605, CI => n620, CO => 
                           n602, S0 => n603);
   U2231 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2791, Z => n1322);
   U2232 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1012, D1 => n4569, S1 
                           => n4667, D2 => n4572, S2 => n4669, D3 => n4577, S3 
                           => n4670, Z => n2791);
   U2233 : HS65_LH_FA1X4 port map( A0 => n1158, B0 => n542, CI => n558, CO => 
                           n539, S0 => n540);
   U2234 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2994, Z => n1158);
   U2235 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1023, D1 => n4526, S1 
                           => n4648, D2 => n4518, S2 => n4645, D3 => n4521, S3 
                           => n4646, Z => n2994);
   U2236 : HS65_LH_FA1X4 port map( A0 => n1091, B0 => n493, CI => n508, CO => 
                           n491, S0 => n492);
   U2237 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3077, Z => n1091);
   U2238 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1026, D1 => n4495, S1 
                           => n4639, D2 => n4498, S2 => n4641, D3 => n4504, S3 
                           => n4642, Z => n3077);
   U2239 : HS65_LH_FA1X4 port map( A0 => n1254, B0 => n536, CI => n552, CO => 
                           n533, S0 => n534);
   U2240 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2874, Z => n1254);
   U2241 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1014, D1 => n4550, S1 
                           => n4662, D2 => n4553, S2 => n4665, D3 => n4558, S3 
                           => n4666, Z => n2874);
   U2242 : HS65_LH_FA1X4 port map( A0 => n1155, B0 => n490, CI => n504, CO => 
                           n487, S0 => n488);
   U2243 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2997, Z => n1155);
   U2244 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1020, D1 => n4526, S1 
                           => n4655, D2 => n4518, S2 => n4651, D3 => n4521, S3 
                           => n4652, Z => n2997);
   U2245 : HS65_LH_FA1X4 port map( A0 => n1098, B0 => n1066, CI => n634, CO => 
                           n616, S0 => n617);
   U2246 : HS65_LH_MX41X7 port map( D0 => n1036, S0 => n4492, D1 => n4622, S1 
                           => n4608, D2 => n4620, S2 => n4604, D3 => n4618, S3 
                           => n4609, Z => n1066);
   U2247 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3070, Z => n1098);
   U2248 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1033, D1 => n4496, S1 
                           => n4625, D2 => n4499, S2 => n4627, D3 => n4504, S3 
                           => n4628, Z => n3070);
   U2249 : HS65_LH_FA1X4 port map( A0 => n1130, B0 => n617, CI => n632, CO => 
                           n614, S0 => n615);
   U2250 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3030, Z => n1130);
   U2251 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1030, D1 => n4507, S1 
                           => n4630, D2 => n4510, S2 => n4633, D3 => n4515, S3 
                           => n4634, Z => n3030);
   U2252 : HS65_LH_FA1X4 port map( A0 => n1162, B0 => n615, CI => n630, CO => 
                           n612, S0 => n613);
   U2253 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2990, Z => n1162);
   U2254 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1027, D1 => n4526, S1 
                           => n4640, D2 => n4518, S2 => n4637, D3 => n4521, S3 
                           => n4638, Z => n2990);
   U2255 : HS65_LH_FA1X4 port map( A0 => n1354, B0 => n603, CI => n618, CO => 
                           n600, S0 => n601);
   U2256 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2751, Z => n1354);
   U2257 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1009, D1 => n4580, S1 
                           => n4672, D2 => n4583, S2 => n4675, D3 => n4588, S3 
                           => n4677, Z => n2751);
   U2258 : HS65_LH_FA1X4 port map( A0 => n1190, B0 => n540, CI => n556, CO => 
                           n537, S0 => n538);
   U2259 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2954, Z => n1190);
   U2260 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1020, D1 => n4529, S1 
                           => n4651, D2 => n4532, S2 => n4653, D3 => n4537, S3 
                           => n4654, Z => n2954);
   U2261 : HS65_LH_FA1X4 port map( A0 => n1219, B0 => n486, CI => n500, CO => 
                           n483, S0 => n484);
   U2262 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2917, Z => n1219);
   U2263 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1014, D1 => n4539, S1 
                           => n4663, D2 => n4542, S2 => n4665, D3 => n4547, S3 
                           => n4666, Z => n2917);
   U2264 : HS65_LH_FA1X4 port map( A0 => n1120, B0 => n445, CI => n458, CO => 
                           n442, S0 => n443);
   U2265 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3040, Z => n1120);
   U2266 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1020, D1 => n4507, S1 
                           => n4650, D2 => n4510, S2 => n4653, D3 => n4515, S3 
                           => n4654, Z => n3040);
   U2267 : HS65_LH_FA1X4 port map( A0 => n1184, B0 => n441, CI => n454, CO => 
                           n438, S0 => n439);
   U2268 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2960, Z => n1184);
   U2269 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1014, D1 => n4528, S1 
                           => n4663, D2 => n4531, S2 => n4665, D3 => n4536, S3 
                           => n4666, Z => n2960);
   U2270 : HS65_LH_FA1X4 port map( A0 => n1085, B0 => n406, CI => n417, CO => 
                           n404, S0 => n405);
   U2271 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3083, Z => n1085);
   U2272 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1020, D1 => n4495, S1 
                           => n4651, D2 => n4498, S2 => n4653, D3 => n4503, S3 
                           => n4654, Z => n3083);
   U2273 : HS65_LH_FA1X4 port map( A0 => n1149, B0 => n403, CI => n413, CO => 
                           n400, S0 => n401);
   U2274 : HS65_LHS_XOR2X6 port map( A => n4701, B => n3003, Z => n1149);
   U2275 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1014, D1 => n4526, S1 
                           => n4667, D2 => n4518, S2 => n4663, D3 => n4521, S3 
                           => n4664, Z => n3003);
   U2276 : HS65_LH_FA1X4 port map( A0 => n1114, B0 => n370, CI => n379, CO => 
                           n367, S0 => n368);
   U2277 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3046, Z => n1114);
   U2278 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1014, D1 => n4506, S1 
                           => n4663, D2 => n4509, S2 => n4665, D3 => n4514, S3 
                           => n4666, Z => n3046);
   U2279 : HS65_LH_FA1X4 port map( A0 => n1079, B0 => n343, CI => n350, CO => 
                           n341, S0 => n342);
   U2280 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3089, Z => n1079);
   U2281 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1014, D1 => n4495, S1 
                           => n4663, D2 => n4499, S2 => n4665, D3 => n4503, S3 
                           => n4666, Z => n3089);
   U2282 : HS65_LH_FA1X4 port map( A0 => n597, B0 => n614, CI => n1161, CO => 
                           n594, S0 => n595);
   U2283 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2991, Z => n1161);
   U2284 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1026, D1 => n4525, S1 
                           => n4642, D2 => n4517, S2 => n4639, D3 => n4520, S3 
                           => n4640, Z => n2991);
   U2285 : HS65_LH_FA1X4 port map( A0 => n579, B0 => n1128, CI => n1160, CO => 
                           n576, S0 => n577);
   U2286 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2992, Z => n1160);
   U2287 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3032, Z => n1128);
   U2288 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1025, D1 => n4525, S1 
                           => n4644, D2 => n4517, S2 => n4641, D3 => n4520, S3 
                           => n4642, Z => n2992);
   U2289 : HS65_LH_FA1X4 port map( A0 => n593, B0 => n610, CI => n1225, CO => 
                           n590, S0 => n591);
   U2290 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2911, Z => n1225);
   U2291 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1020, D1 => n4539, S1 
                           => n4650, D2 => n4542, S2 => n4653, D3 => n4547, S3 
                           => n4654, Z => n2911);
   U2292 : HS65_LH_FA1X4 port map( A0 => n562, B0 => n545, CI => n1094, CO => 
                           n543, S0 => n544);
   U2293 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3074, Z => n1094);
   U2294 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1029, D1 => n4496, S1 
                           => n4632, D2 => n4500, S2 => n4635, D3 => n4505, S3 
                           => n4636, Z => n3074);
   U2295 : HS65_LH_FA1X4 port map( A0 => n575, B0 => n1192, CI => n1224, CO => 
                           n572, S0 => n573);
   U2296 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2912, Z => n1224);
   U2297 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2952, Z => n1192);
   U2298 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1019, D1 => n4539, S1 
                           => n4653, D2 => n4542, S2 => n4655, D3 => n4547, S3 
                           => n4656, Z => n2912);
   U2299 : HS65_LH_FA1X4 port map( A0 => n527, B0 => n543, CI => n1125, CO => 
                           n524, S0 => n525);
   U2300 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3035, Z => n1125);
   U2301 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1025, D1 => n4507, S1 
                           => n4640, D2 => n4510, S2 => n4643, D3 => n4515, S3 
                           => n4644, Z => n3035);
   U2302 : HS65_LH_FA1X4 port map( A0 => n554, B0 => n538, CI => n1222, CO => 
                           n535, S0 => n536);
   U2303 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2914, Z => n1222);
   U2304 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1017, D1 => n4539, S1 
                           => n4656, D2 => n4542, S2 => n4659, D3 => n4547, S3 
                           => n4660, Z => n2914);
   U2305 : HS65_LH_FA1X4 port map( A0 => n523, B0 => n539, CI => n1189, CO => 
                           n520, S0 => n521);
   U2306 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2955, Z => n1189);
   U2307 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1019, D1 => n4528, S1 
                           => n4652, D2 => n4531, S2 => n4655, D3 => n4536, S3 
                           => n4656, Z => n2955);
   U2308 : HS65_LH_FA1X4 port map( A0 => n567, B0 => n1320, CI => n1352, CO => 
                           n564, S0 => n565);
   U2309 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2755, Z => n1352);
   U2310 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2793, Z => n1320);
   U2311 : HS65_LH_OAI21X3 port map( A => n4719, B => n4587, C => n2756, Z => 
                           n2755);
   U2312 : HS65_LH_FA1X4 port map( A0 => n506, B0 => n492, CI => n1123, CO => 
                           n489, S0 => n490);
   U2313 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3037, Z => n1123);
   U2314 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1023, D1 => n4507, S1 
                           => n4644, D2 => n4511, S2 => n4647, D3 => n4516, S3 
                           => n4648, Z => n3037);
   U2315 : HS65_LH_FA1X4 port map( A0 => n333, B0 => n339, CI => n1142, CO => 
                           n330, S0 => n331);
   U2316 : HS65_LHS_XOR2X6 port map( A => a(23), B => n3012, Z => n1142);
   U2317 : HS65_LH_OAI21X3 port map( A => n4719, B => n4524, C => n3013, Z => 
                           n3012);
   U2318 : HS65_LH_OAI22X6 port map( A => n4676, B => n3014, C => n4517, D => 
                           n3014, Z => n3013);
   U2319 : HS65_LH_FA1X4 port map( A0 => n314, B0 => n318, CI => n1107, CO => 
                           n311, S0 => n312);
   U2320 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3055, Z => n1107);
   U2321 : HS65_LH_OAI21X3 port map( A => n4719, B => n4513, C => n3056, Z => 
                           n3055);
   U2322 : HS65_LH_OAI22X6 port map( A => n4676, B => n3057, C => n4506, D => 
                           n3057, Z => n3056);
   U2323 : HS65_LH_FA1X4 port map( A0 => n4710, B0 => n1058, CI => n1090, CO =>
                           n476, S0 => n477);
   U2324 : HS65_LH_MX41X7 port map( D0 => n1028, S0 => n4491, D1 => n4638, S1 
                           => n4607, D2 => n4636, S2 => n4603, D3 => n4634, S3 
                           => n4609, Z => n1058);
   U2325 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3078, Z => n1090);
   U2326 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1025, D1 => n4495, S1 
                           => n4640, D2 => n4498, S2 => n4643, D3 => n4503, S3 
                           => n4644, Z => n3078);
   U2327 : HS65_LH_FA1X4 port map( A0 => n550, B0 => n534, CI => n1286, CO => 
                           n531, S0 => n532);
   U2328 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2834, Z => n1286);
   U2329 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1011, D1 => n4613, S1 
                           => n4673, D2 => n4565, S2 => n4671, D3 => n4562, S3 
                           => n4668, Z => n2834);
   U2330 : HS65_LH_FA1X4 port map( A0 => n519, B0 => n535, CI => n1253, CO => 
                           n516, S0 => n517);
   U2331 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2875, Z => n1253);
   U2332 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1013, D1 => n4550, S1 
                           => n4665, D2 => n4553, S2 => n4667, D3 => n4558, S3 
                           => n4668, Z => n2875);
   U2333 : HS65_LH_FA1X4 port map( A0 => n502, B0 => n488, CI => n1187, CO => 
                           n485, S0 => n486);
   U2334 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2957, Z => n1187);
   U2335 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1017, D1 => n4529, S1 
                           => n4656, D2 => n4533, S2 => n4659, D3 => n4538, S3 
                           => n4660, Z => n2957);
   U2336 : HS65_LH_FA1X4 port map( A0 => n475, B0 => n489, CI => n1154, CO => 
                           n472, S0 => n473);
   U2337 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2998, Z => n1154);
   U2338 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1019, D1 => n4525, S1 
                           => n4657, D2 => n4517, S2 => n4653, D3 => n4520, S3 
                           => n4654, Z => n2998);
   U2339 : HS65_LH_FA1X4 port map( A0 => n515, B0 => n531, CI => n1317, CO => 
                           n512, S0 => n513);
   U2340 : HS65_LHS_XOR2X6 port map( A => a(8), B => n2798, Z => n1317);
   U2341 : HS65_LH_OAI21X3 port map( A => n4719, B => n4576, C => n2799, Z => 
                           n2798);
   U2342 : HS65_LH_OAI22X6 port map( A => n4676, B => n2800, C => n4569, D => 
                           n2800, Z => n2799);
   U2343 : HS65_LH_FA1X4 port map( A0 => n460, B0 => n447, CI => n1088, CO => 
                           n444, S0 => n445);
   U2344 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3080, Z => n1088);
   U2345 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1023, D1 => n4496, S1 
                           => n4644, D2 => n4499, S2 => n4647, D3 => n4504, S3 
                           => n4648, Z => n3080);
   U2346 : HS65_LH_FA1X4 port map( A0 => n498, B0 => n484, CI => n1251, CO => 
                           n481, S0 => n482);
   U2347 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2877, Z => n1251);
   U2348 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1011, D1 => n4550, S1 
                           => n4668, D2 => n4553, S2 => n4671, D3 => n4558, S3 
                           => n4672, Z => n2877);
   U2349 : HS65_LH_FA1X4 port map( A0 => n471, B0 => n485, CI => n1218, CO => 
                           n468, S0 => n469);
   U2350 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2918, Z => n1218);
   U2351 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1013, D1 => n4539, S1 
                           => n4664, D2 => n4542, S2 => n4667, D3 => n4547, S3 
                           => n4668, Z => n2918);
   U2352 : HS65_LH_FA1X4 port map( A0 => n456, B0 => n443, CI => n1152, CO => 
                           n440, S0 => n441);
   U2353 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3000, Z => n1152);
   U2354 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1017, D1 => n4527, S1 
                           => n4661, D2 => n4518, S2 => n4657, D3 => n4522, S3 
                           => n4658, Z => n3000);
   U2355 : HS65_LH_FA1X4 port map( A0 => n432, B0 => n444, CI => n1119, CO => 
                           n429, S0 => n430);
   U2356 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3041, Z => n1119);
   U2357 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1019, D1 => n4506, S1 
                           => n4653, D2 => n4509, S2 => n4655, D3 => n4514, S3 
                           => n4656, Z => n3041);
   U2358 : HS65_LH_FA1X4 port map( A0 => n467, B0 => n481, CI => n1282, CO => 
                           n464, S0 => n465);
   U2359 : HS65_LHS_XOR2X6 port map( A => a(11), B => n2840, Z => n1282);
   U2360 : HS65_LH_OAI21X3 port map( A => n4719, B => n4568, C => n2841, Z => 
                           n2840);
   U2361 : HS65_LH_OAI22X6 port map( A => n4676, B => n2842, C => n4561, D => 
                           n2842, Z => n2841);
   U2362 : HS65_LH_FA1X4 port map( A0 => n452, B0 => n439, CI => n1216, CO => 
                           n436, S0 => n437);
   U2363 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2920, Z => n1216);
   U2364 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1011, D1 => n4539, S1 
                           => n4668, D2 => n4542, S2 => n4671, D3 => n4547, S3 
                           => n4672, Z => n2920);
   U2365 : HS65_LH_FA1X4 port map( A0 => n428, B0 => n440, CI => n1183, CO => 
                           n425, S0 => n426);
   U2366 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2961, Z => n1183);
   U2367 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1013, D1 => n4529, S1 
                           => n4664, D2 => n4532, S2 => n4667, D3 => n4537, S3 
                           => n4668, Z => n2961);
   U2368 : HS65_LH_FA1X4 port map( A0 => n415, B0 => n405, CI => n1117, CO => 
                           n402, S0 => n403);
   U2369 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3043, Z => n1117);
   U2370 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1017, D1 => n4506, S1 
                           => n4657, D2 => n4509, S2 => n4659, D3 => n4514, S3 
                           => n4660, Z => n3043);
   U2371 : HS65_LH_FA1X4 port map( A0 => n424, B0 => n436, CI => n1247, CO => 
                           n421, S0 => n422);
   U2372 : HS65_LHS_XOR2X6 port map( A => a(14), B => n2883, Z => n1247);
   U2373 : HS65_LH_OAI21X3 port map( A => n4719, B => n4557, C => n2884, Z => 
                           n2883);
   U2374 : HS65_LH_OAI22X6 port map( A => n4676, B => n2885, C => n4550, D => 
                           n2885, Z => n2884);
   U2375 : HS65_LH_FA1X4 port map( A0 => n4711, B0 => n1053, CI => n1084, CO =>
                           n393, S0 => n394);
   U2376 : HS65_LH_MX41X7 port map( D0 => n1022, S0 => n4491, D1 => n4646, S1 
                           => n4610, D2 => n4648, S2 => n4602, D3 => n4650, S3 
                           => n4606, Z => n1053);
   U2377 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3084, Z => n1084);
   U2378 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1019, D1 => n4495, S1 
                           => n4653, D2 => n4498, S2 => n4655, D3 => n4503, S3 
                           => n4656, Z => n3084);
   U2379 : HS65_LH_FA1X4 port map( A0 => n411, B0 => n401, CI => n1181, CO => 
                           n398, S0 => n399);
   U2380 : HS65_LHS_XOR2X6 port map( A => a(20), B => n2963, Z => n1181);
   U2381 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1011, D1 => n4529, S1 
                           => n4669, D2 => n4532, S2 => n4671, D3 => n4538, S3 
                           => n4672, Z => n2963);
   U2382 : HS65_LH_FA1X4 port map( A0 => n392, B0 => n402, CI => n1148, CO => 
                           n389, S0 => n390);
   U2383 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3004, Z => n1148);
   U2384 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1013, D1 => n4525, S1 
                           => n4669, D2 => n4517, S2 => n4665, D3 => n4520, S3 
                           => n4666, Z => n3004);
   U2385 : HS65_LH_FA1X4 port map( A0 => n381, B0 => n372, CI => n1082, CO => 
                           n369, S0 => n370);
   U2386 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3086, Z => n1082);
   U2387 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1017, D1 => n4496, S1 
                           => n4657, D2 => n4499, S2 => n4659, D3 => n4504, S3 
                           => n4660, Z => n3086);
   U2388 : HS65_LH_FA1X4 port map( A0 => n388, B0 => n398, CI => n1212, CO => 
                           n385, S0 => n386);
   U2389 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2926, Z => n1212);
   U2390 : HS65_LH_OAI21X3 port map( A => n4719, B => n4546, C => n2927, Z => 
                           n2926);
   U2391 : HS65_LH_OAI22X6 port map( A => n4676, B => n2928, C => n4539, D => 
                           n2928, Z => n2927);
   U2392 : HS65_LH_FA1X4 port map( A0 => n377, B0 => n368, CI => n1146, CO => 
                           n365, S0 => n366);
   U2393 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3006, Z => n1146);
   U2394 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1011, D1 => n4525, S1 
                           => n4673, D2 => n4517, S2 => n4669, D3 => n4520, S3 
                           => n4670, Z => n3006);
   U2395 : HS65_LH_FA1X4 port map( A0 => n361, B0 => n369, CI => n1113, CO => 
                           n358, S0 => n359);
   U2396 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3047, Z => n1113);
   U2397 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1013, D1 => n4506, S1 
                           => n4665, D2 => n4509, S2 => n4667, D3 => n4514, S3 
                           => n4668, Z => n3047);
   U2398 : HS65_LH_FA1X4 port map( A0 => n357, B0 => n365, CI => n1177, CO => 
                           n354, S0 => n355);
   U2399 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2969, Z => n1177);
   U2400 : HS65_LH_OAI21X3 port map( A => n4719, B => n4535, C => n2970, Z => 
                           n2969);
   U2401 : HS65_LH_OAI22X6 port map( A => n4676, B => n2971, C => n4528, D => 
                           n2971, Z => n2970);
   U2402 : HS65_LH_FA1X4 port map( A0 => n348, B0 => n342, CI => n1111, CO => 
                           n339, S0 => n340);
   U2403 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3049, Z => n1111);
   U2404 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1011, D1 => n4506, S1 
                           => n4669, D2 => n4509, S2 => n4671, D3 => n4514, S3 
                           => n4672, Z => n3049);
   U2405 : HS65_LH_FA1X4 port map( A0 => n4712, B0 => n1048, CI => n1078, CO =>
                           n334, S0 => n335);
   U2406 : HS65_LH_MX41X7 port map( D0 => n1016, S0 => n4491, D1 => n4658, S1 
                           => n4610, D2 => n4660, S2 => n4602, D3 => n4662, S3 
                           => n4606, Z => n1048);
   U2407 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3090, Z => n1078);
   U2408 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1013, D1 => n4495, S1 
                           => n4665, D2 => n4498, S2 => n4667, D3 => n4503, S3 
                           => n4668, Z => n3090);
   U2409 : HS65_LH_FA1X4 port map( A0 => n326, B0 => n321, CI => n1076, CO => 
                           n318, S0 => n319);
   U2410 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3092, Z => n1076);
   U2411 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1011, D1 => n4496, S1 
                           => n4668, D2 => n4499, S2 => n4671, D3 => n4504, S3 
                           => n4672, Z => n3092);
   U2412 : HS65_LH_FA1X4 port map( A0 => n4716, B0 => n1043, CI => n1072, CO =>
                           n299, S0 => n300);
   U2413 : HS65_LH_MX41X7 port map( D0 => n1010, S0 => n4491, D1 => n4670, S1 
                           => n4610, D2 => n4672, S2 => n4603, D3 => n4674, S3 
                           => n4607, Z => n1043);
   U2414 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3098, Z => n1072);
   U2415 : HS65_LH_OAI21X3 port map( A => n4719, B => n4502, C => n3099, Z => 
                           n3098);
   U2416 : HS65_LH_FA1X4 port map( A0 => n293, B0 => n292, CI => n228, CO => 
                           n227, S0 => product(62));
   U2417 : HS65_LH_HA1X4 port map( A0 => n4680, B0 => n1419, CO => n289, S0 => 
                           product(0));
   U2418 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2676, Z => n1419);
   U2419 : HS65_LH_AO22X9 port map( A => n4616, B => n4600, C => n4493, D => 
                           n4616, Z => n2676);
   U2420 : HS65_LH_HA1X4 port map( A0 => n1418, B0 => n289, CO => n288, S0 => 
                           product(1));
   U2421 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2678, Z => n1418);
   U2422 : HS65_LH_AO222X4 port map( A => n4617, B => n4596, C => n4598, D => 
                           n4619, E => n4493, F => n1038, Z => n2678);
   U2423 : HS65_LH_IVX9 port map( A => n4687, Z => n4685);
   U2424 : HS65_LH_IVX9 port map( A => n4693, Z => n4692);
   U2425 : HS65_LH_IVX9 port map( A => n4687, Z => n4686);
   U2426 : HS65_LH_IVX9 port map( A => n4693, Z => n4691);
   U2427 : HS65_LH_IVX9 port map( A => n4696, Z => n4695);
   U2428 : HS65_LH_IVX9 port map( A => n4696, Z => n4694);
   U2429 : HS65_LH_IVX9 port map( A => n4708, Z => n4706);
   U2430 : HS65_LH_IVX9 port map( A => n4708, Z => n4707);
   U2431 : HS65_LH_IVX9 port map( A => n4699, Z => n4697);
   U2432 : HS65_LH_IVX9 port map( A => n4699, Z => n4698);
   U2433 : HS65_LH_IVX9 port map( A => n4690, Z => n4688);
   U2434 : HS65_LH_IVX9 port map( A => n4690, Z => n4689);
   U2435 : HS65_LH_IVX9 port map( A => n4705, Z => n4704);
   U2436 : HS65_LH_IVX9 port map( A => n4705, Z => n4703);
   U2437 : HS65_LH_IVX9 port map( A => n4702, Z => n4700);
   U2438 : HS65_LH_IVX9 port map( A => n4702, Z => n4701);
   U2439 : HS65_LH_MX41X7 port map( D0 => n1025, S0 => n4491, D1 => n4644, S1 
                           => n4607, D2 => n4642, S2 => n4603, D3 => n4640, S3 
                           => n4609, Z => n419);
   U2440 : HS65_LH_MX41X7 port map( D0 => n1019, S0 => n4491, D1 => n4652, S1 
                           => n4610, D2 => n4654, S2 => n4603, D3 => n4656, S3 
                           => n4607, Z => n352);
   U2441 : HS65_LH_MX41X7 port map( D0 => n1013, S0 => n4490, D1 => n4664, S1 
                           => n4610, D2 => n4666, S2 => n4602, D3 => n4668, S3 
                           => n4606, Z => n309);
   U2442 : HS65_LH_IVX9 port map( A => n4684, Z => n4683);
   U2443 : HS65_LH_IVX9 port map( A => a(5), Z => n4684);
   U2444 : HS65_LH_HA1X4 port map( A0 => n1417, B0 => n288, CO => n287, S0 => 
                           product(2));
   U2445 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2680, Z => n1417);
   U2446 : HS65_LH_MX41X7 port map( D0 => n1037, S0 => n4493, D1 => n4591, S1 
                           => n4616, D2 => n4594, S2 => n4619, D3 => n4620, S3 
                           => n4598, Z => n2680);
   U2447 : HS65_LH_FA1X4 port map( A0 => n1416, B0 => n941, CI => n287, CO => 
                           n286, S0 => product(3));
   U2448 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2682, Z => n1416);
   U2449 : HS65_LH_MX41X7 port map( D0 => n1036, S0 => n4493, D1 => n4591, S1 
                           => n4618, D2 => n4620, S2 => n4595, D3 => n4622, S3 
                           => n4599, Z => n2682);
   U2450 : HS65_LH_FA1X4 port map( A0 => n1415, B0 => n939, CI => n286, CO => 
                           n285, S0 => product(4));
   U2451 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2683, Z => n1415);
   U2452 : HS65_LH_MX41X7 port map( D0 => n1035, S0 => n4493, D1 => n4591, S1 
                           => n4621, D2 => n4622, S2 => n4595, D3 => n4624, S3 
                           => n4599, Z => n2683);
   U2453 : HS65_LH_FA1X4 port map( A0 => n1414, B0 => n937, CI => n285, CO => 
                           n284, S0 => product(5));
   U2454 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2684, Z => n1414);
   U2455 : HS65_LH_MX41X7 port map( D0 => n1034, S0 => n4494, D1 => n4622, S1 
                           => n4592, D2 => n4624, S2 => n4596, D3 => n4626, S3 
                           => n4600, Z => n2684);
   U2456 : HS65_LH_FA1X4 port map( A0 => n1413, B0 => n933, CI => n284, CO => 
                           n283, S0 => product(6));
   U2457 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2685, Z => n1413);
   U2458 : HS65_LH_MX41X7 port map( D0 => n1033, S0 => n4493, D1 => n4624, S1 
                           => n4592, D2 => n4626, S2 => n4595, D3 => n4628, S3 
                           => n4599, Z => n2685);
   U2459 : HS65_LH_FA1X4 port map( A0 => n1380, B0 => n931, CI => n932, CO => 
                           n928, S0 => n929);
   U2460 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2725, Z => n1380);
   U2461 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1035, D1 => n4581, S1 
                           => n4621, D2 => n4584, S2 => n4623, D3 => n4590, S3 
                           => n4624, Z => n2725);
   U2462 : HS65_LH_FA1X4 port map( A0 => n1412, B0 => n929, CI => n283, CO => 
                           n282, S0 => product(7));
   U2463 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2686, Z => n1412);
   U2464 : HS65_LH_MX41X7 port map( D0 => n1032, S0 => n4493, D1 => n4626, S1 
                           => n4592, D2 => n4628, S2 => n4595, D3 => n4630, S3 
                           => n4599, Z => n2686);
   U2465 : HS65_LH_FA1X4 port map( A0 => n1379, B0 => n927, CI => n928, CO => 
                           n924, S0 => n925);
   U2466 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2726, Z => n1379);
   U2467 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1034, D1 => n4580, S1 
                           => n4622, D2 => n4585, S2 => n4625, D3 => n4590, S3 
                           => n4626, Z => n2726);
   U2468 : HS65_LH_FA1X4 port map( A0 => n1411, B0 => n925, CI => n282, CO => 
                           n281, S0 => product(8));
   U2469 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2687, Z => n1411);
   U2470 : HS65_LH_MX41X7 port map( D0 => n1031, S0 => n4493, D1 => n4628, S1 
                           => n4592, D2 => n4630, S2 => n4595, D3 => n4632, S3 
                           => n4599, Z => n2687);
   U2471 : HS65_LH_FA1X4 port map( A0 => n1345, B0 => n917, CI => n920, CO => 
                           n914, S0 => n915);
   U2472 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2768, Z => n1345);
   U2473 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1035, D1 => n4570, S1 
                           => n4621, D2 => n4573, S2 => n4623, D3 => n4579, S3 
                           => n4624, Z => n2768);
   U2474 : HS65_LH_FA1X4 port map( A0 => n1378, B0 => n921, CI => n924, CO => 
                           n918, S0 => n919);
   U2475 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2727, Z => n1378);
   U2476 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1033, D1 => n4580, S1 
                           => n4624, D2 => n4583, S2 => n4627, D3 => n4588, S3 
                           => n4628, Z => n2727);
   U2477 : HS65_LH_FA1X4 port map( A0 => n1410, B0 => n919, CI => n281, CO => 
                           n280, S0 => product(9));
   U2478 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2688, Z => n1410);
   U2479 : HS65_LH_MX41X7 port map( D0 => n1030, S0 => n4493, D1 => n4630, S1 
                           => n4591, D2 => n4632, S2 => n4595, D3 => n4634, S3 
                           => n4599, Z => n2688);
   U2480 : HS65_LH_FA1X4 port map( A0 => n1344, B0 => n911, CI => n914, CO => 
                           n908, S0 => n909);
   U2481 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2769, Z => n1344);
   U2482 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1034, D1 => n4569, S1 
                           => n4623, D2 => n4574, S2 => n4625, D3 => n4579, S3 
                           => n4626, Z => n2769);
   U2483 : HS65_LH_FA1X4 port map( A0 => n1377, B0 => n915, CI => n918, CO => 
                           n912, S0 => n913);
   U2484 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2728, Z => n1377);
   U2485 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1032, D1 => n4580, S1 
                           => n4627, D2 => n4583, S2 => n4629, D3 => n4588, S3 
                           => n4630, Z => n2728);
   U2486 : HS65_LH_FA1X4 port map( A0 => n1409, B0 => n913, CI => n280, CO => 
                           n279, S0 => product(10));
   U2487 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2689, Z => n1409);
   U2488 : HS65_LH_MX41X7 port map( D0 => n1029, S0 => n4493, D1 => n4632, S1 
                           => n4592, D2 => n4634, S2 => n4595, D3 => n4636, S3 
                           => n4599, Z => n2689);
   U2489 : HS65_LH_FA1X4 port map( A0 => n1310, B0 => n897, CI => n902, CO => 
                           n894, S0 => n895);
   U2490 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2810, Z => n1310);
   U2491 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1035, D1 => n4612, S1 
                           => n4624, D2 => n4565, S2 => n4623, D3 => n4562, S3 
                           => n4620, Z => n2810);
   U2492 : HS65_LH_FA1X4 port map( A0 => n1343, B0 => n903, CI => n908, CO => 
                           n900, S0 => n901);
   U2493 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2770, Z => n1343);
   U2494 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1033, D1 => n4569, S1 
                           => n4624, D2 => n4572, S2 => n4627, D3 => n4577, S3 
                           => n4628, Z => n2770);
   U2495 : HS65_LH_FA1X4 port map( A0 => n1376, B0 => n909, CI => n912, CO => 
                           n906, S0 => n907);
   U2496 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2729, Z => n1376);
   U2497 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1031, D1 => n4580, S1 
                           => n4629, D2 => n4583, S2 => n4631, D3 => n4588, S3 
                           => n4632, Z => n2729);
   U2498 : HS65_LH_FA1X4 port map( A0 => n1408, B0 => n907, CI => n279, CO => 
                           n278, S0 => product(11));
   U2499 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2690, Z => n1408);
   U2500 : HS65_LH_MX41X7 port map( D0 => n1028, S0 => n4493, D1 => n4634, S1 
                           => n4592, D2 => n4636, S2 => n4595, D3 => n4638, S3 
                           => n4599, Z => n2690);
   U2501 : HS65_LH_FA1X4 port map( A0 => n1309, B0 => n889, CI => n894, CO => 
                           n886, S0 => n887);
   U2502 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2811, Z => n1309);
   U2503 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1034, D1 => n4613, S1 
                           => n4626, D2 => n4566, S2 => n4625, D3 => n4561, S3 
                           => n4622, Z => n2811);
   U2504 : HS65_LH_FA1X4 port map( A0 => n1342, B0 => n895, CI => n900, CO => 
                           n892, S0 => n893);
   U2505 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2771, Z => n1342);
   U2506 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1032, D1 => n4569, S1 
                           => n4627, D2 => n4572, S2 => n4629, D3 => n4577, S3 
                           => n4630, Z => n2771);
   U2507 : HS65_LH_FA1X4 port map( A0 => n1375, B0 => n901, CI => n906, CO => 
                           n898, S0 => n899);
   U2508 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2730, Z => n1375);
   U2509 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1030, D1 => n4580, S1 
                           => n4631, D2 => n4583, S2 => n4633, D3 => n4588, S3 
                           => n4634, Z => n2730);
   U2510 : HS65_LH_FA1X4 port map( A0 => n1407, B0 => n899, CI => n278, CO => 
                           n277, S0 => product(12));
   U2511 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2691, Z => n1407);
   U2512 : HS65_LH_MX41X7 port map( D0 => n1027, S0 => n4494, D1 => n4636, S1 
                           => n4592, D2 => n4638, S2 => n4595, D3 => n4598, S3 
                           => n4640, Z => n2691);
   U2513 : HS65_LH_FA1X4 port map( A0 => n1275, B0 => n871, CI => n878, CO => 
                           n868, S0 => n869);
   U2514 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2853, Z => n1275);
   U2515 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1035, D1 => n4551, S1 
                           => n4621, D2 => n4554, S2 => n4623, D3 => n4560, S3 
                           => n4624, Z => n2853);
   U2516 : HS65_LH_FA1X4 port map( A0 => n1308, B0 => n879, CI => n886, CO => 
                           n876, S0 => n877);
   U2517 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2812, Z => n1308);
   U2518 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1033, D1 => n4611, S1 
                           => n4629, D2 => n4564, S2 => n4627, D3 => n4561, S3 
                           => n4624, Z => n2812);
   U2519 : HS65_LH_FA1X4 port map( A0 => n1341, B0 => n887, CI => n892, CO => 
                           n884, S0 => n885);
   U2520 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2772, Z => n1341);
   U2521 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1031, D1 => n4569, S1 
                           => n4629, D2 => n4572, S2 => n4631, D3 => n4577, S3 
                           => n4632, Z => n2772);
   U2522 : HS65_LH_FA1X4 port map( A0 => n1374, B0 => n893, CI => n898, CO => 
                           n890, S0 => n891);
   U2523 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2731, Z => n1374);
   U2524 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1029, D1 => n4580, S1 
                           => n4633, D2 => n4583, S2 => n4635, D3 => n4588, S3 
                           => n4636, Z => n2731);
   U2525 : HS65_LH_FA1X4 port map( A0 => n1406, B0 => n891, CI => n277, CO => 
                           n276, S0 => product(13));
   U2526 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2692, Z => n1406);
   U2527 : HS65_LH_MX41X7 port map( D0 => n1026, S0 => n4493, D1 => n4638, S1 
                           => n4591, D2 => n4594, S2 => n4641, D3 => n4598, S3 
                           => n4642, Z => n2692);
   U2528 : HS65_LH_FA1X4 port map( A0 => n1274, B0 => n861, CI => n868, CO => 
                           n858, S0 => n859);
   U2529 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2854, Z => n1274);
   U2530 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1034, D1 => n4550, S1 
                           => n4623, D2 => n4555, S2 => n4625, D3 => n4560, S3 
                           => n4626, Z => n2854);
   U2531 : HS65_LH_FA1X4 port map( A0 => n1307, B0 => n869, CI => n876, CO => 
                           n866, S0 => n867);
   U2532 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2813, Z => n1307);
   U2533 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1032, D1 => n4611, S1 
                           => n4631, D2 => n4564, S2 => n4629, D3 => n4561, S3 
                           => n4626, Z => n2813);
   U2534 : HS65_LH_FA1X4 port map( A0 => n1340, B0 => n877, CI => n884, CO => 
                           n874, S0 => n875);
   U2535 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2773, Z => n1340);
   U2536 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1030, D1 => n4569, S1 
                           => n4631, D2 => n4572, S2 => n4633, D3 => n4577, S3 
                           => n4634, Z => n2773);
   U2537 : HS65_LH_FA1X4 port map( A0 => n1373, B0 => n885, CI => n890, CO => 
                           n882, S0 => n883);
   U2538 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2732, Z => n1373);
   U2539 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1028, D1 => n4580, S1 
                           => n4635, D2 => n4583, S2 => n4637, D3 => n4588, S3 
                           => n4638, Z => n2732);
   U2540 : HS65_LH_FA1X4 port map( A0 => n1405, B0 => n883, CI => n276, CO => 
                           n275, S0 => product(14));
   U2541 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2693, Z => n1405);
   U2542 : HS65_LH_MX41X7 port map( D0 => n4493, S0 => n1025, D1 => n4591, S1 
                           => n4641, D2 => n4594, S2 => n4643, D3 => n4598, S3 
                           => n4644, Z => n2693);
   U2543 : HS65_LH_FA1X4 port map( A0 => n1240, B0 => n839, CI => n848, CO => 
                           n836, S0 => n837);
   U2544 : HS65_LHS_XOR2X6 port map( A => a(17), B => n2896, Z => n1240);
   U2545 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1035, D1 => n4540, S1 
                           => n4621, D2 => n4543, S2 => n4623, D3 => n4549, S3 
                           => n4624, Z => n2896);
   U2546 : HS65_LH_FA1X4 port map( A0 => n1273, B0 => n849, CI => n858, CO => 
                           n846, S0 => n847);
   U2547 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2855, Z => n1273);
   U2548 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1033, D1 => n4551, S1 
                           => n4625, D2 => n4554, S2 => n4627, D3 => n4559, S3 
                           => n4628, Z => n2855);
   U2549 : HS65_LH_FA1X4 port map( A0 => n1306, B0 => n859, CI => n866, CO => 
                           n856, S0 => n857);
   U2550 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2814, Z => n1306);
   U2551 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1031, D1 => n4611, S1 
                           => n4633, D2 => n4564, S2 => n4631, D3 => n4561, S3 
                           => n4628, Z => n2814);
   U2552 : HS65_LH_FA1X4 port map( A0 => n1339, B0 => n867, CI => n874, CO => 
                           n864, S0 => n865);
   U2553 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2774, Z => n1339);
   U2554 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1029, D1 => n4569, S1 
                           => n4633, D2 => n4572, S2 => n4635, D3 => n4577, S3 
                           => n4636, Z => n2774);
   U2555 : HS65_LH_FA1X4 port map( A0 => n1372, B0 => n875, CI => n882, CO => 
                           n872, S0 => n873);
   U2556 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2733, Z => n1372);
   U2557 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1027, D1 => n4581, S1 
                           => n4637, D2 => n4584, S2 => n4639, D3 => n4590, S3 
                           => n4640, Z => n2733);
   U2558 : HS65_LH_FA1X4 port map( A0 => n1404, B0 => n873, CI => n275, CO => 
                           n274, S0 => product(15));
   U2559 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2694, Z => n1404);
   U2560 : HS65_LH_MX41X7 port map( D0 => n1024, S0 => n4494, D1 => n4591, S1 
                           => n4643, D2 => n4594, S2 => n4645, D3 => n4646, S3 
                           => n4599, Z => n2694);
   U2561 : HS65_LH_FA1X4 port map( A0 => n1239, B0 => n827, CI => n836, CO => 
                           n824, S0 => n825);
   U2562 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2897, Z => n1239);
   U2563 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1034, D1 => n4539, S1 
                           => n4623, D2 => n4544, S2 => n4625, D3 => n4549, S3 
                           => n4626, Z => n2897);
   U2564 : HS65_LH_FA1X4 port map( A0 => n1272, B0 => n837, CI => n846, CO => 
                           n834, S0 => n835);
   U2565 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2856, Z => n1272);
   U2566 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1032, D1 => n4550, S1 
                           => n4627, D2 => n4554, S2 => n4629, D3 => n4559, S3 
                           => n4630, Z => n2856);
   U2567 : HS65_LH_FA1X4 port map( A0 => n1305, B0 => n847, CI => n856, CO => 
                           n844, S0 => n845);
   U2568 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2815, Z => n1305);
   U2569 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1030, D1 => n4611, S1 
                           => n4635, D2 => n4564, S2 => n4633, D3 => n4561, S3 
                           => n4630, Z => n2815);
   U2570 : HS65_LH_FA1X4 port map( A0 => n1338, B0 => n857, CI => n864, CO => 
                           n854, S0 => n855);
   U2571 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2775, Z => n1338);
   U2572 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1028, D1 => n4569, S1 
                           => n4635, D2 => n4572, S2 => n4637, D3 => n4577, S3 
                           => n4638, Z => n2775);
   U2573 : HS65_LH_FA1X4 port map( A0 => n1371, B0 => n865, CI => n872, CO => 
                           n862, S0 => n863);
   U2574 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2734, Z => n1371);
   U2575 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1026, D1 => n4581, S1 
                           => n4638, D2 => n4584, S2 => n4641, D3 => n4589, S3 
                           => n4642, Z => n2734);
   U2576 : HS65_LH_FA1X4 port map( A0 => n1403, B0 => n863, CI => n274, CO => 
                           n273, S0 => product(16));
   U2577 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2695, Z => n1403);
   U2578 : HS65_LH_MX41X7 port map( D0 => n1023, S0 => n4493, D1 => n4591, S1 
                           => n4645, D2 => n4646, S2 => n4595, D3 => n4648, S3 
                           => n4599, Z => n2695);
   U2579 : HS65_LH_FA1X4 port map( A0 => n1205, B0 => n801, CI => n812, CO => 
                           n798, S0 => n799);
   U2580 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2939, Z => n1205);
   U2581 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1035, D1 => n4529, S1 
                           => n4620, D2 => n4532, S2 => n4623, D3 => n4537, S3 
                           => n4624, Z => n2939);
   U2582 : HS65_LH_FA1X4 port map( A0 => n1238, B0 => n813, CI => n824, CO => 
                           n810, S0 => n811);
   U2583 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2898, Z => n1238);
   U2584 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1033, D1 => n4540, S1 
                           => n4625, D2 => n4543, S2 => n4627, D3 => n4548, S3 
                           => n4628, Z => n2898);
   U2585 : HS65_LH_FA1X4 port map( A0 => n1271, B0 => n825, CI => n834, CO => 
                           n822, S0 => n823);
   U2586 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2857, Z => n1271);
   U2587 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1031, D1 => n4550, S1 
                           => n4628, D2 => n4553, S2 => n4631, D3 => n4559, S3 
                           => n4632, Z => n2857);
   U2588 : HS65_LH_FA1X4 port map( A0 => n1304, B0 => n835, CI => n844, CO => 
                           n832, S0 => n833);
   U2589 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2816, Z => n1304);
   U2590 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1029, D1 => n4611, S1 
                           => n4637, D2 => n4564, S2 => n4635, D3 => n4561, S3 
                           => n4632, Z => n2816);
   U2591 : HS65_LH_FA1X4 port map( A0 => n1337, B0 => n845, CI => n854, CO => 
                           n842, S0 => n843);
   U2592 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2776, Z => n1337);
   U2593 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1027, D1 => n4570, S1 
                           => n4637, D2 => n4573, S2 => n4639, D3 => n4578, S3 
                           => n4640, Z => n2776);
   U2594 : HS65_LH_FA1X4 port map( A0 => n1370, B0 => n855, CI => n862, CO => 
                           n852, S0 => n853);
   U2595 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2735, Z => n1370);
   U2596 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1025, D1 => n4581, S1 
                           => n4641, D2 => n4584, S2 => n4643, D3 => n4589, S3 
                           => n4644, Z => n2735);
   U2597 : HS65_LH_FA1X4 port map( A0 => n1402, B0 => n853, CI => n273, CO => 
                           n272, S0 => product(17));
   U2598 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2696, Z => n1402);
   U2599 : HS65_LH_MX41X7 port map( D0 => n1022, S0 => n4493, D1 => n4646, S1 
                           => n4592, D2 => n4648, S2 => n4595, D3 => n4650, S3 
                           => n4598, Z => n2696);
   U2600 : HS65_LH_FA1X4 port map( A0 => n1237, B0 => n799, CI => n810, CO => 
                           n796, S0 => n797);
   U2601 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2899, Z => n1237);
   U2602 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1032, D1 => n4540, S1 
                           => n4627, D2 => n4543, S2 => n4629, D3 => n4548, S3 
                           => n4630, Z => n2899);
   U2603 : HS65_LH_FA1X4 port map( A0 => n1270, B0 => n811, CI => n822, CO => 
                           n808, S0 => n809);
   U2604 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2858, Z => n1270);
   U2605 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1030, D1 => n4550, S1 
                           => n4631, D2 => n4553, S2 => n4633, D3 => n4558, S3 
                           => n4634, Z => n2858);
   U2606 : HS65_LH_FA1X4 port map( A0 => n1303, B0 => n823, CI => n832, CO => 
                           n820, S0 => n821);
   U2607 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2817, Z => n1303);
   U2608 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1028, D1 => n4611, S1 
                           => n4638, D2 => n4564, S2 => n4637, D3 => n4561, S3 
                           => n4634, Z => n2817);
   U2609 : HS65_LH_FA1X4 port map( A0 => n1336, B0 => n833, CI => n842, CO => 
                           n830, S0 => n831);
   U2610 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2777, Z => n1336);
   U2611 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1026, D1 => n4570, S1 
                           => n4639, D2 => n4573, S2 => n4641, D3 => n4578, S3 
                           => n4642, Z => n2777);
   U2612 : HS65_LH_FA1X4 port map( A0 => n1369, B0 => n843, CI => n852, CO => 
                           n840, S0 => n841);
   U2613 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2736, Z => n1369);
   U2614 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1024, D1 => n4580, S1 
                           => n4643, D2 => n4583, S2 => n4645, D3 => n4588, S3 
                           => n4646, Z => n2736);
   U2615 : HS65_LH_FA1X4 port map( A0 => n1401, B0 => n841, CI => n272, CO => 
                           n271, S0 => product(18));
   U2616 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2697, Z => n1401);
   U2617 : HS65_LH_MX41X7 port map( D0 => n1021, S0 => n4493, D1 => n4648, S1 
                           => n4591, D2 => n4650, S2 => n4594, D3 => n4598, S3 
                           => n4652, Z => n2697);
   U2618 : HS65_LH_FA1X4 port map( A0 => n1170, B0 => n757, CI => n770, CO => 
                           n754, S0 => n755);
   U2619 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2982, Z => n1170);
   U2620 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1035, D1 => n4527, S1 
                           => n4625, D2 => n4518, S2 => n4621, D3 => n4521, S3 
                           => n4622, Z => n2982);
   U2621 : HS65_LH_FA1X4 port map( A0 => n1203, B0 => n771, CI => n784, CO => 
                           n768, S0 => n769);
   U2622 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2941, Z => n1203);
   U2623 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1033, D1 => n4529, S1 
                           => n4625, D2 => n4532, S2 => n4627, D3 => n4537, S3 
                           => n4628, Z => n2941);
   U2624 : HS65_LH_FA1X4 port map( A0 => n1236, B0 => n785, CI => n796, CO => 
                           n782, S0 => n783);
   U2625 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2900, Z => n1236);
   U2626 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1031, D1 => n4540, S1 
                           => n4628, D2 => n4543, S2 => n4631, D3 => n4548, S3 
                           => n4632, Z => n2900);
   U2627 : HS65_LH_FA1X4 port map( A0 => n1269, B0 => n797, CI => n808, CO => 
                           n794, S0 => n795);
   U2628 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2859, Z => n1269);
   U2629 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1029, D1 => n4550, S1 
                           => n4633, D2 => n4553, S2 => n4635, D3 => n4558, S3 
                           => n4636, Z => n2859);
   U2630 : HS65_LH_FA1X4 port map( A0 => n1302, B0 => n809, CI => n820, CO => 
                           n806, S0 => n807);
   U2631 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2818, Z => n1302);
   U2632 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1027, D1 => n4612, S1 
                           => n4640, D2 => n4565, S2 => n4639, D3 => n4562, S3 
                           => n4636, Z => n2818);
   U2633 : HS65_LH_FA1X4 port map( A0 => n1335, B0 => n821, CI => n830, CO => 
                           n818, S0 => n819);
   U2634 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2778, Z => n1335);
   U2635 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1025, D1 => n4570, S1 
                           => n4641, D2 => n4573, S2 => n4643, D3 => n4578, S3 
                           => n4644, Z => n2778);
   U2636 : HS65_LH_FA1X4 port map( A0 => n1368, B0 => n831, CI => n840, CO => 
                           n828, S0 => n829);
   U2637 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2737, Z => n1368);
   U2638 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1023, D1 => n4581, S1 
                           => n4645, D2 => n4584, S2 => n4647, D3 => n4589, S3 
                           => n4648, Z => n2737);
   U2639 : HS65_LH_FA1X4 port map( A0 => n1400, B0 => n829, CI => n271, CO => 
                           n270, S0 => product(19));
   U2640 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2698, Z => n1400);
   U2641 : HS65_LH_MX41X7 port map( D0 => n1020, S0 => n4494, D1 => n4650, S1 
                           => n4592, D2 => n4594, S2 => n4653, D3 => n4598, S3 
                           => n4654, Z => n2698);
   U2642 : HS65_LH_FA1X4 port map( A0 => n1169, B0 => n741, CI => n754, CO => 
                           n738, S0 => n739);
   U2643 : HS65_LHS_XOR2X6 port map( A => a(23), B => n2983, Z => n1169);
   U2644 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1034, D1 => n4527, S1 
                           => n4627, D2 => n4517, S2 => n4623, D3 => n4522, S3 
                           => n4624, Z => n2983);
   U2645 : HS65_LH_FA1X4 port map( A0 => n1202, B0 => n755, CI => n768, CO => 
                           n752, S0 => n753);
   U2646 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2942, Z => n1202);
   U2647 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1032, D1 => n4528, S1 
                           => n4626, D2 => n4532, S2 => n4629, D3 => n4537, S3 
                           => n4630, Z => n2942);
   U2648 : HS65_LH_FA1X4 port map( A0 => n1235, B0 => n769, CI => n782, CO => 
                           n766, S0 => n767);
   U2649 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2901, Z => n1235);
   U2650 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1030, D1 => n4540, S1 
                           => n4631, D2 => n4543, S2 => n4633, D3 => n4548, S3 
                           => n4634, Z => n2901);
   U2651 : HS65_LH_FA1X4 port map( A0 => n1268, B0 => n783, CI => n794, CO => 
                           n780, S0 => n781);
   U2652 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2860, Z => n1268);
   U2653 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1028, D1 => n4550, S1 
                           => n4635, D2 => n4553, S2 => n4637, D3 => n4558, S3 
                           => n4638, Z => n2860);
   U2654 : HS65_LH_FA1X4 port map( A0 => n1301, B0 => n795, CI => n806, CO => 
                           n792, S0 => n793);
   U2655 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2819, Z => n1301);
   U2656 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1026, D1 => n4612, S1 
                           => n4642, D2 => n4565, S2 => n4641, D3 => n4562, S3 
                           => n4638, Z => n2819);
   U2657 : HS65_LH_FA1X4 port map( A0 => n1334, B0 => n807, CI => n818, CO => 
                           n804, S0 => n805);
   U2658 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2779, Z => n1334);
   U2659 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1024, D1 => n4569, S1 
                           => n4643, D2 => n4572, S2 => n4645, D3 => n4577, S3 
                           => n4646, Z => n2779);
   U2660 : HS65_LH_FA1X4 port map( A0 => n1367, B0 => n819, CI => n828, CO => 
                           n816, S0 => n817);
   U2661 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2738, Z => n1367);
   U2662 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1022, D1 => n4581, S1 
                           => n4646, D2 => n4584, S2 => n4649, D3 => n4589, S3 
                           => n4650, Z => n2738);
   U2663 : HS65_LH_FA1X4 port map( A0 => n1399, B0 => n817, CI => n270, CO => 
                           n269, S0 => product(20));
   U2664 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2699, Z => n1399);
   U2665 : HS65_LH_MX41X7 port map( D0 => n4493, S0 => n1019, D1 => n4591, S1 
                           => n4653, D2 => n4594, S2 => n4655, D3 => n4598, S3 
                           => n4656, Z => n2699);
   U2666 : HS65_LH_FA1X4 port map( A0 => n1135, B0 => n707, CI => n722, CO => 
                           n704, S0 => n705);
   U2667 : HS65_LHS_XOR2X6 port map( A => a(26), B => n3025, Z => n1135);
   U2668 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1035, D1 => n4507, S1 
                           => n4621, D2 => n4510, S2 => n4623, D3 => n4516, S3 
                           => n4624, Z => n3025);
   U2669 : HS65_LH_FA1X4 port map( A0 => n1168, B0 => n723, CI => n738, CO => 
                           n720, S0 => n721);
   U2670 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2984, Z => n1168);
   U2671 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1033, D1 => n4526, S1 
                           => n4628, D2 => n4518, S2 => n4625, D3 => n4521, S3 
                           => n4626, Z => n2984);
   U2672 : HS65_LH_FA1X4 port map( A0 => n1201, B0 => n739, CI => n752, CO => 
                           n736, S0 => n737);
   U2673 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2943, Z => n1201);
   U2674 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1031, D1 => n4528, S1 
                           => n4629, D2 => n4531, S2 => n4631, D3 => n4537, S3 
                           => n4632, Z => n2943);
   U2675 : HS65_LH_FA1X4 port map( A0 => n1234, B0 => n753, CI => n766, CO => 
                           n750, S0 => n751);
   U2676 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2902, Z => n1234);
   U2677 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1029, D1 => n4539, S1 
                           => n4633, D2 => n4543, S2 => n4635, D3 => n4548, S3 
                           => n4636, Z => n2902);
   U2678 : HS65_LH_FA1X4 port map( A0 => n1267, B0 => n767, CI => n780, CO => 
                           n764, S0 => n765);
   U2679 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2861, Z => n1267);
   U2680 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1027, D1 => n4551, S1 
                           => n4637, D2 => n4554, S2 => n4639, D3 => n4559, S3 
                           => n4640, Z => n2861);
   U2681 : HS65_LH_FA1X4 port map( A0 => n1300, B0 => n781, CI => n792, CO => 
                           n778, S0 => n779);
   U2682 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2820, Z => n1300);
   U2683 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1025, D1 => n4612, S1 
                           => n4644, D2 => n4565, S2 => n4643, D3 => n4562, S3 
                           => n4640, Z => n2820);
   U2684 : HS65_LH_FA1X4 port map( A0 => n1333, B0 => n793, CI => n804, CO => 
                           n790, S0 => n791);
   U2685 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2780, Z => n1333);
   U2686 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1023, D1 => n4570, S1 
                           => n4645, D2 => n4573, S2 => n4647, D3 => n4578, S3 
                           => n4648, Z => n2780);
   U2687 : HS65_LH_FA1X4 port map( A0 => n1366, B0 => n805, CI => n816, CO => 
                           n802, S0 => n803);
   U2688 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2739, Z => n1366);
   U2689 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1021, D1 => n4581, S1 
                           => n4649, D2 => n4584, S2 => n4651, D3 => n4589, S3 
                           => n4652, Z => n2739);
   U2690 : HS65_LH_FA1X4 port map( A0 => n1398, B0 => n803, CI => n269, CO => 
                           n268, S0 => product(21));
   U2691 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2700, Z => n1398);
   U2692 : HS65_LH_MX41X7 port map( D0 => n1018, S0 => n4494, D1 => n4591, S1 
                           => n4655, D2 => n4594, S2 => n4657, D3 => n4658, S3 
                           => n4599, Z => n2700);
   U2693 : HS65_LH_FA1X4 port map( A0 => n1101, B0 => n1069, CI => n688, CO => 
                           n670, S0 => n671);
   U2694 : HS65_LH_AO22X9 port map( A => n4606, B => n4617, C => n4490, D => 
                           n4617, Z => n1069);
   U2695 : HS65_LHS_XOR2X6 port map( A => a(29), B => n3067, Z => n1101);
   U2696 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1036, D1 => n4496, S1 
                           => n4618, D2 => n4500, S2 => n4621, D3 => n4505, S3 
                           => n4622, Z => n3067);
   U2697 : HS65_LH_FA1X4 port map( A0 => n1134, B0 => n689, CI => n704, CO => 
                           n686, S0 => n687);
   U2698 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3026, Z => n1134);
   U2699 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1034, D1 => n4506, S1 
                           => n4623, D2 => n4511, S2 => n4625, D3 => n4516, S3 
                           => n4626, Z => n3026);
   U2700 : HS65_LH_FA1X4 port map( A0 => n1167, B0 => n705, CI => n720, CO => 
                           n702, S0 => n703);
   U2701 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2985, Z => n1167);
   U2702 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1032, D1 => n4526, S1 
                           => n4631, D2 => n4518, S2 => n4627, D3 => n4521, S3 
                           => n4628, Z => n2985);
   U2703 : HS65_LH_FA1X4 port map( A0 => n1200, B0 => n721, CI => n736, CO => 
                           n718, S0 => n719);
   U2704 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2944, Z => n1200);
   U2705 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1030, D1 => n4528, S1 
                           => n4630, D2 => n4531, S2 => n4633, D3 => n4537, S3 
                           => n4634, Z => n2944);
   U2706 : HS65_LH_FA1X4 port map( A0 => n1233, B0 => n737, CI => n750, CO => 
                           n734, S0 => n735);
   U2707 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2903, Z => n1233);
   U2708 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1028, D1 => n4539, S1 
                           => n4635, D2 => n4542, S2 => n4637, D3 => n4548, S3 
                           => n4638, Z => n2903);
   U2709 : HS65_LH_FA1X4 port map( A0 => n1266, B0 => n751, CI => n764, CO => 
                           n748, S0 => n749);
   U2710 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2862, Z => n1266);
   U2711 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1026, D1 => n4551, S1 
                           => n4639, D2 => n4554, S2 => n4641, D3 => n4559, S3 
                           => n4642, Z => n2862);
   U2712 : HS65_LH_FA1X4 port map( A0 => n1299, B0 => n765, CI => n778, CO => 
                           n762, S0 => n763);
   U2713 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2821, Z => n1299);
   U2714 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1024, D1 => n4566, S1 
                           => n4645, D2 => n4611, S2 => n4647, D3 => n4561, S3 
                           => n4642, Z => n2821);
   U2715 : HS65_LH_FA1X4 port map( A0 => n1332, B0 => n779, CI => n790, CO => 
                           n776, S0 => n777);
   U2716 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2781, Z => n1332);
   U2717 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1022, D1 => n4570, S1 
                           => n4647, D2 => n4573, S2 => n4649, D3 => n4578, S3 
                           => n4650, Z => n2781);
   U2718 : HS65_LH_FA1X4 port map( A0 => n1365, B0 => n791, CI => n802, CO => 
                           n788, S0 => n789);
   U2719 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2740, Z => n1365);
   U2720 : HS65_LH_MX41X7 port map( D0 => n2719, S0 => n1020, D1 => n4581, S1 
                           => n4651, D2 => n4584, S2 => n4653, D3 => n4589, S3 
                           => n4654, Z => n2740);
   U2721 : HS65_LH_FA1X4 port map( A0 => n1397, B0 => n789, CI => n268, CO => 
                           n267, S0 => product(22));
   U2722 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2701, Z => n1397);
   U2723 : HS65_LH_MX41X7 port map( D0 => n1017, S0 => n4494, D1 => n4591, S1 
                           => n4656, D2 => n4658, S2 => n4596, D3 => n4660, S3 
                           => n4600, Z => n2701);
   U2724 : HS65_LH_FA1X4 port map( A0 => n1100, B0 => n1068, CI => n670, CO => 
                           n652, S0 => n653);
   U2725 : HS65_LH_AO222X4 port map( A => n4608, B => n4619, C => n4602, D => 
                           n4617, E => n4490, F => n1038, Z => n1068);
   U2726 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3068, Z => n1100);
   U2727 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1035, D1 => n4496, S1 
                           => n4620, D2 => n4499, S2 => n4623, D3 => n4505, S3 
                           => n4624, Z => n3068);
   U2728 : HS65_LH_FA1X4 port map( A0 => n1133, B0 => n671, CI => n686, CO => 
                           n668, S0 => n669);
   U2729 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3027, Z => n1133);
   U2730 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1033, D1 => n4507, S1 
                           => n4625, D2 => n4510, S2 => n4627, D3 => n4515, S3 
                           => n4628, Z => n3027);
   U2731 : HS65_LH_FA1X4 port map( A0 => n1166, B0 => n687, CI => n702, CO => 
                           n684, S0 => n685);
   U2732 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2986, Z => n1166);
   U2733 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1031, D1 => n4526, S1 
                           => n4633, D2 => n4517, S2 => n4629, D3 => n4521, S3 
                           => n4630, Z => n2986);
   U2734 : HS65_LH_FA1X4 port map( A0 => n1199, B0 => n703, CI => n718, CO => 
                           n700, S0 => n701);
   U2735 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2945, Z => n1199);
   U2736 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1029, D1 => n4528, S1 
                           => n4632, D2 => n4531, S2 => n4635, D3 => n4536, S3 
                           => n4636, Z => n2945);
   U2737 : HS65_LH_FA1X4 port map( A0 => n1232, B0 => n719, CI => n734, CO => 
                           n716, S0 => n717);
   U2738 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2904, Z => n1232);
   U2739 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1027, D1 => n4540, S1 
                           => n4637, D2 => n4543, S2 => n4639, D3 => n4549, S3 
                           => n4640, Z => n2904);
   U2740 : HS65_LH_FA1X4 port map( A0 => n1265, B0 => n735, CI => n748, CO => 
                           n732, S0 => n733);
   U2741 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2863, Z => n1265);
   U2742 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1025, D1 => n4551, S1 
                           => n4641, D2 => n4554, S2 => n4643, D3 => n4559, S3 
                           => n4644, Z => n2863);
   U2743 : HS65_LH_FA1X4 port map( A0 => n1298, B0 => n749, CI => n762, CO => 
                           n746, S0 => n747);
   U2744 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2822, Z => n1298);
   U2745 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1023, D1 => n4566, S1 
                           => n4646, D2 => n4611, S2 => n4649, D3 => n4561, S3 
                           => n4644, Z => n2822);
   U2746 : HS65_LH_FA1X4 port map( A0 => n1331, B0 => n763, CI => n776, CO => 
                           n760, S0 => n761);
   U2747 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2782, Z => n1331);
   U2748 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1021, D1 => n4570, S1 
                           => n4649, D2 => n4573, S2 => n4651, D3 => n4578, S3 
                           => n4652, Z => n2782);
   U2749 : HS65_LH_FA1X4 port map( A0 => n1364, B0 => n777, CI => n788, CO => 
                           n774, S0 => n775);
   U2750 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2741, Z => n1364);
   U2751 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1019, D1 => n4581, S1 
                           => n4652, D2 => n4584, S2 => n4655, D3 => n4589, S3 
                           => n4656, Z => n2741);
   U2752 : HS65_LH_FA1X4 port map( A0 => n1396, B0 => n775, CI => n267, CO => 
                           n266, S0 => product(23));
   U2753 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2702, Z => n1396);
   U2754 : HS65_LH_MX41X7 port map( D0 => n1016, S0 => n4494, D1 => n4658, S1 
                           => n4592, D2 => n4660, S2 => n4596, D3 => n4662, S3 
                           => n4600, Z => n2702);
   U2755 : HS65_LH_FA1X4 port map( A0 => n1099, B0 => n1067, CI => n652, CO => 
                           n634, S0 => n635);
   U2756 : HS65_LH_MX41X7 port map( D0 => n1037, S0 => n4492, D1 => n4620, S1 
                           => n4608, D2 => n4618, S2 => n4604, D3 => n4616, S3 
                           => n4609, Z => n1067);
   U2757 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3069, Z => n1099);
   U2758 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1034, D1 => n4496, S1 
                           => n4622, D2 => n4499, S2 => n4625, D3 => n4505, S3 
                           => n4626, Z => n3069);
   U2759 : HS65_LH_FA1X4 port map( A0 => n1132, B0 => n653, CI => n668, CO => 
                           n650, S0 => n651);
   U2760 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3028, Z => n1132);
   U2761 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1032, D1 => n4507, S1 
                           => n4626, D2 => n4510, S2 => n4629, D3 => n4515, S3 
                           => n4630, Z => n3028);
   U2762 : HS65_LH_FA1X4 port map( A0 => n1165, B0 => n669, CI => n684, CO => 
                           n666, S0 => n667);
   U2763 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2987, Z => n1165);
   U2764 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1030, D1 => n4526, S1 
                           => n4634, D2 => n4517, S2 => n4631, D3 => n4521, S3 
                           => n4632, Z => n2987);
   U2765 : HS65_LH_FA1X4 port map( A0 => n1198, B0 => n685, CI => n700, CO => 
                           n682, S0 => n683);
   U2766 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2946, Z => n1198);
   U2767 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1028, D1 => n4528, S1 
                           => n4634, D2 => n4531, S2 => n4637, D3 => n4536, S3 
                           => n4638, Z => n2946);
   U2768 : HS65_LH_FA1X4 port map( A0 => n1231, B0 => n701, CI => n716, CO => 
                           n698, S0 => n699);
   U2769 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2905, Z => n1231);
   U2770 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1026, D1 => n4540, S1 
                           => n4638, D2 => n4543, S2 => n4641, D3 => n4548, S3 
                           => n4642, Z => n2905);
   U2771 : HS65_LH_FA1X4 port map( A0 => n1264, B0 => n717, CI => n732, CO => 
                           n714, S0 => n715);
   U2772 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2864, Z => n1264);
   U2773 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1024, D1 => n4550, S1 
                           => n4643, D2 => n4553, S2 => n4645, D3 => n4558, S3 
                           => n4646, Z => n2864);
   U2774 : HS65_LH_FA1X4 port map( A0 => n1297, B0 => n733, CI => n746, CO => 
                           n730, S0 => n731);
   U2775 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2823, Z => n1297);
   U2776 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1022, D1 => n4611, S1 
                           => n4651, D2 => n4564, S2 => n4649, D3 => n4561, S3 
                           => n4646, Z => n2823);
   U2777 : HS65_LH_FA1X4 port map( A0 => n1330, B0 => n747, CI => n760, CO => 
                           n744, S0 => n745);
   U2778 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2783, Z => n1330);
   U2779 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1020, D1 => n4570, S1 
                           => n4651, D2 => n4573, S2 => n4653, D3 => n4578, S3 
                           => n4654, Z => n2783);
   U2780 : HS65_LH_FA1X4 port map( A0 => n1363, B0 => n761, CI => n774, CO => 
                           n758, S0 => n759);
   U2781 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2742, Z => n1363);
   U2782 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1018, D1 => n4580, S1 
                           => n4654, D2 => n4583, S2 => n4657, D3 => n4588, S3 
                           => n4658, Z => n2742);
   U2783 : HS65_LH_FA1X4 port map( A0 => n1395, B0 => n759, CI => n266, CO => 
                           n265, S0 => product(24));
   U2784 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2703, Z => n1395);
   U2785 : HS65_LH_MX41X7 port map( D0 => n1015, S0 => n4494, D1 => n4660, S1 
                           => n4592, D2 => n4662, S2 => n4596, D3 => n4598, S3 
                           => n4664, Z => n2703);
   U2786 : HS65_LH_FA1X4 port map( A0 => n1131, B0 => n635, CI => n650, CO => 
                           n632, S0 => n633);
   U2787 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3029, Z => n1131);
   U2788 : HS65_LH_MX41X7 port map( D0 => n3019, S0 => n1031, D1 => n4507, S1 
                           => n4629, D2 => n4510, S2 => n4631, D3 => n4515, S3 
                           => n4632, Z => n3029);
   U2789 : HS65_LH_FA1X4 port map( A0 => n1164, B0 => n651, CI => n666, CO => 
                           n648, S0 => n649);
   U2790 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2988, Z => n1164);
   U2791 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1029, D1 => n4526, S1 
                           => n4636, D2 => n4517, S2 => n4633, D3 => n4520, S3 
                           => n4634, Z => n2988);
   U2792 : HS65_LH_FA1X4 port map( A0 => n1197, B0 => n667, CI => n682, CO => 
                           n664, S0 => n665);
   U2793 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2947, Z => n1197);
   U2794 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1027, D1 => n4529, S1 
                           => n4636, D2 => n4532, S2 => n4639, D3 => n4537, S3 
                           => n4640, Z => n2947);
   U2795 : HS65_LH_FA1X4 port map( A0 => n1230, B0 => n683, CI => n698, CO => 
                           n680, S0 => n681);
   U2796 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2906, Z => n1230);
   U2797 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1025, D1 => n4540, S1 
                           => n4641, D2 => n4543, S2 => n4643, D3 => n4548, S3 
                           => n4644, Z => n2906);
   U2798 : HS65_LH_FA1X4 port map( A0 => n1263, B0 => n699, CI => n714, CO => 
                           n696, S0 => n697);
   U2799 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2865, Z => n1263);
   U2800 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1023, D1 => n4551, S1 
                           => n4645, D2 => n4554, S2 => n4647, D3 => n4559, S3 
                           => n4648, Z => n2865);
   U2801 : HS65_LH_FA1X4 port map( A0 => n1296, B0 => n715, CI => n730, CO => 
                           n712, S0 => n713);
   U2802 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2824, Z => n1296);
   U2803 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1021, D1 => n4612, S1 
                           => n4653, D2 => n4565, S2 => n4651, D3 => n4562, S3 
                           => n4648, Z => n2824);
   U2804 : HS65_LH_FA1X4 port map( A0 => n1329, B0 => n731, CI => n744, CO => 
                           n728, S0 => n729);
   U2805 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2784, Z => n1329);
   U2806 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1019, D1 => n4570, S1 
                           => n4652, D2 => n4573, S2 => n4655, D3 => n4578, S3 
                           => n4656, Z => n2784);
   U2807 : HS65_LH_FA1X4 port map( A0 => n1362, B0 => n745, CI => n758, CO => 
                           n742, S0 => n743);
   U2808 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2743, Z => n1362);
   U2809 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1017, D1 => n4581, S1 
                           => n4656, D2 => n4584, S2 => n4659, D3 => n4589, S3 
                           => n4660, Z => n2743);
   U2810 : HS65_LH_FA1X4 port map( A0 => n1394, B0 => n743, CI => n265, CO => 
                           n264, S0 => product(25));
   U2811 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2704, Z => n1394);
   U2812 : HS65_LH_MX41X7 port map( D0 => n1014, S0 => n4494, D1 => n4662, S1 
                           => n4592, D2 => n4594, S2 => n4665, D3 => n4598, S3 
                           => n4666, Z => n2704);
   U2813 : HS65_LH_FA1X4 port map( A0 => n1163, B0 => n633, CI => n648, CO => 
                           n630, S0 => n631);
   U2814 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2989, Z => n1163);
   U2815 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1028, D1 => n4526, S1 
                           => n4639, D2 => n4518, S2 => n4635, D3 => n4521, S3 
                           => n4636, Z => n2989);
   U2816 : HS65_LH_FA1X4 port map( A0 => n1196, B0 => n649, CI => n664, CO => 
                           n646, S0 => n647);
   U2817 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2948, Z => n1196);
   U2818 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1026, D1 => n4529, S1 
                           => n4639, D2 => n4532, S2 => n4641, D3 => n4537, S3 
                           => n4642, Z => n2948);
   U2819 : HS65_LH_FA1X4 port map( A0 => n1229, B0 => n665, CI => n680, CO => 
                           n662, S0 => n663);
   U2820 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2907, Z => n1229);
   U2821 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1024, D1 => n4539, S1 
                           => n4643, D2 => n4542, S2 => n4645, D3 => n4547, S3 
                           => n4646, Z => n2907);
   U2822 : HS65_LH_FA1X4 port map( A0 => n1262, B0 => n681, CI => n696, CO => 
                           n678, S0 => n679);
   U2823 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2866, Z => n1262);
   U2824 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1022, D1 => n4551, S1 
                           => n4647, D2 => n4554, S2 => n4649, D3 => n4559, S3 
                           => n4650, Z => n2866);
   U2825 : HS65_LH_FA1X4 port map( A0 => n1295, B0 => n697, CI => n712, CO => 
                           n694, S0 => n695);
   U2826 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2825, Z => n1295);
   U2827 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1020, D1 => n4612, S1 
                           => n4654, D2 => n4565, S2 => n4653, D3 => n4562, S3 
                           => n4650, Z => n2825);
   U2828 : HS65_LH_FA1X4 port map( A0 => n1328, B0 => n713, CI => n728, CO => 
                           n710, S0 => n711);
   U2829 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2785, Z => n1328);
   U2830 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1018, D1 => n4569, S1 
                           => n4655, D2 => n4572, S2 => n4657, D3 => n4577, S3 
                           => n4658, Z => n2785);
   U2831 : HS65_LH_FA1X4 port map( A0 => n1361, B0 => n729, CI => n742, CO => 
                           n726, S0 => n727);
   U2832 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2744, Z => n1361);
   U2833 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1016, D1 => n4581, S1 
                           => n4659, D2 => n4584, S2 => n4661, D3 => n4589, S3 
                           => n4662, Z => n2744);
   U2834 : HS65_LH_FA1X4 port map( A0 => n1393, B0 => n727, CI => n264, CO => 
                           n263, S0 => product(26));
   U2835 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2705, Z => n1393);
   U2836 : HS65_LH_MX41X7 port map( D0 => n4493, S0 => n1013, D1 => n4591, S1 
                           => n4665, D2 => n4594, S2 => n4667, D3 => n4598, S3 
                           => n4668, Z => n2705);
   U2837 : HS65_LH_FA1X4 port map( A0 => n1195, B0 => n631, CI => n646, CO => 
                           n628, S0 => n629);
   U2838 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2949, Z => n1195);
   U2839 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1025, D1 => n4529, S1 
                           => n4640, D2 => n4532, S2 => n4643, D3 => n4537, S3 
                           => n4644, Z => n2949);
   U2840 : HS65_LH_FA1X4 port map( A0 => n1228, B0 => n647, CI => n662, CO => 
                           n644, S0 => n645);
   U2841 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2908, Z => n1228);
   U2842 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1023, D1 => n4540, S1 
                           => n4645, D2 => n4543, S2 => n4647, D3 => n4548, S3 
                           => n4648, Z => n2908);
   U2843 : HS65_LH_FA1X4 port map( A0 => n1261, B0 => n663, CI => n678, CO => 
                           n660, S0 => n661);
   U2844 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2867, Z => n1261);
   U2845 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1021, D1 => n4551, S1 
                           => n4649, D2 => n4554, S2 => n4651, D3 => n4559, S3 
                           => n4652, Z => n2867);
   U2846 : HS65_LH_FA1X4 port map( A0 => n1294, B0 => n679, CI => n694, CO => 
                           n676, S0 => n677);
   U2847 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2826, Z => n1294);
   U2848 : HS65_LH_MX41X7 port map( D0 => n2804, S0 => n1019, D1 => n4612, S1 
                           => n4657, D2 => n4565, S2 => n4655, D3 => n4562, S3 
                           => n4652, Z => n2826);
   U2849 : HS65_LH_FA1X4 port map( A0 => n1327, B0 => n695, CI => n710, CO => 
                           n692, S0 => n693);
   U2850 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2786, Z => n1327);
   U2851 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1017, D1 => n4569, S1 
                           => n4657, D2 => n4573, S2 => n4659, D3 => n4578, S3 
                           => n4660, Z => n2786);
   U2852 : HS65_LH_FA1X4 port map( A0 => n1360, B0 => n711, CI => n726, CO => 
                           n708, S0 => n709);
   U2853 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2745, Z => n1360);
   U2854 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1015, D1 => n4580, S1 
                           => n4661, D2 => n4583, S2 => n4663, D3 => n4588, S3 
                           => n4664, Z => n2745);
   U2855 : HS65_LH_FA1X4 port map( A0 => n1392, B0 => n709, CI => n263, CO => 
                           n262, S0 => product(27));
   U2856 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2706, Z => n1392);
   U2857 : HS65_LH_MX41X7 port map( D0 => n1012, S0 => n4494, D1 => n4591, S1 
                           => n4667, D2 => n4594, S2 => n4669, D3 => n4670, S3 
                           => n4600, Z => n2706);
   U2858 : HS65_LH_FA1X4 port map( A0 => n1227, B0 => n629, CI => n644, CO => 
                           n626, S0 => n627);
   U2859 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2909, Z => n1227);
   U2860 : HS65_LH_MX41X7 port map( D0 => n2890, S0 => n1022, D1 => n4540, S1 
                           => n4646, D2 => n4543, S2 => n4649, D3 => n4548, S3 
                           => n4650, Z => n2909);
   U2861 : HS65_LH_FA1X4 port map( A0 => n1260, B0 => n645, CI => n660, CO => 
                           n642, S0 => n643);
   U2862 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2868, Z => n1260);
   U2863 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1020, D1 => n4551, S1 
                           => n4651, D2 => n4554, S2 => n4653, D3 => n4559, S3 
                           => n4654, Z => n2868);
   U2864 : HS65_LH_FA1X4 port map( A0 => n1293, B0 => n661, CI => n676, CO => 
                           n658, S0 => n659);
   U2865 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2827, Z => n1293);
   U2866 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1018, D1 => n4612, S1 
                           => n4658, D2 => n4565, S2 => n4657, D3 => n4562, S3 
                           => n4654, Z => n2827);
   U2867 : HS65_LH_FA1X4 port map( A0 => n1326, B0 => n677, CI => n692, CO => 
                           n674, S0 => n675);
   U2868 : HS65_LHS_XOR2X6 port map( A => n4686, B => n2787, Z => n1326);
   U2869 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1016, D1 => n4569, S1 
                           => n4659, D2 => n4572, S2 => n4661, D3 => n4578, S3 
                           => n4662, Z => n2787);
   U2870 : HS65_LH_FA1X4 port map( A0 => n1359, B0 => n693, CI => n708, CO => 
                           n690, S0 => n691);
   U2871 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2746, Z => n1359);
   U2872 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1014, D1 => n4580, S1 
                           => n4662, D2 => n4583, S2 => n4665, D3 => n4588, S3 
                           => n4666, Z => n2746);
   U2873 : HS65_LH_FA1X4 port map( A0 => n1391, B0 => n691, CI => n262, CO => 
                           n261, S0 => product(28));
   U2874 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2707, Z => n1391);
   U2875 : HS65_LH_MX41X7 port map( D0 => n1011, S0 => n4494, D1 => n4591, S1 
                           => n4669, D2 => n4670, S2 => n4595, D3 => n4672, S3 
                           => n4599, Z => n2707);
   U2876 : HS65_LH_FA1X4 port map( A0 => n1259, B0 => n627, CI => n642, CO => 
                           n624, S0 => n625);
   U2877 : HS65_LHS_XOR2X6 port map( A => n4692, B => n2869, Z => n1259);
   U2878 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1019, D1 => n4551, S1 
                           => n4652, D2 => n4554, S2 => n4655, D3 => n4559, S3 
                           => n4656, Z => n2869);
   U2879 : HS65_LH_FA1X4 port map( A0 => n1292, B0 => n643, CI => n658, CO => 
                           n640, S0 => n641);
   U2880 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2828, Z => n1292);
   U2881 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1017, D1 => n4612, S1 
                           => n4660, D2 => n4565, S2 => n4659, D3 => n4562, S3 
                           => n4656, Z => n2828);
   U2882 : HS65_LH_FA1X4 port map( A0 => n1325, B0 => n659, CI => n674, CO => 
                           n656, S0 => n657);
   U2883 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2788, Z => n1325);
   U2884 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1015, D1 => n4569, S1 
                           => n4661, D2 => n4572, S2 => n4663, D3 => n4577, S3 
                           => n4664, Z => n2788);
   U2885 : HS65_LH_FA1X4 port map( A0 => n1358, B0 => n675, CI => n690, CO => 
                           n672, S0 => n673);
   U2886 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2747, Z => n1358);
   U2887 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1013, D1 => n4580, S1 
                           => n4664, D2 => n4584, S2 => n4667, D3 => n4589, S3 
                           => n4668, Z => n2747);
   U2888 : HS65_LH_FA1X4 port map( A0 => n1390, B0 => n673, CI => n261, CO => 
                           n260, S0 => product(29));
   U2889 : HS65_LHS_XOR2X6 port map( A => a(2), B => n2708, Z => n1390);
   U2890 : HS65_LH_MX41X7 port map( D0 => n1010, S0 => n4494, D1 => n4670, S1 
                           => n4592, D2 => n4672, S2 => n4595, D3 => n4674, S3 
                           => n4600, Z => n2708);
   U2891 : HS65_LH_FA1X4 port map( A0 => n1291, B0 => n625, CI => n640, CO => 
                           n622, S0 => n623);
   U2892 : HS65_LHS_XOR2X6 port map( A => n4689, B => n2829, Z => n1291);
   U2893 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1016, D1 => n4612, S1 
                           => n4663, D2 => n4564, S2 => n4661, D3 => n4562, S3 
                           => n4658, Z => n2829);
   U2894 : HS65_LH_FA1X4 port map( A0 => n1324, B0 => n641, CI => n656, CO => 
                           n638, S0 => n639);
   U2895 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2789, Z => n1324);
   U2896 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1014, D1 => n4569, S1 
                           => n4662, D2 => n4572, S2 => n4665, D3 => n4577, S3 
                           => n4666, Z => n2789);
   U2897 : HS65_LH_FA1X4 port map( A0 => n1357, B0 => n657, CI => n672, CO => 
                           n654, S0 => n655);
   U2898 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2748, Z => n1357);
   U2899 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1012, D1 => n4580, S1 
                           => n4667, D2 => n4584, S2 => n4669, D3 => n4589, S3 
                           => n4670, Z => n2748);
   U2900 : HS65_LH_FA1X4 port map( A0 => n1389, B0 => n655, CI => n260, CO => 
                           n259, S0 => product(30));
   U2901 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2709, Z => n1389);
   U2902 : HS65_LH_MX41X7 port map( D0 => n1009, S0 => n4494, D1 => n4672, S1 
                           => n4592, D2 => n4674, S2 => n4595, D3 => n4676, S3 
                           => n4599, Z => n2709);
   U2903 : HS65_LH_FA1X4 port map( A0 => n1323, B0 => n623, CI => n638, CO => 
                           n620, S0 => n621);
   U2904 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2790, Z => n1323);
   U2905 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1013, D1 => n4569, S1 
                           => n4664, D2 => n4573, S2 => n4667, D3 => n4578, S3 
                           => n4668, Z => n2790);
   U2906 : HS65_LH_FA1X4 port map( A0 => n1356, B0 => n639, CI => n654, CO => 
                           n636, S0 => n637);
   U2907 : HS65_LHS_XOR2X6 port map( A => n4683, B => n2749, Z => n1356);
   U2908 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1011, D1 => n4580, S1 
                           => n4669, D2 => n4583, S2 => n4671, D3 => n4589, S3 
                           => n4672, Z => n2749);
   U2909 : HS65_LH_FA1X4 port map( A0 => n1388, B0 => n637, CI => n259, CO => 
                           n258, S0 => product(31));
   U2910 : HS65_LHS_XOR2X6 port map( A => n4680, B => n2710, Z => n1388);
   U2911 : HS65_LH_MX41X7 port map( D0 => n1008, S0 => n4493, D1 => n4674, S1 
                           => n4591, D2 => n4676, S2 => n4594, D3 => n4598, S3 
                           => n4678, Z => n2710);
   U2912 : HS65_LH_FA1X4 port map( A0 => n1355, B0 => n621, CI => n636, CO => 
                           n618, S0 => n619);
   U2913 : HS65_LHS_XOR2X6 port map( A => a(5), B => n2750, Z => n1355);
   U2914 : HS65_LH_MX41X7 port map( D0 => n4586, S0 => n1010, D1 => n4580, S1 
                           => n4671, D2 => n4583, S2 => n4673, D3 => n4588, S3 
                           => n4674, Z => n2750);
   U2915 : HS65_LH_FA1X4 port map( A0 => n1204, B0 => n787, CI => n798, CO => 
                           n784, S0 => n785);
   U2916 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2940, Z => n1204);
   U2917 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1034, D1 => n4528, S1 
                           => n4623, D2 => n4533, S2 => n4625, D3 => n4538, S3 
                           => n4626, Z => n2940);
   U2918 : HS65_LH_FA1X4 port map( A0 => n599, B0 => n616, CI => n1129, CO => 
                           n596, S0 => n597);
   U2919 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3031, Z => n1129);
   U2920 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1029, D1 => n4506, S1 
                           => n4632, D2 => n4510, S2 => n4635, D3 => n4515, S3 
                           => n4636, Z => n3031);
   U2921 : HS65_LH_FA1X4 port map( A0 => n477, B0 => n491, CI => n1122, CO => 
                           n474, S0 => n475);
   U2922 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3038, Z => n1122);
   U2923 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1022, D1 => n4506, S1 
                           => n4647, D2 => n4509, S2 => n4649, D3 => n4514, S3 
                           => n4650, Z => n3038);
   U2924 : HS65_LH_FA1X4 port map( A0 => n473, B0 => n487, CI => n1186, CO => 
                           n470, S0 => n471);
   U2925 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2958, Z => n1186);
   U2926 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1016, D1 => n4528, S1 
                           => n4659, D2 => n4531, S2 => n4661, D3 => n4536, S3 
                           => n4662, Z => n2958);
   U2927 : HS65_LH_FA1X4 port map( A0 => n581, B0 => n1096, CI => n596, CO => 
                           n578, S0 => n579);
   U2928 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3072, Z => n1096);
   U2929 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1031, D1 => n4496, S1 
                           => n4629, D2 => n4499, S2 => n4631, D3 => n4504, S3 
                           => n4632, Z => n3072);
   U2930 : HS65_LH_FA1X4 port map( A0 => n595, B0 => n612, CI => n1193, CO => 
                           n592, S0 => n593);
   U2931 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2951, Z => n1193);
   U2932 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1023, D1 => n4528, S1 
                           => n4644, D2 => n4531, S2 => n4647, D3 => n4536, S3 
                           => n4648, Z => n2951);
   U2933 : HS65_LH_FA1X4 port map( A0 => n563, B0 => n1095, CI => n578, CO => 
                           n560, S0 => n561);
   U2934 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3073, Z => n1095);
   U2935 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1030, D1 => n4496, S1 
                           => n4630, D2 => n4499, S2 => n4633, D3 => n4504, S3 
                           => n4634, Z => n3073);
   U2936 : HS65_LH_FA1X4 port map( A0 => n561, B0 => n1127, CI => n1159, CO => 
                           n558, S0 => n559);
   U2937 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2993, Z => n1159);
   U2938 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3033, Z => n1127);
   U2939 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1024, D1 => n4525, S1 
                           => n4647, D2 => n4517, S2 => n4643, D3 => n4520, S3 
                           => n4644, Z => n2993);
   U2940 : HS65_LH_FA1X4 port map( A0 => n591, B0 => n608, CI => n1257, CO => 
                           n588, S0 => n589);
   U2941 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2871, Z => n1257);
   U2942 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1017, D1 => n4550, S1 
                           => n4656, D2 => n4553, S2 => n4659, D3 => n4558, S3 
                           => n4660, Z => n2871);
   U2943 : HS65_LH_FA1X4 port map( A0 => n589, B0 => n606, CI => n1289, CO => 
                           n586, S0 => n587);
   U2944 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2831, Z => n1289);
   U2945 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1014, D1 => n4611, S1 
                           => n4666, D2 => n4564, S2 => n4665, D3 => n4561, S3 
                           => n4662, Z => n2831);
   U2946 : HS65_LH_FA1X4 port map( A0 => n587, B0 => n604, CI => n1321, CO => 
                           n584, S0 => n585);
   U2947 : HS65_LHS_XOR2X6 port map( A => n4685, B => n2792, Z => n1321);
   U2948 : HS65_LH_MX41X7 port map( D0 => n4575, S0 => n1011, D1 => n4569, S1 
                           => n4668, D2 => n4572, S2 => n4671, D3 => n4577, S3 
                           => n4672, Z => n2792);
   U2949 : HS65_LH_FA1X4 port map( A0 => n551, B0 => n1287, CI => n566, CO => 
                           n548, S0 => n549);
   U2950 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2833, Z => n1287);
   U2951 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1012, D1 => n4611, S1 
                           => n4670, D2 => n4564, S2 => n4669, D3 => n4561, S3 
                           => n4666, Z => n2833);
   U2952 : HS65_LH_FA1X4 port map( A0 => n521, B0 => n537, CI => n1221, CO => 
                           n518, S0 => n519);
   U2953 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2915, Z => n1221);
   U2954 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1016, D1 => n4539, S1 
                           => n4659, D2 => n4542, S2 => n4661, D3 => n4547, S3 
                           => n4662, Z => n2915);
   U2955 : HS65_LH_FA1X4 port map( A0 => n517, B0 => n533, CI => n1285, CO => 
                           n514, S0 => n515);
   U2956 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2835, Z => n1285);
   U2957 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1010, D1 => n4611, S1 
                           => n4674, D2 => n4564, S2 => n4673, D3 => n4561, S3 
                           => n4670, Z => n2835);
   U2958 : HS65_LH_FA1X4 port map( A0 => n469, B0 => n483, CI => n1250, CO => 
                           n466, S0 => n467);
   U2959 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2878, Z => n1250);
   U2960 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1010, D1 => n4550, S1 
                           => n4671, D2 => n4554, S2 => n4673, D3 => n4559, S3 
                           => n4674, Z => n2878);
   U2961 : HS65_LH_FA1X4 port map( A0 => n430, B0 => n442, CI => n1151, CO => 
                           n427, S0 => n428);
   U2962 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3001, Z => n1151);
   U2963 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1016, D1 => n4525, S1 
                           => n4663, D2 => n4517, S2 => n4659, D3 => n4520, S3 
                           => n4660, Z => n3001);
   U2964 : HS65_LH_FA1X4 port map( A0 => n426, B0 => n438, CI => n1215, CO => 
                           n423, S0 => n424);
   U2965 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2921, Z => n1215);
   U2966 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1010, D1 => n4539, S1 
                           => n4670, D2 => n4542, S2 => n4673, D3 => n4547, S3 
                           => n4674, Z => n2921);
   U2967 : HS65_LH_FA1X4 port map( A0 => n394, B0 => n404, CI => n1116, CO => 
                           n391, S0 => n392);
   U2968 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3044, Z => n1116);
   U2969 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1016, D1 => n4506, S1 
                           => n4658, D2 => n4509, S2 => n4661, D3 => n4514, S3 
                           => n4662, Z => n3044);
   U2970 : HS65_LH_FA1X4 port map( A0 => n390, B0 => n400, CI => n1180, CO => 
                           n387, S0 => n388);
   U2971 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2964, Z => n1180);
   U2972 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1010, D1 => n4529, S1 
                           => n4671, D2 => n4532, S2 => n4673, D3 => n4537, S3 
                           => n4674, Z => n2964);
   U2973 : HS65_LH_FA1X4 port map( A0 => n359, B0 => n367, CI => n1145, CO => 
                           n356, S0 => n357);
   U2974 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3007, Z => n1145);
   U2975 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1010, D1 => n4525, S1 
                           => n4675, D2 => n4517, S2 => n4671, D3 => n4520, S3 
                           => n4672, Z => n3007);
   U2976 : HS65_LH_FA1X4 port map( A0 => n335, B0 => n341, CI => n1110, CO => 
                           n332, S0 => n333);
   U2977 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3050, Z => n1110);
   U2978 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1010, D1 => n4506, S1 
                           => n4671, D2 => n4509, S2 => n4673, D3 => n4514, S3 
                           => n4674, Z => n3050);
   U2979 : HS65_LH_FA1X4 port map( A0 => n571, B0 => n1256, CI => n586, CO => 
                           n568, S0 => n569);
   U2980 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2872, Z => n1256);
   U2981 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1016, D1 => n4550, S1 
                           => n4659, D2 => n4553, S2 => n4661, D3 => n4558, S3 
                           => n4662, Z => n2872);
   U2982 : HS65_LH_FA1X4 port map( A0 => n525, B0 => n541, CI => n1157, CO => 
                           n522, S0 => n523);
   U2983 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2995, Z => n1157);
   U2984 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1022, D1 => n4525, S1 
                           => n4650, D2 => n4517, S2 => n4647, D3 => n4520, S3 
                           => n4648, Z => n2995);
   U2985 : HS65_LH_FA1X4 port map( A0 => n601, B0 => n1386, CI => n257, CO => 
                           n256, S0 => product(33));
   U2986 : HS65_LHS_XOR2X6 port map( A => n4682, B => n2716, Z => n1386);
   U2987 : HS65_LH_AOI22X6 port map( A => n4493, B => n1006, C => n4591, D => 
                           n4678, Z => n2716);
   U2988 : HS65_LH_FA1X4 port map( A0 => n569, B0 => n1288, CI => n584, CO => 
                           n566, S0 => n567);
   U2989 : HS65_LHS_XOR2X6 port map( A => n4688, B => n2832, Z => n1288);
   U2990 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1013, D1 => n4612, S1 
                           => n4668, D2 => n4565, S2 => n4667, D3 => n4561, S3 
                           => n4664, Z => n2832);
   U2991 : HS65_LH_FA1X4 port map( A0 => n4709, B0 => n1061, CI => n1093, CO =>
                           n526, S0 => n527);
   U2992 : HS65_LH_MX41X7 port map( D0 => n1031, S0 => n4490, D1 => n4632, S1 
                           => n4607, D2 => n4630, S2 => n4602, D3 => n4628, S3 
                           => n4609, Z => n1061);
   U2993 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3075, Z => n1093);
   U2994 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1028, D1 => n4495, S1 
                           => n4635, D2 => n4498, S2 => n4637, D3 => n4503, S3 
                           => n4638, Z => n3075);
   U2995 : HS65_LH_FA1X4 port map( A0 => n4713, B0 => n446, CI => n1087, CO => 
                           n431, S0 => n432);
   U2996 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3081, Z => n1087);
   U2997 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1022, D1 => n4495, S1 
                           => n4647, D2 => n4498, S2 => n4649, D3 => n4503, S3 
                           => n4650, Z => n3081);
   U2998 : HS65_LH_FA1X4 port map( A0 => n4714, B0 => n371, CI => n1081, CO => 
                           n360, S0 => n361);
   U2999 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3087, Z => n1081);
   U3000 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1016, D1 => n4495, S1 
                           => n4659, D2 => n4498, S2 => n4661, D3 => n4503, S3 
                           => n4662, Z => n3087);
   U3001 : HS65_LH_FA1X4 port map( A0 => n4715, B0 => n320, CI => n1075, CO => 
                           n313, S0 => n314);
   U3002 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3093, Z => n1075);
   U3003 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1010, D1 => n4495, S1 
                           => n4671, D2 => n4498, S2 => n4673, D3 => n4504, S3 
                           => n4674, Z => n3093);
   U3004 : HS65_LH_FA1X4 port map( A0 => n1065, B0 => n4680, CI => n1097, CO =>
                           n598, S0 => n599);
   U3005 : HS65_LH_MX41X7 port map( D0 => n1035, S0 => n4492, D1 => n4624, S1 
                           => n4608, D2 => n4622, S2 => n4604, D3 => n4620, S3 
                           => n4609, Z => n1065);
   U3006 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3071, Z => n1097);
   U3007 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1032, D1 => n4496, S1 
                           => n4627, D2 => n4499, S2 => n4629, D3 => n4504, S3 
                           => n4630, Z => n3071);
   U3008 : HS65_LH_FA1X4 port map( A0 => n1064, B0 => n4680, CI => n598, CO => 
                           n580, S0 => n581);
   U3009 : HS65_LH_MX41X7 port map( D0 => n1034, S0 => n4490, D1 => n4626, S1 
                           => n4608, D2 => n4624, S2 => n4602, D3 => n4622, S3 
                           => n4609, Z => n1064);
   U3010 : HS65_LH_FA1X4 port map( A0 => n1060, B0 => n4709, CI => n526, CO => 
                           n508, S0 => n509);
   U3011 : HS65_LH_MX41X7 port map( D0 => n1030, S0 => n4491, D1 => n4634, S1 
                           => n4607, D2 => n4632, S2 => n4603, D3 => n4630, S3 
                           => n4609, Z => n1060);
   U3012 : HS65_LH_FA1X4 port map( A0 => n1055, B0 => n4713, CI => n431, CO => 
                           n417, S0 => n418);
   U3013 : HS65_LH_MX41X7 port map( D0 => n1024, S0 => n4491, D1 => n4644, S1 
                           => n4602, D2 => n4642, S2 => n4610, D3 => n4646, S3 
                           => n4606, Z => n1055);
   U3014 : HS65_LH_FA1X4 port map( A0 => n1050, B0 => n4714, CI => n360, CO => 
                           n350, S0 => n351);
   U3015 : HS65_LH_MX41X7 port map( D0 => n1018, S0 => n4490, D1 => n4654, S1 
                           => n4609, D2 => n4656, S2 => n4602, D3 => n4658, S3 
                           => n4606, Z => n1050);
   U3016 : HS65_LH_FA1X4 port map( A0 => n1045, B0 => n4715, CI => n313, CO => 
                           n307, S0 => n308);
   U3017 : HS65_LH_MX41X7 port map( D0 => n1012, S0 => n4491, D1 => n4666, S1 
                           => n4610, D2 => n4668, S2 => n4603, D3 => n4670, S3 
                           => n4607, Z => n1045);
   U3018 : HS65_LH_MX41X7 port map( D0 => n4567, S0 => n1009, D1 => n4612, S1 
                           => n4677, D2 => n4564, S2 => n4675, D3 => n4561, S3 
                           => n4672, Z => n2836);
   U3019 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1028, D1 => n4507, S1 
                           => n4634, D2 => n4510, S2 => n4637, D3 => n4515, S3 
                           => n4638, Z => n3032);
   U3020 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1027, D1 => n4507, S1 
                           => n4636, D2 => n4510, S2 => n4639, D3 => n4515, S3 
                           => n4640, Z => n3033);
   U3021 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1022, D1 => n4528, S1 
                           => n4647, D2 => n4531, S2 => n4649, D3 => n4536, S3 
                           => n4650, Z => n2952);
   U3022 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1021, D1 => n4528, S1 
                           => n4649, D2 => n4532, S2 => n4651, D3 => n4536, S3 
                           => n4652, Z => n2953);
   U3023 : HS65_LH_MX41X7 port map( D0 => n3062, S0 => n1027, D1 => n4496, S1 
                           => n4637, D2 => n4499, S2 => n4639, D3 => n4504, S3 
                           => n4640, Z => n3076);
   U3024 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1010, D1 => n4570, S1 
                           => n4670, D2 => n4573, S2 => n4673, D3 => n4578, S3 
                           => n4674, Z => n2793);
   U3025 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1015, D1 => n4539, S1 
                           => n4661, D2 => n4542, S2 => n4663, D3 => n4547, S3 
                           => n4664, Z => n2916);
   U3026 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1021, D1 => n4506, S1 
                           => n4648, D2 => n4509, S2 => n4651, D3 => n4515, S3 
                           => n4652, Z => n3039);
   U3027 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1015, D1 => n4528, S1 
                           => n4660, D2 => n4531, S2 => n4663, D3 => n4536, S3 
                           => n4664, Z => n2959);
   U3028 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1021, D1 => n4495, S1 
                           => n4648, D2 => n4499, S2 => n4651, D3 => n4504, S3 
                           => n4652, Z => n3082);
   U3029 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1009, D1 => n4539, S1 
                           => n4672, D2 => n4542, S2 => n4675, D3 => n4547, S3 
                           => n4676, Z => n2922);
   U3030 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1015, D1 => n4506, S1 
                           => n4661, D2 => n4509, S2 => n4663, D3 => n4514, S3 
                           => n4664, Z => n3045);
   U3031 : HS65_LH_MX41X7 port map( D0 => n2933, S0 => n1009, D1 => n4529, S1 
                           => n4672, D2 => n4532, S2 => n4675, D3 => n4537, S3 
                           => n4677, Z => n2965);
   U3032 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1015, D1 => n4495, S1 
                           => n4660, D2 => n4498, S2 => n4663, D3 => n4503, S3 
                           => n4664, Z => n3088);
   U3033 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1009, D1 => n4506, S1 
                           => n4673, D2 => n4509, S2 => n4675, D3 => n4514, S3 
                           => n4676, Z => n3051);
   U3034 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1009, D1 => n4496, S1 
                           => n4673, D2 => n4499, S2 => n4675, D3 => n4504, S3 
                           => n4676, Z => n3094);
   U3035 : HS65_LH_MX41X7 port map( D0 => n2762, S0 => n1009, D1 => n4570, S1 
                           => n4673, D2 => n4573, S2 => n4675, D3 => n4579, S3 
                           => n4677, Z => n2794);
   U3036 : HS65_LH_MX41X7 port map( D0 => n2847, S0 => n1009, D1 => n4551, S1 
                           => n4673, D2 => n4554, S2 => n4675, D3 => n4560, S3 
                           => n4677, Z => n2879);
   U3037 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1021, D1 => n4526, S1 
                           => n4652, D2 => n4518, S2 => n4649, D3 => n4521, S3 
                           => n4650, Z => n2996);
   U3038 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1015, D1 => n4525, S1 
                           => n4664, D2 => n4517, S2 => n4661, D3 => n4520, S3 
                           => n4662, Z => n3002);
   U3039 : HS65_LH_MX41X7 port map( D0 => n2976, S0 => n1009, D1 => n4526, S1 
                           => n4677, D2 => n4518, S2 => n4673, D3 => n4521, S3 
                           => n4674, Z => n3008);
   U3040 : HS65_LH_FA1X4 port map( A0 => n4622, B0 => n4624, CI => n1003, CO =>
                           n1002, S0 => n1035);
   U3041 : HS65_LH_FA1X4 port map( A0 => n4624, B0 => n4626, CI => n1002, CO =>
                           n1001, S0 => n1034);
   U3042 : HS65_LH_FA1X4 port map( A0 => n4626, B0 => n4628, CI => n1001, CO =>
                           n1000, S0 => n1033);
   U3043 : HS65_LH_FA1X4 port map( A0 => n4628, B0 => n4630, CI => n1000, CO =>
                           n999, S0 => n1032);
   U3044 : HS65_LH_FA1X4 port map( A0 => n4630, B0 => n4632, CI => n999, CO => 
                           n998, S0 => n1031);
   U3045 : HS65_LH_FA1X4 port map( A0 => n4632, B0 => n4634, CI => n998, CO => 
                           n997, S0 => n1030);
   U3046 : HS65_LH_FA1X4 port map( A0 => n4634, B0 => n4636, CI => n997, CO => 
                           n996, S0 => n1029);
   U3047 : HS65_LH_FA1X4 port map( A0 => n4636, B0 => n4638, CI => n996, CO => 
                           n995, S0 => n1028);
   U3048 : HS65_LH_FA1X4 port map( A0 => n4638, B0 => n4640, CI => n995, CO => 
                           n994, S0 => n1027);
   U3049 : HS65_LH_FA1X4 port map( A0 => n4640, B0 => n4642, CI => n994, CO => 
                           n993, S0 => n1026);
   U3050 : HS65_LH_FA1X4 port map( A0 => n4642, B0 => n4644, CI => n993, CO => 
                           n992, S0 => n1025);
   U3051 : HS65_LH_FA1X4 port map( A0 => n4644, B0 => n4646, CI => n992, CO => 
                           n991, S0 => n1024);
   U3052 : HS65_LH_FA1X4 port map( A0 => n4646, B0 => n4648, CI => n991, CO => 
                           n990, S0 => n1023);
   U3053 : HS65_LH_FA1X4 port map( A0 => n4648, B0 => n4650, CI => n990, CO => 
                           n989, S0 => n1022);
   U3054 : HS65_LH_FA1X4 port map( A0 => n4650, B0 => n4652, CI => n989, CO => 
                           n988, S0 => n1021);
   U3055 : HS65_LH_FA1X4 port map( A0 => n4652, B0 => n4654, CI => n988, CO => 
                           n987, S0 => n1020);
   U3056 : HS65_LH_FA1X4 port map( A0 => n4654, B0 => n4656, CI => n987, CO => 
                           n986, S0 => n1019);
   U3057 : HS65_LH_FA1X4 port map( A0 => n4656, B0 => n4658, CI => n986, CO => 
                           n985, S0 => n1018);
   U3058 : HS65_LH_FA1X4 port map( A0 => n4658, B0 => n4660, CI => n985, CO => 
                           n984, S0 => n1017);
   U3059 : HS65_LH_FA1X4 port map( A0 => n4662, B0 => n4664, CI => n983, CO => 
                           n982, S0 => n1015);
   U3060 : HS65_LH_FA1X4 port map( A0 => n4664, B0 => n4666, CI => n982, CO => 
                           n981, S0 => n1014);
   U3061 : HS65_LH_FA1X4 port map( A0 => n4666, B0 => n4668, CI => n981, CO => 
                           n980, S0 => n1013);
   U3062 : HS65_LH_FA1X4 port map( A0 => n4668, B0 => n4670, CI => n980, CO => 
                           n979, S0 => n1012);
   U3063 : HS65_LH_FA1X4 port map( A0 => n4670, B0 => n4672, CI => n979, CO => 
                           n978, S0 => n1011);
   U3064 : HS65_LH_FA1X4 port map( A0 => n4672, B0 => n4674, CI => n978, CO => 
                           n977, S0 => n1010);
   U3065 : HS65_LH_FA1X4 port map( A0 => n297, B0 => n4708, CI => n1041, CO => 
                           n293, S0 => n294);
   U3066 : HS65_LH_MX41X7 port map( D0 => n1008, S0 => n4492, D1 => n4674, S1 
                           => n4609, D2 => n4676, S2 => n4604, D3 => n4606, S3 
                           => n4679, Z => n1041);
   U3067 : HS65_LH_FA1X4 port map( A0 => n557, B0 => n1191, CI => n1223, CO => 
                           n554, S0 => n555);
   U3068 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2913, Z => n1223);
   U3069 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2953, Z => n1191);
   U3070 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1018, D1 => n4539, S1 
                           => n4655, D2 => n4542, S2 => n4657, D3 => n4547, S3 
                           => n4658, Z => n2913);
   U3071 : HS65_LH_FA1X4 port map( A0 => n509, B0 => n1092, CI => n1124, CO => 
                           n506, S0 => n507);
   U3072 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3036, Z => n1124);
   U3073 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3076, Z => n1092);
   U3074 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1024, D1 => n4506, S1 
                           => n4642, D2 => n4509, S2 => n4645, D3 => n4515, S3 
                           => n4646, Z => n3036);
   U3075 : HS65_LH_FA1X4 port map( A0 => n553, B0 => n1255, CI => n568, CO => 
                           n550, S0 => n551);
   U3076 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2873, Z => n1255);
   U3077 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1015, D1 => n4550, S1 
                           => n4661, D2 => n4553, S2 => n4663, D3 => n4558, S3 
                           => n4664, Z => n2873);
   U3078 : HS65_LH_FA1X4 port map( A0 => n505, B0 => n1156, CI => n1188, CO => 
                           n502, S0 => n503);
   U3079 : HS65_LHS_XOR2X6 port map( A => n4698, B => n2956, Z => n1188);
   U3080 : HS65_LHS_XOR2X6 port map( A => n4701, B => n2996, Z => n1156);
   U3081 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1018, D1 => n4528, S1 
                           => n4655, D2 => n4531, S2 => n4657, D3 => n4536, S3 
                           => n4658, Z => n2956);
   U3082 : HS65_LH_FA1X4 port map( A0 => n501, B0 => n1220, CI => n1252, CO => 
                           n498, S0 => n499);
   U3083 : HS65_LHS_XOR2X6 port map( A => n4691, B => n2876, Z => n1252);
   U3084 : HS65_LHS_XOR2X6 port map( A => n4695, B => n2916, Z => n1220);
   U3085 : HS65_LH_MX41X7 port map( D0 => n4556, S0 => n1012, D1 => n4550, S1 
                           => n4667, D2 => n4553, S2 => n4669, D3 => n4558, S3 
                           => n4670, Z => n2876);
   U3086 : HS65_LH_FA1X4 port map( A0 => n459, B0 => n1121, CI => n1153, CO => 
                           n456, S0 => n457);
   U3087 : HS65_LHS_XOR2X6 port map( A => n4700, B => n2999, Z => n1153);
   U3088 : HS65_LHS_XOR2X6 port map( A => n4704, B => n3039, Z => n1121);
   U3089 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1018, D1 => n4525, S1 
                           => n4658, D2 => n4517, S2 => n4655, D3 => n4520, S3 
                           => n4656, Z => n2999);
   U3090 : HS65_LH_FA1X4 port map( A0 => n455, B0 => n1185, CI => n1217, CO => 
                           n452, S0 => n453);
   U3091 : HS65_LHS_XOR2X6 port map( A => n4694, B => n2919, Z => n1217);
   U3092 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2959, Z => n1185);
   U3093 : HS65_LH_MX41X7 port map( D0 => n4545, S0 => n1012, D1 => n4539, S1 
                           => n4666, D2 => n4543, S2 => n4669, D3 => n4548, S3 
                           => n4670, Z => n2919);
   U3094 : HS65_LH_FA1X4 port map( A0 => n418, B0 => n1086, CI => n1118, CO => 
                           n415, S0 => n416);
   U3095 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3042, Z => n1118);
   U3096 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3082, Z => n1086);
   U3097 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1018, D1 => n4506, S1 
                           => n4654, D2 => n4509, S2 => n4657, D3 => n4514, S3 
                           => n4658, Z => n3042);
   U3098 : HS65_LH_FA1X4 port map( A0 => n414, B0 => n1150, CI => n1182, CO => 
                           n411, S0 => n412);
   U3099 : HS65_LHS_XOR2X6 port map( A => n4697, B => n2962, Z => n1182);
   U3100 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3002, Z => n1150);
   U3101 : HS65_LH_MX41X7 port map( D0 => n4534, S0 => n1012, D1 => n4528, S1 
                           => n4666, D2 => n4531, S2 => n4669, D3 => n4536, S3 
                           => n4670, Z => n2962);
   U3102 : HS65_LH_FA1X4 port map( A0 => n380, B0 => n1115, CI => n1147, CO => 
                           n377, S0 => n378);
   U3103 : HS65_LHS_XOR2X6 port map( A => n4700, B => n3005, Z => n1147);
   U3104 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3045, Z => n1115);
   U3105 : HS65_LH_MX41X7 port map( D0 => n4523, S0 => n1012, D1 => n4525, S1 
                           => n4671, D2 => n4518, S2 => n4667, D3 => n4521, S3 
                           => n4668, Z => n3005);
   U3106 : HS65_LH_FA1X4 port map( A0 => n351, B0 => n1080, CI => n1112, CO => 
                           n348, S0 => n349);
   U3107 : HS65_LHS_XOR2X6 port map( A => n4703, B => n3048, Z => n1112);
   U3108 : HS65_LHS_XOR2X6 port map( A => n4707, B => n3088, Z => n1080);
   U3109 : HS65_LH_MX41X7 port map( D0 => n4512, S0 => n1012, D1 => n4506, S1 
                           => n4666, D2 => n4510, S2 => n4669, D3 => n4514, S3 
                           => n4670, Z => n3048);
   U3110 : HS65_LH_FA1X4 port map( A0 => n1063, B0 => n4680, CI => n580, CO => 
                           n562, S0 => n563);
   U3111 : HS65_LH_MX41X7 port map( D0 => n1033, S0 => n4492, D1 => n4628, S1 
                           => n4608, D2 => n4626, S2 => n4603, D3 => n4624, S3 
                           => n4609, Z => n1063);
   U3112 : HS65_LH_FA1X4 port map( A0 => n1057, B0 => n4710, CI => n1089, CO =>
                           n460, S0 => n461);
   U3113 : HS65_LH_MX41X7 port map( D0 => n1027, S0 => n4491, D1 => n4606, S1 
                           => n4640, D2 => n4638, S2 => n4603, D3 => n4636, S3 
                           => n4609, Z => n1057);
   U3114 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3079, Z => n1089);
   U3115 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1024, D1 => n4495, S1 
                           => n4642, D2 => n4498, S2 => n4645, D3 => n4503, S3 
                           => n4646, Z => n3079);
   U3116 : HS65_LH_FA1X4 port map( A0 => n1052, B0 => n4711, CI => n1083, CO =>
                           n381, S0 => n382);
   U3117 : HS65_LH_MX41X7 port map( D0 => n1021, S0 => n4490, D1 => n4648, S1 
                           => n4610, D2 => n4650, S2 => n4602, D3 => n4652, S3 
                           => n4606, Z => n1052);
   U3118 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3085, Z => n1083);
   U3119 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1018, D1 => n4495, S1 
                           => n4654, D2 => n4498, S2 => n4657, D3 => n4503, S3 
                           => n4658, Z => n3085);
   U3120 : HS65_LH_FA1X4 port map( A0 => n1047, B0 => n4712, CI => n1077, CO =>
                           n326, S0 => n327);
   U3121 : HS65_LH_MX41X7 port map( D0 => n1015, S0 => n4490, D1 => n4660, S1 
                           => n4610, D2 => n4662, S2 => n4602, D3 => n4664, S3 
                           => n4606, Z => n1047);
   U3122 : HS65_LHS_XOR2X6 port map( A => n4706, B => n3091, Z => n1077);
   U3123 : HS65_LH_MX41X7 port map( D0 => n4501, S0 => n1012, D1 => n4495, S1 
                           => n4666, D2 => n4498, S2 => n4669, D3 => n4503, S3 
                           => n4670, Z => n3091);
   U3124 : HS65_LH_FA1X4 port map( A0 => n1042, B0 => n4716, CI => n1071, CO =>
                           n295, S0 => n296);
   U3125 : HS65_LH_MX41X7 port map( D0 => n1009, S0 => n4490, D1 => n4672, S1 
                           => n4609, D2 => n4674, S2 => n4602, D3 => n4676, S3 
                           => n4606, Z => n1042);
   U3126 : HS65_LHS_XOR2X6 port map( A => n4708, B => n3102, Z => n1071);
   U3127 : HS65_LH_AOI22X6 port map( A => n4501, B => n1006, C => n4495, D => 
                           n4678, Z => n3102);
   U3128 : HS65_LH_IVX9 port map( A => a(8), Z => n4687);
   U3129 : HS65_LH_IVX9 port map( A => a(14), Z => n4693);
   U3130 : HS65_LH_IVX9 port map( A => a(17), Z => n4696);
   U3131 : HS65_LH_IVX9 port map( A => a(29), Z => n4708);
   U3132 : HS65_LH_IVX9 port map( A => a(20), Z => n4699);
   U3133 : HS65_LH_IVX9 port map( A => a(11), Z => n4690);
   U3134 : HS65_LH_IVX9 port map( A => a(26), Z => n4705);
   U3135 : HS65_LH_IVX9 port map( A => a(23), Z => n4702);
   U3136 : HS65_LH_IVX9 port map( A => n4587, Z => n4586);
   U3137 : HS65_LH_IVX9 port map( A => n4576, Z => n4575);
   U3138 : HS65_LH_IVX9 port map( A => n4568, Z => n4567);
   U3139 : HS65_LH_IVX9 port map( A => n4557, Z => n4556);
   U3140 : HS65_LH_IVX9 port map( A => n4546, Z => n4545);
   U3141 : HS65_LH_IVX9 port map( A => n4535, Z => n4534);
   U3142 : HS65_LH_IVX9 port map( A => n4524, Z => n4523);
   U3143 : HS65_LH_IVX9 port map( A => n4513, Z => n4512);
   U3144 : HS65_LH_IVX9 port map( A => n4502, Z => n4501);
   U3145 : HS65_LH_BFX9 port map( A => b(30), Z => n4676);
   U3146 : HS65_LH_AND2X4 port map( A => n4594, B => n4679, Z => n2715);
   U3147 : HS65_LH_BFX9 port map( A => n2723, Z => n4580);
   U3148 : HS65_LH_BFX9 port map( A => n2766, Z => n4569);
   U3149 : HS65_LH_BFX9 port map( A => n2851, Z => n4550);
   U3150 : HS65_LH_BFX9 port map( A => n2894, Z => n4539);
   U3151 : HS65_LH_BFX9 port map( A => n2937, Z => n4528);
   U3152 : HS65_LH_BFX9 port map( A => n3023, Z => n4506);
   U3153 : HS65_LH_BFX9 port map( A => n3066, Z => n4495);
   U3154 : HS65_LH_BFX9 port map( A => n2808, Z => n4561);
   U3155 : HS65_LH_BFX9 port map( A => n2980, Z => n4517);
   U3156 : HS65_LH_BFX9 port map( A => b(31), Z => n4678);
   U3157 : HS65_LH_BFX9 port map( A => n2980, Z => n4518);
   U3158 : HS65_LH_BFX9 port map( A => n2723, Z => n4581);
   U3159 : HS65_LH_BFX9 port map( A => n3066, Z => n4496);
   U3160 : HS65_LH_BFX9 port map( A => n2894, Z => n4540);
   U3161 : HS65_LH_BFX9 port map( A => n2766, Z => n4570);
   U3162 : HS65_LH_BFX9 port map( A => n3023, Z => n4507);
   U3163 : HS65_LH_BFX9 port map( A => n2851, Z => n4551);
   U3164 : HS65_LH_BFX9 port map( A => n2937, Z => n4529);
   U3165 : HS65_LH_BFX9 port map( A => n2808, Z => n4562);
   U3166 : HS65_LH_BFX9 port map( A => b(3), Z => n4622);
   U3167 : HS65_LH_BFX9 port map( A => b(23), Z => n4662);
   U3168 : HS65_LH_BFX9 port map( A => b(2), Z => n4620);
   U3169 : HS65_LH_BFX9 port map( A => b(22), Z => n4660);
   U3170 : HS65_LH_BFX9 port map( A => b(29), Z => n4674);
   U3171 : HS65_LH_BFX9 port map( A => b(0), Z => n4614);
   U3172 : HS65_LH_BFX9 port map( A => b(1), Z => n4618);
   U3173 : HS65_LH_BFX9 port map( A => n4718, Z => n4493);
   U3174 : HS65_LH_BFX9 port map( A => n2417, Z => n4611);
   U3175 : HS65_LH_BFX9 port map( A => n2417, Z => n4612);
   U3176 : HS65_LH_BFX9 port map( A => n2975, Z => n4526);
   U3177 : HS65_LH_BFX9 port map( A => n2975, Z => n4525);
   U3178 : HS65_LH_BFX9 port map( A => n2932, Z => n4537);
   U3179 : HS65_LH_BFX9 port map( A => n2718, Z => n4589);
   U3180 : HS65_LH_BFX9 port map( A => n2846, Z => n4559);
   U3181 : HS65_LH_BFX9 port map( A => n3061, Z => n4504);
   U3182 : HS65_LH_BFX9 port map( A => n2761, Z => n4577);
   U3183 : HS65_LH_BFX9 port map( A => n2761, Z => n4578);
   U3184 : HS65_LH_BFX9 port map( A => n2718, Z => n4588);
   U3185 : HS65_LH_BFX9 port map( A => n3018, Z => n4515);
   U3186 : HS65_LH_BFX9 port map( A => n2889, Z => n4547);
   U3187 : HS65_LH_BFX9 port map( A => n2846, Z => n4558);
   U3188 : HS65_LH_BFX9 port map( A => n2889, Z => n4548);
   U3189 : HS65_LH_BFX9 port map( A => n2932, Z => n4536);
   U3190 : HS65_LH_BFX9 port map( A => n3018, Z => n4514);
   U3191 : HS65_LH_BFX9 port map( A => n3061, Z => n4503);
   U3192 : HS65_LH_BFX9 port map( A => n4717, Z => n4491);
   U3193 : HS65_LH_BFX9 port map( A => b(31), Z => n4679);
   U3194 : HS65_LH_BFX9 port map( A => n4717, Z => n4490);
   U3195 : HS65_LH_BFX9 port map( A => b(3), Z => n4623);
   U3196 : HS65_LH_BFX9 port map( A => b(2), Z => n4621);
   U3197 : HS65_LH_BFX9 port map( A => b(23), Z => n4663);
   U3198 : HS65_LH_BFX9 port map( A => b(30), Z => n4677);
   U3199 : HS65_LH_BFX9 port map( A => b(22), Z => n4661);
   U3200 : HS65_LH_BFX9 port map( A => b(29), Z => n4675);
   U3201 : HS65_LH_BFX9 port map( A => b(1), Z => n4619);
   U3202 : HS65_LH_BFX9 port map( A => n4718, Z => n4494);
   U3203 : HS65_LH_BFX9 port map( A => n4582, Z => n4584);
   U3204 : HS65_LH_BFX9 port map( A => n4571, Z => n4573);
   U3205 : HS65_LH_BFX9 port map( A => n4563, Z => n4565);
   U3206 : HS65_LH_BFX9 port map( A => n4552, Z => n4554);
   U3207 : HS65_LH_BFX9 port map( A => n4497, Z => n4499);
   U3208 : HS65_LH_BFX9 port map( A => n4571, Z => n4572);
   U3209 : HS65_LH_BFX9 port map( A => n4563, Z => n4564);
   U3210 : HS65_LH_BFX9 port map( A => n4582, Z => n4583);
   U3211 : HS65_LH_BFX9 port map( A => n4541, Z => n4542);
   U3212 : HS65_LH_BFX9 port map( A => n4552, Z => n4553);
   U3213 : HS65_LH_BFX9 port map( A => n4541, Z => n4543);
   U3214 : HS65_LH_BFX9 port map( A => n4508, Z => n4509);
   U3215 : HS65_LH_BFX9 port map( A => n4530, Z => n4532);
   U3216 : HS65_LH_BFX9 port map( A => n4530, Z => n4531);
   U3217 : HS65_LH_BFX9 port map( A => n4508, Z => n4510);
   U3218 : HS65_LH_BFX9 port map( A => n4497, Z => n4498);
   U3219 : HS65_LH_BFX9 port map( A => n4601, Z => n4602);
   U3220 : HS65_LH_BFX9 port map( A => n4519, Z => n4520);
   U3221 : HS65_LH_BFX9 port map( A => n4519, Z => n4521);
   U3222 : HS65_LH_BFX9 port map( A => n4601, Z => n4603);
   U3223 : HS65_LH_BFX9 port map( A => n2975, Z => n4527);
   U3224 : HS65_LH_BFX9 port map( A => n2718, Z => n4590);
   U3225 : HS65_LH_BFX9 port map( A => n2761, Z => n4579);
   U3226 : HS65_LH_BFX9 port map( A => n2846, Z => n4560);
   U3227 : HS65_LH_BFX9 port map( A => n2889, Z => n4549);
   U3228 : HS65_LH_BFX9 port map( A => n2932, Z => n4538);
   U3229 : HS65_LH_BFX9 port map( A => n3018, Z => n4516);
   U3230 : HS65_LH_BFX9 port map( A => n3061, Z => n4505);
   U3231 : HS65_LH_BFX9 port map( A => n2417, Z => n4613);
   U3232 : HS65_LH_BFX9 port map( A => n4717, Z => n4492);
   U3233 : HS65_LH_BFX9 port map( A => n4582, Z => n4585);
   U3234 : HS65_LH_BFX9 port map( A => n4571, Z => n4574);
   U3235 : HS65_LH_BFX9 port map( A => n4552, Z => n4555);
   U3236 : HS65_LH_BFX9 port map( A => n4541, Z => n4544);
   U3237 : HS65_LH_BFX9 port map( A => n4530, Z => n4533);
   U3238 : HS65_LH_BFX9 port map( A => n4508, Z => n4511);
   U3239 : HS65_LH_BFX9 port map( A => n4497, Z => n4500);
   U3240 : HS65_LH_BFX9 port map( A => n4563, Z => n4566);
   U3241 : HS65_LH_BFX9 port map( A => n4519, Z => n4522);
   U3242 : HS65_LH_BFX9 port map( A => n4601, Z => n4604);
   U3243 : HS65_LH_IVX9 port map( A => n2673, Z => n4717);
   U3244 : HS65_LH_IVX9 port map( A => n2713, Z => n4718);
   U3245 : HS65_LH_IVX9 port map( A => n2719, Z => n4587);
   U3246 : HS65_LH_NOR2AX3 port map( A => n2753, B => n2754, Z => n2719);
   U3247 : HS65_LH_IVX9 port map( A => n2762, Z => n4576);
   U3248 : HS65_LH_NOR2AX3 port map( A => n2796, B => n2797, Z => n2762);
   U3249 : HS65_LH_IVX9 port map( A => n2804, Z => n4568);
   U3250 : HS65_LH_NOR2AX3 port map( A => n2838, B => n2839, Z => n2804);
   U3251 : HS65_LH_IVX9 port map( A => n2847, Z => n4557);
   U3252 : HS65_LH_NOR2AX3 port map( A => n2881, B => n2882, Z => n2847);
   U3253 : HS65_LH_IVX9 port map( A => n2890, Z => n4546);
   U3254 : HS65_LH_NOR2AX3 port map( A => n2924, B => n2925, Z => n2890);
   U3255 : HS65_LH_IVX9 port map( A => n2933, Z => n4535);
   U3256 : HS65_LH_NOR2AX3 port map( A => n2967, B => n2968, Z => n2933);
   U3257 : HS65_LH_IVX9 port map( A => n2976, Z => n4524);
   U3258 : HS65_LH_NOR2AX3 port map( A => n3010, B => n3011, Z => n2976);
   U3259 : HS65_LH_IVX9 port map( A => n3019, Z => n4513);
   U3260 : HS65_LH_NOR2AX3 port map( A => n3053, B => n3054, Z => n3019);
   U3261 : HS65_LH_IVX9 port map( A => n3062, Z => n4502);
   U3262 : HS65_LH_NOR2AX3 port map( A => n3096, B => n3097, Z => n3062);
   U3263 : HS65_LH_IVX9 port map( A => n4682, Z => n4680);
   U3264 : HS65_LH_IVX9 port map( A => a(2), Z => n4682);
   U3265 : HS65_LH_IVX9 port map( A => n4682, Z => n4681);
   U3266 : HS65_LH_FA1X4 port map( A0 => n1387, B0 => n619, CI => n258, CO => 
                           n257, S0 => product(32));
   U3267 : HS65_LHS_XOR2X6 port map( A => n4681, B => n2712, Z => n1387);
   U3268 : HS65_LH_OAI21X3 port map( A => n4719, B => n2713, C => n2714, Z => 
                           n2712);
   U3269 : HS65_LH_OAI22X6 port map( A => n4676, B => n2715, C => n4591, D => 
                           n2715, Z => n2714);
   U3270 : HS65_LH_OA12X9 port map( A => n2673, B => n4719, C => n2674, Z => 
                           n292);
   U3271 : HS65_LH_OAI22X6 port map( A => n4676, B => n2675, C => n4609, D => 
                           n2675, Z => n2674);
   U3272 : HS65_LH_AND2X4 port map( A => n4678, B => n4602, Z => n2675);
   U3273 : HS65_LH_BFX9 port map( A => n2670, Z => n4609);
   U3274 : HS65_LH_BFX9 port map( A => n2681, Z => n4591);
   U3275 : HS65_LH_BFX9 port map( A => n2672, Z => n4601);
   U3276 : HS65_LH_NOR2AX3 port map( A => n3104, B => n3103, Z => n2672);
   U3277 : HS65_LH_BFX9 port map( A => n2721, Z => n4582);
   U3278 : HS65_LH_NOR2X6 port map( A => n2753, B => n2758, Z => n2721);
   U3279 : HS65_LH_BFX9 port map( A => n2764, Z => n4571);
   U3280 : HS65_LH_NOR2X6 port map( A => n2796, B => n2801, Z => n2764);
   U3281 : HS65_LH_BFX9 port map( A => n2806, Z => n4563);
   U3282 : HS65_LH_NOR2X6 port map( A => n2838, B => n2843, Z => n2806);
   U3283 : HS65_LH_BFX9 port map( A => n2849, Z => n4552);
   U3284 : HS65_LH_NOR2X6 port map( A => n2881, B => n2886, Z => n2849);
   U3285 : HS65_LH_BFX9 port map( A => n2892, Z => n4541);
   U3286 : HS65_LH_NOR2X6 port map( A => n2924, B => n2929, Z => n2892);
   U3287 : HS65_LH_BFX9 port map( A => n2935, Z => n4530);
   U3288 : HS65_LH_NOR2X6 port map( A => n2967, B => n2972, Z => n2935);
   U3289 : HS65_LH_BFX9 port map( A => n2978, Z => n4519);
   U3290 : HS65_LH_NOR2X6 port map( A => n3010, B => n3015, Z => n2978);
   U3291 : HS65_LH_BFX9 port map( A => n3021, Z => n4508);
   U3292 : HS65_LH_NOR2X6 port map( A => n3053, B => n3058, Z => n3021);
   U3293 : HS65_LH_BFX9 port map( A => n3064, Z => n4497);
   U3294 : HS65_LH_NOR2X6 port map( A => n3096, B => n3101, Z => n3064);
   U3295 : HS65_LH_BFX9 port map( A => n2681, Z => n4592);
   U3296 : HS65_LH_BFX9 port map( A => b(27), Z => n4670);
   U3297 : HS65_LH_BFX9 port map( A => b(19), Z => n4654);
   U3298 : HS65_LH_BFX9 port map( A => b(15), Z => n4646);
   U3299 : HS65_LH_BFX9 port map( A => b(4), Z => n4624);
   U3300 : HS65_LH_BFX9 port map( A => b(5), Z => n4626);
   U3301 : HS65_LH_BFX9 port map( A => b(17), Z => n4650);
   U3302 : HS65_LH_BFX9 port map( A => b(7), Z => n4630);
   U3303 : HS65_LH_BFX9 port map( A => b(11), Z => n4638);
   U3304 : HS65_LH_BFX9 port map( A => b(21), Z => n4658);
   U3305 : HS65_LH_BFX9 port map( A => b(9), Z => n4634);
   U3306 : HS65_LH_BFX9 port map( A => b(28), Z => n4672);
   U3307 : HS65_LH_BFX9 port map( A => b(25), Z => n4666);
   U3308 : HS65_LH_BFX9 port map( A => b(18), Z => n4652);
   U3309 : HS65_LH_BFX9 port map( A => b(26), Z => n4668);
   U3310 : HS65_LH_BFX9 port map( A => b(13), Z => n4642);
   U3311 : HS65_LH_BFX9 port map( A => b(24), Z => n4664);
   U3312 : HS65_LH_BFX9 port map( A => b(20), Z => n4656);
   U3313 : HS65_LH_BFX9 port map( A => b(6), Z => n4628);
   U3314 : HS65_LH_BFX9 port map( A => b(10), Z => n4636);
   U3315 : HS65_LH_BFX9 port map( A => b(8), Z => n4632);
   U3316 : HS65_LH_BFX9 port map( A => b(16), Z => n4648);
   U3317 : HS65_LH_BFX9 port map( A => b(12), Z => n4640);
   U3318 : HS65_LH_BFX9 port map( A => b(14), Z => n4644);
   U3319 : HS65_LH_BFX9 port map( A => n2670, Z => n4610);
   U3320 : HS65_LH_BFX9 port map( A => b(27), Z => n4671);
   U3321 : HS65_LH_BFX9 port map( A => b(19), Z => n4655);
   U3322 : HS65_LH_BFX9 port map( A => b(25), Z => n4667);
   U3323 : HS65_LH_BFX9 port map( A => b(15), Z => n4647);
   U3324 : HS65_LH_BFX9 port map( A => b(4), Z => n4625);
   U3325 : HS65_LH_BFX9 port map( A => b(5), Z => n4627);
   U3326 : HS65_LH_BFX9 port map( A => b(17), Z => n4651);
   U3327 : HS65_LH_BFX9 port map( A => b(7), Z => n4631);
   U3328 : HS65_LH_BFX9 port map( A => b(11), Z => n4639);
   U3329 : HS65_LH_BFX9 port map( A => b(21), Z => n4659);
   U3330 : HS65_LH_BFX9 port map( A => b(12), Z => n4641);
   U3331 : HS65_LH_BFX9 port map( A => b(9), Z => n4635);
   U3332 : HS65_LH_BFX9 port map( A => b(28), Z => n4673);
   U3333 : HS65_LH_BFX9 port map( A => b(13), Z => n4643);
   U3334 : HS65_LH_BFX9 port map( A => b(18), Z => n4653);
   U3335 : HS65_LH_BFX9 port map( A => b(26), Z => n4669);
   U3336 : HS65_LH_BFX9 port map( A => b(24), Z => n4665);
   U3337 : HS65_LH_BFX9 port map( A => b(20), Z => n4657);
   U3338 : HS65_LH_BFX9 port map( A => b(14), Z => n4645);
   U3339 : HS65_LH_BFX9 port map( A => b(6), Z => n4629);
   U3340 : HS65_LH_BFX9 port map( A => b(10), Z => n4637);
   U3341 : HS65_LH_BFX9 port map( A => b(8), Z => n4633);
   U3342 : HS65_LH_BFX9 port map( A => b(16), Z => n4649);
   U3343 : HS65_LH_BFX9 port map( A => n4593, Z => n4594);
   U3344 : HS65_LH_BFX9 port map( A => n4597, Z => n4598);
   U3345 : HS65_LH_BFX9 port map( A => n4593, Z => n4595);
   U3346 : HS65_LH_BFX9 port map( A => n4605, Z => n4606);
   U3347 : HS65_LH_BFX9 port map( A => n4597, Z => n4599);
   U3348 : HS65_LH_BFX9 port map( A => n4605, Z => n4607);
   U3349 : HS65_LH_BFX9 port map( A => n4597, Z => n4600);
   U3350 : HS65_LH_BFX9 port map( A => n4605, Z => n4608);
   U3351 : HS65_LH_BFX9 port map( A => n4593, Z => n4596);
   U3352 : HS65_LHS_XOR3X2 port map( A => n292, B => n227, C => n2669, Z => 
                           product(63));
   U3353 : HS65_LH_AO22X9 port map( A => n4678, B => n4610, C => n4490, D => 
                           n1006, Z => n2669);
   U3354 : HS65_LHS_XOR2X6 port map( A => n4706, B => a(30), Z => n3103);
   U3355 : HS65_LHS_XOR2X6 port map( A => n4685, B => a(9), Z => n2838);
   U3356 : HS65_LHS_XOR2X6 port map( A => n4691, B => a(15), Z => n2924);
   U3357 : HS65_LHS_XOR2X6 port map( A => n4680, B => a(3), Z => n2753);
   U3358 : HS65_LHS_XOR2X6 port map( A => n4695, B => a(18), Z => n2967);
   U3359 : HS65_LHS_XOR2X6 port map( A => n4688, B => a(12), Z => n2881);
   U3360 : HS65_LHS_XOR2X6 port map( A => n4697, B => a(21), Z => n3010);
   U3361 : HS65_LHS_XOR2X6 port map( A => n4703, B => a(27), Z => n3096);
   U3362 : HS65_LHS_XOR2X6 port map( A => n4700, B => a(24), Z => n3053);
   U3363 : HS65_LHS_XOR2X6 port map( A => a(5), B => a(6), Z => n2796);
   U3364 : HS65_LHS_XOR2X6 port map( A => n4681, B => a(1), Z => n2711);
   U3365 : HS65_LHS_XNOR2X6 port map( A => a(8), B => a(7), Z => n2797);
   U3366 : HS65_LHS_XNOR2X6 port map( A => a(14), B => a(13), Z => n2882);
   U3367 : HS65_LHS_XNOR2X6 port map( A => a(11), B => a(10), Z => n2839);
   U3368 : HS65_LHS_XNOR2X6 port map( A => a(17), B => a(16), Z => n2925);
   U3369 : HS65_LHS_XNOR2X6 port map( A => a(20), B => a(19), Z => n2968);
   U3370 : HS65_LHS_XNOR2X6 port map( A => a(26), B => a(25), Z => n3054);
   U3371 : HS65_LHS_XNOR2X6 port map( A => a(29), B => a(28), Z => n3097);
   U3372 : HS65_LHS_XNOR2X6 port map( A => a(23), B => a(22), Z => n3011);
   U3373 : HS65_LHS_XNOR2X6 port map( A => a(5), B => a(4), Z => n2754);
   U3374 : HS65_LHS_XOR2X6 port map( A => a(31), B => a(30), Z => n3104);
   U3375 : HS65_LHS_XNOR2X6 port map( A => a(4), B => a(3), Z => n2758);
   U3376 : HS65_LHS_XNOR2X6 port map( A => a(7), B => a(6), Z => n2801);
   U3377 : HS65_LHS_XNOR2X6 port map( A => a(9), B => a(10), Z => n2843);
   U3378 : HS65_LHS_XNOR2X6 port map( A => a(13), B => a(12), Z => n2886);
   U3379 : HS65_LHS_XNOR2X6 port map( A => a(16), B => a(15), Z => n2929);
   U3380 : HS65_LHS_XNOR2X6 port map( A => a(19), B => a(18), Z => n2972);
   U3381 : HS65_LHS_XNOR2X6 port map( A => a(22), B => a(21), Z => n3015);
   U3382 : HS65_LHS_XNOR2X6 port map( A => a(25), B => a(24), Z => n3058);
   U3383 : HS65_LHS_XNOR2X6 port map( A => a(28), B => a(27), Z => n3101);
   U3384 : HS65_LH_NAND2X7 port map( A => a(0), B => n2711, Z => n2713);
   U3385 : HS65_LH_NAND2X7 port map( A => a(31), B => n3103, Z => n2673);
   U3386 : HS65_LH_BFX9 port map( A => n2677, Z => n4597);
   U3387 : HS65_LH_NOR2AX3 port map( A => a(0), B => n2711, Z => n2677);
   U3388 : HS65_LH_BFX9 port map( A => n2671, Z => n4605);
   U3389 : HS65_LH_NOR2AX3 port map( A => n3103, B => a(31), Z => n2671);
   U3390 : HS65_LH_BFX9 port map( A => n2679, Z => n4593);
   U3391 : HS65_LH_NOR2AX3 port map( A => a(1), B => a(0), Z => n2679);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_add_0;

architecture SYN_rpl of alu_DW01_add_0 is

   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1 : std_logic;

begin
   
   U1_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => B(30), CI => 
                           carry_30_port, CO => carry_31_port, S0 => SUM(30));
   U1_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => B(28), CI => 
                           carry_28_port, CO => carry_29_port, S0 => SUM(28));
   U1_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => B(27), CI => 
                           carry_27_port, CO => carry_28_port, S0 => SUM(27));
   U1_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => B(25), CI => 
                           carry_25_port, CO => carry_26_port, S0 => SUM(25));
   U1_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => B(24), CI => 
                           carry_24_port, CO => carry_25_port, S0 => SUM(24));
   U1_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => B(22), CI => 
                           carry_22_port, CO => carry_23_port, S0 => SUM(22));
   U1_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => B(21), CI => 
                           carry_21_port, CO => carry_22_port, S0 => SUM(21));
   U1_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => B(19), CI => 
                           carry_19_port, CO => carry_20_port, S0 => SUM(19));
   U1_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => B(18), CI => 
                           carry_18_port, CO => carry_19_port, S0 => SUM(18));
   U1_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => B(12), CI => 
                           carry_12_port, CO => carry_13_port, S0 => SUM(12));
   U1_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => B(10), CI => 
                           carry_10_port, CO => carry_11_port, S0 => SUM(10));
   U1_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => B(9), CI => carry_9_port, 
                           CO => carry_10_port, S0 => SUM(9));
   U1_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => B(7), CI => carry_7_port, 
                           CO => carry_8_port, S0 => SUM(7));
   U1_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => B(6), CI => carry_6_port, 
                           CO => carry_7_port, S0 => SUM(6));
   U1_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => B(4), CI => carry_4_port, 
                           CO => carry_5_port, S0 => SUM(4));
   U1_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => B(3), CI => carry_3_port, 
                           CO => carry_4_port, S0 => SUM(3));
   U1_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => B(16), CI => 
                           carry_16_port, CO => carry_17_port, S0 => SUM(16));
   U1_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => B(1), CI => n1, CO => 
                           carry_2_port, S0 => SUM(1));
   U1_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => B(15), CI => 
                           carry_15_port, CO => carry_16_port, S0 => SUM(15));
   U1_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => B(13), CI => 
                           carry_13_port, CO => carry_14_port, S0 => SUM(13));
   U1_31 : HS65_LHS_XOR3X2 port map( A => A(31), B => B(31), C => carry_31_port
                           , Z => SUM(31));
   U1_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => B(2), CI => carry_2_port, 
                           CO => carry_3_port, S0 => SUM(2));
   U1_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => B(23), CI => 
                           carry_23_port, CO => carry_24_port, S0 => SUM(23));
   U1_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => B(29), CI => 
                           carry_29_port, CO => carry_30_port, S0 => SUM(29));
   U1_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => B(26), CI => 
                           carry_26_port, CO => carry_27_port, S0 => SUM(26));
   U1_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => B(20), CI => 
                           carry_20_port, CO => carry_21_port, S0 => SUM(20));
   U1_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => B(17), CI => 
                           carry_17_port, CO => carry_18_port, S0 => SUM(17));
   U1_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => B(11), CI => 
                           carry_11_port, CO => carry_12_port, S0 => SUM(11));
   U1_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => B(5), CI => carry_5_port, 
                           CO => carry_6_port, S0 => SUM(5));
   U1_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => B(8), CI => carry_8_port, 
                           CO => carry_9_port, S0 => SUM(8));
   U1_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => B(14), CI => 
                           carry_14_port, CO => carry_15_port, S0 => SUM(14));
   U1 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => SUM(0));
   U2 : HS65_LH_AND2X4 port map( A => A(0), B => B(0), Z => n1);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end alu_DW01_cmp6_0;

architecture SYN_rpl of alu_DW01_cmp6_0 is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2AX7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND4X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   signal LT_port, EQ_port, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n364, n365, n366, n367, n368, 
      n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405 : 
      std_logic;

begin
   LT <= LT_port;
   EQ <= EQ_port;
   
   U1 : HS65_LH_NAND2X7 port map( A => A(5), B => n366, Z => n106);
   U2 : HS65_LH_NAND2X7 port map( A => A(29), B => n381, Z => n62);
   U3 : HS65_LH_NAND2X7 port map( A => A(11), B => n369, Z => n54);
   U4 : HS65_LH_NAND2X7 port map( A => A(20), B => n375, Z => n74);
   U5 : HS65_LH_NAND2X7 port map( A => A(23), B => n377, Z => n72);
   U6 : HS65_LH_NAND2X7 port map( A => A(17), B => n373, Z => n69);
   U7 : HS65_LH_IVX9 port map( A => B(3), Z => n365);
   U8 : HS65_LH_IVX9 port map( A => B(2), Z => n364);
   U9 : HS65_LH_IVX9 port map( A => B(23), Z => n377);
   U10 : HS65_LH_IVX9 port map( A => B(29), Z => n381);
   U11 : HS65_LH_IVX9 port map( A => A(8), Z => n383);
   U12 : HS65_LH_IVX9 port map( A => B(31), Z => n382);
   U13 : HS65_LH_IVX9 port map( A => A(14), Z => n384);
   U14 : HS65_LH_IVX9 port map( A => A(26), Z => n385);
   U15 : HS65_LH_IVX9 port map( A => n115, Z => n403);
   U16 : HS65_LH_NOR4ABX2 port map( A => n76, B => n77, C => n78, D => LT_port,
                           Z => n43);
   U17 : HS65_LH_AND2X4 port map( A => n114, B => n109, Z => n77);
   U18 : HS65_LH_NAND4ABX3 port map( A => n115, B => n401, C => n106, D => n105
                           , Z => n78);
   U19 : HS65_LH_IVX9 port map( A => n102, Z => n401);
   U20 : HS65_LH_NOR4ABX2 port map( A => n55, B => n56, C => n57, D => n58, Z 
                           => n44);
   U21 : HS65_LH_AND4X6 port map( A => n72, B => n73, C => n74, D => n75, Z => 
                           n55);
   U22 : HS65_LH_NAND4ABX3 port map( A => n59, B => n60, C => n61, D => n62, Z 
                           => n58);
   U23 : HS65_LH_NAND4ABX3 port map( A => n64, B => n390, C => n65, D => n66, Z
                           => n57);
   U24 : HS65_LH_NOR4ABX2 port map( A => n68, B => n69, C => n70, D => n71, Z 
                           => n56);
   U25 : HS65_LH_NOR2X6 port map( A => B(18), B => n395, Z => n70);
   U26 : HS65_LH_NAND4ABX3 port map( A => n51, B => n398, C => n52, D => n53, Z
                           => n45);
   U27 : HS65_LH_IVX9 port map( A => n54, Z => n398);
   U28 : HS65_LH_NOR2X6 port map( A => n397, B => B(16), Z => n71);
   U29 : HS65_LH_NOR2X6 port map( A => n389, B => B(30), Z => n60);
   U30 : HS65_LH_NOR2X6 port map( A => n404, B => B(4), Z => n115);
   U31 : HS65_LH_NOR2X6 port map( A => n392, B => B(24), Z => n64);
   U32 : HS65_LH_NOR2X6 port map( A => n383, B => B(8), Z => n51);
   U33 : HS65_LH_IVX9 port map( A => EQ_port, Z => NE);
   U34 : HS65_LH_NOR4ABX2 port map( A => n43, B => n44, C => n45, D => n46, Z 
                           => EQ_port);
   U35 : HS65_LH_OR2X9 port map( A => B(26), B => n385, Z => n66);
   U36 : HS65_LH_NAND2X7 port map( A => A(2), B => n364, Z => n114);
   U37 : HS65_LH_OR2X9 port map( A => B(14), B => n384, Z => n50);
   U38 : HS65_LH_IVX9 port map( A => B(19), Z => n374);
   U39 : HS65_LH_IVX9 port map( A => B(27), Z => n379);
   U40 : HS65_LH_IVX9 port map( A => B(25), Z => n378);
   U41 : HS65_LH_IVX9 port map( A => B(12), Z => n370);
   U42 : HS65_LH_IVX9 port map( A => B(15), Z => n372);
   U43 : HS65_LH_IVX9 port map( A => B(20), Z => n375);
   U44 : HS65_LH_IVX9 port map( A => B(13), Z => n371);
   U45 : HS65_LH_IVX9 port map( A => B(5), Z => n366);
   U46 : HS65_LH_IVX9 port map( A => B(17), Z => n373);
   U47 : HS65_LH_IVX9 port map( A => B(7), Z => n367);
   U48 : HS65_LH_IVX9 port map( A => B(11), Z => n369);
   U49 : HS65_LH_IVX9 port map( A => B(28), Z => n380);
   U50 : HS65_LH_IVX9 port map( A => B(21), Z => n376);
   U51 : HS65_LH_IVX9 port map( A => B(9), Z => n368);
   U52 : HS65_LH_NAND4X9 port map( A => n47, B => n48, C => n49, D => n50, Z =>
                           n46);
   U53 : HS65_LH_IVX9 port map( A => n67, Z => n390);
   U54 : HS65_LH_OAI22X6 port map( A => A(31), B => n382, C => n387, D => n79, 
                           Z => LT_port);
   U55 : HS65_LH_IVX9 port map( A => n76, Z => n387);
   U56 : HS65_LH_AOI32X5 port map( A => n62, B => n388, C => n80, D => B(30), E
                           => n389, Z => n79);
   U57 : HS65_LH_IVX9 port map( A => n60, Z => n388);
   U58 : HS65_LH_OAI212X5 port map( A => A(2), B => n364, C => A(3), D => n365,
                           E => n111, Z => n110);
   U59 : HS65_LH_OAI212X5 port map( A => B(1), B => n112, C => n113, D => n405,
                           E => n114, Z => n111);
   U60 : HS65_LH_AND2X4 port map( A => n113, B => n405, Z => n112);
   U61 : HS65_LH_NOR2AX3 port map( A => B(0), B => A(0), Z => n113);
   U62 : HS65_LH_OAI212X5 port map( A => A(12), B => n370, C => A(13), D => 
                           n371, E => n97, Z => n96);
   U63 : HS65_LH_NAND3X5 port map( A => n47, B => n54, C => n98, Z => n97);
   U64 : HS65_LH_OAI21X3 port map( A => A(11), B => n369, C => n99, Z => n98);
   U65 : HS65_LH_AOI32X5 port map( A => n53, B => n52, C => n100, D => B(10), E
                           => n399, Z => n99);
   U66 : HS65_LH_OAI212X5 port map( A => A(28), B => n380, C => A(29), D => 
                           n381, E => n81, Z => n80);
   U67 : HS65_LH_NAND3X5 port map( A => n61, B => n67, C => n82, Z => n81);
   U68 : HS65_LH_OAI21X3 port map( A => A(27), B => n379, C => n83, Z => n82);
   U69 : HS65_LH_AOI32X5 port map( A => n66, B => n65, C => n84, D => B(26), E 
                           => n385, Z => n83);
   U70 : HS65_LH_AOI32X5 port map( A => n73, B => n75, C => n88, D => B(22), E 
                           => n393, Z => n87);
   U71 : HS65_LH_IVX9 port map( A => A(22), Z => n393);
   U72 : HS65_LH_OAI212X5 port map( A => A(20), B => n375, C => A(21), D => 
                           n376, E => n89, Z => n88);
   U73 : HS65_LH_NAND3X5 port map( A => n74, B => n68, C => n90, Z => n89);
   U74 : HS65_LH_AOI32X5 port map( A => n396, B => n49, C => n94, D => B(16), E
                           => n397, Z => n93);
   U75 : HS65_LH_IVX9 port map( A => n71, Z => n396);
   U76 : HS65_LH_OAI21X3 port map( A => A(15), B => n372, C => n95, Z => n94);
   U77 : HS65_LH_AOI32X5 port map( A => n50, B => n48, C => n96, D => B(14), E 
                           => n384, Z => n95);
   U78 : HS65_LH_AOI32X5 port map( A => n105, B => n106, C => n107, D => B(6), 
                           E => n402, Z => n104);
   U79 : HS65_LH_IVX9 port map( A => A(6), Z => n402);
   U80 : HS65_LH_OAI21X3 port map( A => A(5), B => n366, C => n108, Z => n107);
   U81 : HS65_LH_AOI32X5 port map( A => n403, B => n109, C => n110, D => B(4), 
                           E => n404, Z => n108);
   U82 : HS65_LH_AOI22X6 port map( A => n405, B => n63, C => n63, D => B(1), Z 
                           => n59);
   U83 : HS65_LH_NAND2AX7 port map( A => B(0), B => A(0), Z => n63);
   U84 : HS65_LH_OAI21X3 port map( A => A(25), B => n378, C => n85, Z => n84);
   U85 : HS65_LH_AOI32X5 port map( A => n391, B => n72, C => n86, D => B(24), E
                           => n392, Z => n85);
   U86 : HS65_LH_IVX9 port map( A => n64, Z => n391);
   U87 : HS65_LH_OAI21X3 port map( A => A(23), B => n377, C => n87, Z => n86);
   U88 : HS65_LH_OAI21X3 port map( A => A(9), B => n368, C => n101, Z => n100);
   U89 : HS65_LH_AOI32X5 port map( A => n400, B => n102, C => n103, D => B(8), 
                           E => n383, Z => n101);
   U90 : HS65_LH_IVX9 port map( A => n51, Z => n400);
   U91 : HS65_LH_OAI21X3 port map( A => A(7), B => n367, C => n104, Z => n103);
   U92 : HS65_LH_OAI21X3 port map( A => A(19), B => n374, C => n91, Z => n90);
   U93 : HS65_LH_AOI32X5 port map( A => n394, B => n69, C => n92, D => B(18), E
                           => n395, Z => n91);
   U94 : HS65_LH_IVX9 port map( A => n70, Z => n394);
   U95 : HS65_LH_OAI21X3 port map( A => A(17), B => n373, C => n93, Z => n92);
   U96 : HS65_LH_NAND2AX7 port map( A => B(6), B => A(6), Z => n105);
   U97 : HS65_LH_NAND2AX7 port map( A => B(10), B => A(10), Z => n53);
   U98 : HS65_LH_NAND2AX7 port map( A => B(22), B => A(22), Z => n73);
   U99 : HS65_LH_NAND2X7 port map( A => A(28), B => n380, Z => n61);
   U100 : HS65_LH_NAND2X7 port map( A => A(25), B => n378, Z => n65);
   U101 : HS65_LH_NAND2X7 port map( A => A(9), B => n368, Z => n52);
   U102 : HS65_LH_NAND2X7 port map( A => A(27), B => n379, Z => n67);
   U103 : HS65_LH_NAND2X7 port map( A => A(7), B => n367, Z => n102);
   U104 : HS65_LH_NAND2X7 port map( A => A(19), B => n374, Z => n68);
   U105 : HS65_LH_NAND2X7 port map( A => A(3), B => n365, Z => n109);
   U106 : HS65_LH_NAND2X7 port map( A => A(21), B => n376, Z => n75);
   U107 : HS65_LH_NAND2X7 port map( A => A(31), B => n382, Z => n76);
   U108 : HS65_LH_NAND2X7 port map( A => A(12), B => n370, Z => n47);
   U109 : HS65_LH_NAND2X7 port map( A => A(13), B => n371, Z => n48);
   U110 : HS65_LH_NAND2X7 port map( A => A(15), B => n372, Z => n49);
   U111 : HS65_LH_IVX9 port map( A => A(1), Z => n405);
   U112 : HS65_LH_IVX9 port map( A => A(4), Z => n404);
   U113 : HS65_LH_IVX9 port map( A => A(16), Z => n397);
   U114 : HS65_LH_IVX9 port map( A => A(24), Z => n392);
   U115 : HS65_LH_IVX9 port map( A => A(30), Z => n389);
   U116 : HS65_LH_IVX9 port map( A => A(18), Z => n395);
   U117 : HS65_LH_IVX9 port map( A => A(10), Z => n399);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_sub_0;

architecture SYN_rpl of alu_DW01_sub_0 is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n223, n224, n225,
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253 : std_logic;

begin
   
   U2_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => n252, CI => carry_30_port
                           , CO => carry_31_port, S0 => DIFF(30));
   U2_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => n250, CI => carry_28_port
                           , CO => carry_29_port, S0 => DIFF(28));
   U2_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => n249, CI => carry_27_port
                           , CO => carry_28_port, S0 => DIFF(27));
   U2_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => n244, CI => carry_22_port
                           , CO => carry_23_port, S0 => DIFF(22));
   U2_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => n241, CI => carry_19_port
                           , CO => carry_20_port, S0 => DIFF(19));
   U2_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => n240, CI => carry_18_port
                           , CO => carry_19_port, S0 => DIFF(18));
   U2_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => n238, CI => carry_16_port
                           , CO => carry_17_port, S0 => DIFF(16));
   U2_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => n237, CI => carry_15_port
                           , CO => carry_16_port, S0 => DIFF(15));
   U2_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => n235, CI => carry_13_port
                           , CO => carry_14_port, S0 => DIFF(13));
   U2_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => n234, CI => carry_12_port
                           , CO => carry_13_port, S0 => DIFF(12));
   U2_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => n232, CI => carry_10_port
                           , CO => carry_11_port, S0 => DIFF(10));
   U2_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => n231, CI => carry_9_port, 
                           CO => carry_10_port, S0 => DIFF(9));
   U2_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => n229, CI => carry_7_port, 
                           CO => carry_8_port, S0 => DIFF(7));
   U2_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => n228, CI => carry_6_port, 
                           CO => carry_7_port, S0 => DIFF(6));
   U2_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => n226, CI => carry_4_port, 
                           CO => carry_5_port, S0 => DIFF(4));
   U2_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => n225, CI => carry_3_port, 
                           CO => carry_4_port, S0 => DIFF(3));
   U2_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => n247, CI => carry_25_port
                           , CO => carry_26_port, S0 => DIFF(25));
   U2_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => n243, CI => carry_21_port
                           , CO => carry_22_port, S0 => DIFF(21));
   U2_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => n223, CI => carry_1_port, 
                           CO => carry_2_port, S0 => DIFF(1));
   U2_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => n246, CI => carry_24_port
                           , CO => carry_25_port, S0 => DIFF(24));
   U2_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => n224, CI => carry_2_port, 
                           CO => carry_3_port, S0 => DIFF(2));
   U2_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => n245, CI => carry_23_port
                           , CO => carry_24_port, S0 => DIFF(23));
   U2_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => n248, CI => carry_26_port
                           , CO => carry_27_port, S0 => DIFF(26));
   U2_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => n242, CI => carry_20_port
                           , CO => carry_21_port, S0 => DIFF(20));
   U2_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => n251, CI => carry_29_port
                           , CO => carry_30_port, S0 => DIFF(29));
   U2_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => n239, CI => carry_17_port
                           , CO => carry_18_port, S0 => DIFF(17));
   U2_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => n233, CI => carry_11_port
                           , CO => carry_12_port, S0 => DIFF(11));
   U2_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => n227, CI => carry_5_port, 
                           CO => carry_6_port, S0 => DIFF(5));
   U2_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => n236, CI => carry_14_port
                           , CO => carry_15_port, S0 => DIFF(14));
   U2_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => n230, CI => carry_8_port, 
                           CO => carry_9_port, S0 => DIFF(8));
   U1 : HS65_LH_IVX9 port map( A => B(8), Z => n230);
   U2 : HS65_LH_IVX9 port map( A => B(14), Z => n236);
   U3 : HS65_LH_IVX9 port map( A => B(5), Z => n227);
   U4 : HS65_LH_IVX9 port map( A => B(11), Z => n233);
   U5 : HS65_LH_IVX9 port map( A => B(17), Z => n239);
   U6 : HS65_LH_IVX9 port map( A => B(29), Z => n251);
   U7 : HS65_LH_IVX9 port map( A => B(20), Z => n242);
   U8 : HS65_LH_IVX9 port map( A => B(26), Z => n248);
   U9 : HS65_LH_IVX9 port map( A => B(23), Z => n245);
   U10 : HS65_LH_IVX9 port map( A => B(2), Z => n224);
   U11 : HS65_LHS_XNOR3X2 port map( A => A(31), B => B(31), C => carry_31_port,
                           Z => DIFF(31));
   U12 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => DIFF(0));
   U13 : HS65_LH_IVX9 port map( A => B(24), Z => n246);
   U14 : HS65_LH_IVX9 port map( A => B(1), Z => n223);
   U15 : HS65_LH_NAND2X7 port map( A => n253, B => B(0), Z => carry_1_port);
   U16 : HS65_LH_IVX9 port map( A => A(0), Z => n253);
   U17 : HS65_LH_IVX9 port map( A => B(21), Z => n243);
   U18 : HS65_LH_IVX9 port map( A => B(25), Z => n247);
   U19 : HS65_LH_IVX9 port map( A => B(3), Z => n225);
   U20 : HS65_LH_IVX9 port map( A => B(4), Z => n226);
   U21 : HS65_LH_IVX9 port map( A => B(6), Z => n228);
   U22 : HS65_LH_IVX9 port map( A => B(7), Z => n229);
   U23 : HS65_LH_IVX9 port map( A => B(9), Z => n231);
   U24 : HS65_LH_IVX9 port map( A => B(10), Z => n232);
   U25 : HS65_LH_IVX9 port map( A => B(12), Z => n234);
   U26 : HS65_LH_IVX9 port map( A => B(13), Z => n235);
   U27 : HS65_LH_IVX9 port map( A => B(15), Z => n237);
   U28 : HS65_LH_IVX9 port map( A => B(16), Z => n238);
   U29 : HS65_LH_IVX9 port map( A => B(18), Z => n240);
   U30 : HS65_LH_IVX9 port map( A => B(19), Z => n241);
   U31 : HS65_LH_IVX9 port map( A => B(22), Z => n244);
   U32 : HS65_LH_IVX9 port map( A => B(27), Z => n249);
   U33 : HS65_LH_IVX9 port map( A => B(28), Z => n250);
   U34 : HS65_LH_IVX9 port map( A => B(30), Z => n252);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_cmp_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in 
         std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);

end alu_DW_cmp_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_cmp_0 is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND3X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2AX7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3AX6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI312X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA112X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI211X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   signal n226, n227, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
      n327, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621 : std_logic;

begin
   
   U157 : HS65_LH_AND2X4 port map( A => A(23), B => n587, Z => n284);
   U158 : HS65_LH_IVX9 port map( A => B(1), Z => n580);
   U159 : HS65_LH_OR2X9 port map( A => B(29), B => n599, Z => n294);
   U160 : HS65_LH_IVX9 port map( A => B(2), Z => n581);
   U161 : HS65_LH_IVX9 port map( A => B(23), Z => n587);
   U162 : HS65_LH_IVX9 port map( A => B(3), Z => n582);
   U163 : HS65_LH_IVX9 port map( A => B(22), Z => n586);
   U164 : HS65_LH_IVX9 port map( A => B(30), Z => n592);
   U165 : HS65_LH_IVX9 port map( A => A(14), Z => n596);
   U166 : HS65_LH_IVX9 port map( A => n304, Z => n609);
   U167 : HS65_LH_IVX9 port map( A => A(8), Z => n594);
   U168 : HS65_LH_IVX9 port map( A => A(5), Z => n593);
   U169 : HS65_LH_IVX9 port map( A => A(17), Z => n597);
   U170 : HS65_LH_IVX9 port map( A => A(29), Z => n599);
   U171 : HS65_LH_IVX9 port map( A => A(20), Z => n598);
   U172 : HS65_LH_IVX9 port map( A => A(11), Z => n595);
   U173 : HS65_LH_OAI32X5 port map( A => n273, B => n274, C => n275, D => n276,
                           E => n273, Z => n272);
   U174 : HS65_LH_OA22X9 port map( A => n226, B => n227, C => n227, D => n283, 
                           Z => n274);
   U175 : HS65_LH_CBI4I1X5 port map( A => n600, B => n601, C => n286, D => n287
                           , Z => n273);
   U176 : HS65_LH_AOI212X4 port map( A => n277, B => n278, C => n278, D => n605
                           , E => n279, Z => n275);
   U177 : HS65_LH_OAI21X3 port map( A => n270, B => n271, C => n272, Z => 
                           GE_LT_GT_LE);
   U178 : HS65_LH_AOI312X4 port map( A => n294, B => n603, C => B(28), D => 
                           B(29), E => n599, F => n295, Z => n286);
   U179 : HS65_LH_OAI212X5 port map( A => n299, B => n300, C => n301, D => n299
                           , E => n302, Z => n270);
   U180 : HS65_LH_OA12X9 port map( A => n606, B => B(16), C => n282, Z => n302)
                           ;
   U181 : HS65_LH_CBI4I1X5 port map( A => n307, B => n308, C => n309, D => n310
                           , Z => n300);
   U182 : HS65_LH_NOR3X4 port map( A => n303, B => n304, C => n305, Z => n301);
   U183 : HS65_LH_CBI4I1X5 port map( A => n319, B => n320, C => n321, D => n322
                           , Z => n299);
   U184 : HS65_LH_OAI212X5 port map( A => n323, B => n324, C => n613, D => n323
                           , E => n609, Z => n322);
   U185 : HS65_LH_AOI312X4 port map( A => n325, B => n612, C => B(12), D => 
                           B(13), E => n611, F => n607, Z => n321);
   U186 : HS65_LH_IVX9 port map( A => n305, Z => n613);
   U187 : HS65_LH_OAI211X5 port map( A => B(12), B => n612, C => n325, D => 
                           n610, Z => n304);
   U188 : HS65_LH_IVX9 port map( A => n320, Z => n610);
   U189 : HS65_LH_AOI32X5 port map( A => n282, B => n606, C => B(16), D => 
                           B(17), E => n597, Z => n277);
   U190 : HS65_LH_AOI12X2 port map( A => n590, B => A(26), C => n293, Z => n290
                           );
   U191 : HS65_LH_OAI21X3 port map( A => B(14), B => n596, C => n327, Z => n320
                           );
   U192 : HS65_LH_OAI211X5 port map( A => B(20), B => n598, C => n285, D => 
                           n283, Z => n279);
   U193 : HS65_LH_OAI21X3 port map( A => B(10), B => n614, C => n326, Z => n305
                           );
   U194 : HS65_LH_OAI21X3 port map( A => B(6), B => n618, C => n318, Z => n308)
                           ;
   U195 : HS65_LH_NOR2X6 port map( A => n593, B => B(5), Z => n315);
   U196 : HS65_LH_NAND3AX6 port map( A => n279, B => n280, C => n276, Z => n271
                           );
   U197 : HS65_LH_OA112X9 port map( A => B(28), B => n603, C => n294, D => n296
                           , Z => n291);
   U198 : HS65_LH_OAI21X3 port map( A => B(8), B => n594, C => n306, Z => n303)
                           ;
   U199 : HS65_LH_AO32X4 port map( A => B(10), B => n614, C => n326, D => n595,
                           E => B(11), Z => n323);
   U200 : HS65_LH_OR2X9 port map( A => B(13), B => n611, Z => n325);
   U201 : HS65_LH_IVX9 port map( A => n295, Z => n600);
   U202 : HS65_LH_AND2X4 port map( A => B(31), B => n602, Z => n297);
   U203 : HS65_LH_OR2X9 port map( A => B(17), B => n597, Z => n282);
   U204 : HS65_LH_OR2X9 port map( A => B(21), B => n604, Z => n285);
   U205 : HS65_LH_AO32X4 port map( A => n285, B => n598, C => B(20), D => B(21)
                           , E => n604, Z => n226);
   U206 : HS65_LH_OR2X9 port map( A => B(11), B => n595, Z => n326);
   U207 : HS65_LH_IVX9 port map( A => B(4), Z => n583);
   U208 : HS65_LH_IVX9 port map( A => n319, Z => n607);
   U209 : HS65_LH_IVX9 port map( A => n307, Z => n616);
   U210 : HS65_LH_IVX9 port map( A => B(27), Z => n591);
   U211 : HS65_LH_IVX9 port map( A => B(26), Z => n590);
   U212 : HS65_LH_IVX9 port map( A => B(24), Z => n588);
   U213 : HS65_LH_IVX9 port map( A => B(19), Z => n585);
   U214 : HS65_LH_IVX9 port map( A => B(18), Z => n584);
   U215 : HS65_LH_IVX9 port map( A => n280, Z => n605);
   U216 : HS65_LH_IVX9 port map( A => n296, Z => n601);
   U217 : HS65_LH_OAI32X5 port map( A => n592, B => A(30), C => n297, D => 
                           B(31), E => n602, Z => n295);
   U218 : HS65_LH_OAI32X5 port map( A => n586, B => A(22), C => n284, D => 
                           A(23), E => n587, Z => n227);
   U219 : HS65_LH_AOI312X4 port map( A => n619, B => n620, C => B(4), D => B(5)
                           , E => n593, F => n616, Z => n309);
   U220 : HS65_LH_IVX9 port map( A => A(4), Z => n620);
   U221 : HS65_LH_IVX9 port map( A => n315, Z => n619);
   U222 : HS65_LH_OAI212X5 port map( A => n288, B => n289, C => n290, D => n288
                           , E => n291, Z => n287);
   U223 : HS65_LH_OAI32X5 port map( A => n588, B => A(24), C => n292, D => 
                           A(25), E => n589, Z => n289);
   U224 : HS65_LH_OAI32X5 port map( A => n590, B => A(26), C => n293, D => 
                           A(27), E => n591, Z => n288);
   U225 : HS65_LH_IVX9 port map( A => B(25), Z => n589);
   U226 : HS65_LH_AOI32X5 port map( A => B(14), B => n596, C => n327, D => n608
                           , E => B(15), Z => n319);
   U227 : HS65_LH_IVX9 port map( A => A(15), Z => n608);
   U228 : HS65_LH_AOI32X5 port map( A => B(6), B => n618, C => n318, D => n617,
                           E => B(7), Z => n307);
   U229 : HS65_LH_IVX9 port map( A => A(7), Z => n617);
   U230 : HS65_LH_AOI12X2 port map( A => n584, B => A(18), C => n281, Z => n280
                           );
   U231 : HS65_LH_AOI22X6 port map( A => B(1), B => n621, C => n316, D => B(0),
                           Z => n313);
   U232 : HS65_LH_IVX9 port map( A => A(1), Z => n621);
   U233 : HS65_LH_AOI12X2 port map( A => A(1), B => n580, C => A(0), Z => n316)
                           ;
   U234 : HS65_LH_AOI12X2 port map( A => n586, B => A(22), C => n284, Z => n283
                           );
   U235 : HS65_LH_NOR2AX3 port map( A => A(25), B => B(25), Z => n292);
   U236 : HS65_LH_NAND3AX6 port map( A => n308, B => n311, C => n312, Z => n310
                           );
   U237 : HS65_LH_CBI4I1X5 port map( A => A(2), B => n581, C => n317, D => n314
                           , Z => n311);
   U238 : HS65_LH_AOI212X4 port map( A => n313, B => n314, C => A(4), D => n583
                           , E => n315, Z => n312);
   U239 : HS65_LH_OA32X4 port map( A => n581, B => A(2), C => n317, D => A(3), 
                           E => n582, Z => n314);
   U240 : HS65_LH_AOI12X2 port map( A => n592, B => A(30), C => n297, Z => n296
                           );
   U241 : HS65_LH_OA32X4 port map( A => n584, B => A(18), C => n281, D => A(19)
                           , E => n585, Z => n278);
   U242 : HS65_LH_NAND2AX7 port map( A => B(15), B => A(15), Z => n327);
   U243 : HS65_LH_NAND2AX7 port map( A => B(7), B => A(7), Z => n318);
   U244 : HS65_LH_NAND2AX7 port map( A => B(9), B => A(9), Z => n306);
   U245 : HS65_LH_AND2X4 port map( A => A(27), B => n591, Z => n293);
   U246 : HS65_LH_AO32X4 port map( A => B(8), B => n594, C => n306, D => n615, 
                           E => B(9), Z => n324);
   U247 : HS65_LH_IVX9 port map( A => A(9), Z => n615);
   U248 : HS65_LH_AND3X9 port map( A => n290, B => n291, C => n298, Z => n276);
   U249 : HS65_LH_AOI12X2 port map( A => A(24), B => n588, C => n292, Z => n298
                           );
   U250 : HS65_LH_AND2X4 port map( A => A(3), B => n582, Z => n317);
   U251 : HS65_LH_AND2X4 port map( A => A(19), B => n585, Z => n281);
   U252 : HS65_LH_IVX9 port map( A => A(12), Z => n612);
   U253 : HS65_LH_IVX9 port map( A => A(6), Z => n618);
   U254 : HS65_LH_IVX9 port map( A => A(13), Z => n611);
   U255 : HS65_LH_IVX9 port map( A => A(16), Z => n606);
   U256 : HS65_LH_IVX9 port map( A => A(31), Z => n602);
   U257 : HS65_LH_IVX9 port map( A => A(10), Z => n614);
   U258 : HS65_LH_IVX9 port map( A => A(28), Z => n603);
   U259 : HS65_LH_IVX9 port map( A => A(21), Z => n604);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_ctrl is

   port( alu_ctrl_i : in std_logic_vector (9 downto 0);  alu_ctrl_o : out 
         std_logic_vector (4 downto 0));

end alu_ctrl;

architecture SYN_Behavioral of alu_ctrl is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3AX6
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI33X3
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI33X5
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI211X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI13X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125 : std_logic;

begin
   
   U3 : HS65_LH_NOR2X6 port map( A => n33, B => n116, Z => n22);
   U4 : HS65_LH_NOR2X6 port map( A => n124, B => n125, Z => n19);
   U5 : HS65_LH_AOI12X2 port map( A => n124, B => n125, C => n19, Z => n13);
   U6 : HS65_LH_NAND2X7 port map( A => n26, B => n22, Z => n16);
   U7 : HS65_LH_NAND2X7 port map( A => n118, B => n119, Z => n33);
   U8 : HS65_LH_NOR2X6 port map( A => n25, B => n123, Z => n23);
   U9 : HS65_LH_IVX9 port map( A => n24, Z => n116);
   U10 : HS65_LH_OAI212X5 port map( A => n16, B => n20, C => n12, D => n118, E 
                           => n21, Z => alu_ctrl_o(2));
   U11 : HS65_LH_OAI21X3 port map( A => alu_ctrl_i(1), B => n121, C => n125, Z 
                           => n20);
   U12 : HS65_LH_AOI13X5 port map( A => n13, B => n22, C => n23, D => n117, Z 
                           => n21);
   U13 : HS65_LH_IVX9 port map( A => n18, Z => n117);
   U14 : HS65_LH_OAI212X5 port map( A => alu_ctrl_i(9), B => n27, C => 
                           alu_ctrl_i(0), D => n17, E => n31, Z => 
                           alu_ctrl_o(0));
   U15 : HS65_LH_AOI32X5 port map( A => n22, B => n32, C => n120, D => n24, E 
                           => n33, Z => n31);
   U16 : HS65_LH_IVX9 port map( A => n25, Z => n120);
   U17 : HS65_LH_AO22X9 port map( A => n125, B => alu_ctrl_i(2), C => n123, D 
                           => n19, Z => n32);
   U18 : HS65_LH_OAI211X5 port map( A => n15, B => n16, C => n17, D => n18, Z 
                           => alu_ctrl_o(3));
   U19 : HS65_LH_AOI22X6 port map( A => n19, B => n121, C => alu_ctrl_i(4), D 
                           => n125, Z => n15);
   U20 : HS65_LH_OAI212X5 port map( A => alu_ctrl_i(9), B => n27, C => n125, D 
                           => n17, E => n28, Z => alu_ctrl_o(1));
   U21 : HS65_LH_AOI33X5 port map( A => n29, B => n124, C => n22, D => 
                           alu_ctrl_i(7), E => n24, F => alu_ctrl_i(8), Z => 
                           n28);
   U22 : HS65_LH_OAI33X3 port map( A => n30, B => alu_ctrl_i(5), C => 
                           alu_ctrl_i(2), D => n123, E => alu_ctrl_i(0), F => 
                           n25, Z => n29);
   U23 : HS65_LH_AOI32X5 port map( A => alu_ctrl_i(3), B => alu_ctrl_i(0), C =>
                           alu_ctrl_i(4), D => n125, E => n121, Z => n30);
   U24 : HS65_LH_NOR3X4 port map( A => alu_ctrl_i(3), B => alu_ctrl_i(5), C => 
                           alu_ctrl_i(2), Z => n26);
   U25 : HS65_LH_NAND4ABX3 port map( A => n122, B => n34, C => alu_ctrl_i(5), D
                           => n22, Z => n17);
   U26 : HS65_LH_NAND3X5 port map( A => n123, B => n121, C => alu_ctrl_i(1), Z 
                           => n34);
   U27 : HS65_LH_IVX9 port map( A => alu_ctrl_i(0), Z => n125);
   U28 : HS65_LH_NAND3X5 port map( A => n122, B => n121, C => alu_ctrl_i(5), Z 
                           => n25);
   U29 : HS65_LH_CBI4I1X5 port map( A => n118, B => n11, C => n116, D => n12, Z
                           => alu_ctrl_o(4));
   U30 : HS65_LH_NAND4ABX3 port map( A => n13, B => n14, C => n125, D => 
                           alu_ctrl_i(3), Z => n11);
   U31 : HS65_LH_NAND4ABX3 port map( A => alu_ctrl_i(2), B => alu_ctrl_i(5), C 
                           => n121, D => n119, Z => n14);
   U32 : HS65_LH_NOR2X6 port map( A => alu_ctrl_i(6), B => alu_ctrl_i(9), Z => 
                           n24);
   U33 : HS65_LH_NAND3AX6 port map( A => n33, B => n26, C => n35, Z => n27);
   U34 : HS65_LH_NOR3X4 port map( A => n36, B => alu_ctrl_i(6), C => 
                           alu_ctrl_i(0), Z => n35);
   U35 : HS65_LHS_XOR2X6 port map( A => alu_ctrl_i(4), B => n124, Z => n36);
   U36 : HS65_LH_IVX9 port map( A => alu_ctrl_i(4), Z => n121);
   U37 : HS65_LH_NAND3AX6 port map( A => alu_ctrl_i(9), B => alu_ctrl_i(6), C 
                           => alu_ctrl_i(7), Z => n12);
   U38 : HS65_LH_NAND3X5 port map( A => n24, B => n118, C => alu_ctrl_i(7), Z 
                           => n18);
   U39 : HS65_LH_IVX9 port map( A => alu_ctrl_i(1), Z => n124);
   U40 : HS65_LH_IVX9 port map( A => alu_ctrl_i(8), Z => n118);
   U41 : HS65_LH_IVX9 port map( A => alu_ctrl_i(2), Z => n123);
   U42 : HS65_LH_IVX9 port map( A => alu_ctrl_i(7), Z => n119);
   U43 : HS65_LH_IVX9 port map( A => alu_ctrl_i(3), Z => n122);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu is

   port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 0);
         alu_o : out std_logic_vector (32 downto 0));

end alu;

architecture SYN_behavioral of alu is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI222X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I6X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO312X9
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO33X9
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI33X5
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI222X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI13X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CB4I6X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component alu_DW_mult_uns_0
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component alu_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component alu_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW_cmp_0
      port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in
            std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal HI_LO_c_HI_31_port, HI_LO_c_HI_30_port, HI_LO_c_HI_29_port, 
      HI_LO_c_HI_28_port, HI_LO_c_HI_27_port, HI_LO_c_HI_26_port, 
      HI_LO_c_HI_25_port, HI_LO_c_HI_24_port, HI_LO_c_HI_23_port, 
      HI_LO_c_HI_22_port, HI_LO_c_HI_21_port, HI_LO_c_HI_20_port, 
      HI_LO_c_HI_19_port, HI_LO_c_HI_18_port, HI_LO_c_HI_17_port, 
      HI_LO_c_HI_16_port, HI_LO_c_HI_15_port, HI_LO_c_HI_14_port, 
      HI_LO_c_HI_13_port, HI_LO_c_HI_12_port, HI_LO_c_HI_11_port, 
      HI_LO_c_HI_10_port, HI_LO_c_HI_9_port, HI_LO_c_HI_8_port, 
      HI_LO_c_HI_7_port, HI_LO_c_HI_6_port, HI_LO_c_HI_5_port, 
      HI_LO_c_HI_4_port, HI_LO_c_HI_3_port, HI_LO_c_HI_2_port, 
      HI_LO_c_HI_1_port, HI_LO_c_HI_0_port, HI_LO_c_LO_31_port, 
      HI_LO_c_LO_30_port, HI_LO_c_LO_29_port, HI_LO_c_LO_28_port, 
      HI_LO_c_LO_27_port, HI_LO_c_LO_26_port, HI_LO_c_LO_25_port, 
      HI_LO_c_LO_24_port, HI_LO_c_LO_23_port, HI_LO_c_LO_22_port, 
      HI_LO_c_LO_21_port, HI_LO_c_LO_20_port, HI_LO_c_LO_19_port, 
      HI_LO_c_LO_18_port, HI_LO_c_LO_17_port, HI_LO_c_LO_16_port, 
      HI_LO_c_LO_15_port, HI_LO_c_LO_14_port, HI_LO_c_LO_13_port, 
      HI_LO_c_LO_12_port, HI_LO_c_LO_11_port, HI_LO_c_LO_10_port, 
      HI_LO_c_LO_9_port, HI_LO_c_LO_8_port, HI_LO_c_LO_7_port, 
      HI_LO_c_LO_6_port, HI_LO_c_LO_5_port, HI_LO_c_LO_4_port, 
      HI_LO_c_LO_3_port, HI_LO_c_LO_2_port, HI_LO_c_LO_1_port, 
      HI_LO_c_LO_0_port, N98, N99, N100, N101, N102, N103, N104, N105, N106, 
      N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, 
      N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, 
      N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, 
      N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, 
      N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, 
      N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, 
      N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
      N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
      N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
      N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N647, 
      N648, N713, N714, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n6, n7, n8, n9, n10, n86, n87, 
      n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98_port, n99_port, 
      n100_port, n101_port, n102_port, n103_port, n104_port, n105_port, 
      n106_port, n107_port, n108_port, n109_port, n110_port, n111_port, 
      n112_port, n113_port, n114_port, n115_port, n116_port, n117_port, 
      n118_port, n119_port, n120_port, n121_port, n122_port, n123_port, 
      n124_port, n125_port, n126_port, n127_port, n128_port, n129_port, 
      n130_port, n131_port, n132_port, n133_port, n134_port, n135_port, 
      n136_port, n137_port, n138_port, n139_port, n140_port, n141_port, 
      n142_port, n143_port, n144_port, n145_port, n146_port, n147_port, 
      n148_port, n149_port, n150_port, n151_port, n152_port, n153_port, 
      n154_port, n155_port, n156_port, n157_port, n158_port, n159_port, 
      n160_port, n161_port, n162_port, n163_port, n164_port, n165_port, 
      n166_port, n167_port, n168_port, n169_port, n170_port, n171_port, 
      n172_port, n173_port, n174_port, n175_port, n176_port, n177_port, 
      n178_port, n179_port, n180_port, n181_port, n182_port, n183_port, 
      n184_port, n185_port, n186_port, n187_port, n188_port, n189_port, 
      n190_port, n191_port, n192_port, n193_port, n194_port, n195_port, 
      n196_port, n197_port, n198_port, n199_port, n200_port, n201_port, 
      n202_port, n203_port, n204_port, n205_port, n206_port, n207_port, 
      n208_port, n209_port, n210_port, n211_port, n212_port, n213_port, 
      n214_port, n215_port, n216_port, n217_port, n218_port, n219_port, 
      n220_port, n221_port, n222_port, n223_port, n224_port, n225_port, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n_1014, n_1015, n_1016, n_1017, n_1018
      , n_1019 : std_logic;

begin
   
   HI_LO_c_reg_HI_31_inst : HS65_LH_DFPRQX9 port map( D => n525, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_31_port);
   HI_LO_c_reg_HI_30_inst : HS65_LH_DFPRQX9 port map( D => n524, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_30_port);
   HI_LO_c_reg_HI_29_inst : HS65_LH_DFPRQX9 port map( D => n523, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_29_port);
   HI_LO_c_reg_HI_28_inst : HS65_LH_DFPRQX9 port map( D => n522, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_28_port);
   HI_LO_c_reg_HI_27_inst : HS65_LH_DFPRQX9 port map( D => n521, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_27_port);
   HI_LO_c_reg_HI_26_inst : HS65_LH_DFPRQX9 port map( D => n520, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_26_port);
   HI_LO_c_reg_HI_25_inst : HS65_LH_DFPRQX9 port map( D => n519, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_25_port);
   HI_LO_c_reg_HI_24_inst : HS65_LH_DFPRQX9 port map( D => n518, CP => clk, RN 
                           => n1748, Q => HI_LO_c_HI_24_port);
   HI_LO_c_reg_HI_23_inst : HS65_LH_DFPRQX9 port map( D => n517, CP => clk, RN 
                           => n1748, Q => HI_LO_c_HI_23_port);
   HI_LO_c_reg_HI_22_inst : HS65_LH_DFPRQX9 port map( D => n516, CP => clk, RN 
                           => n1748, Q => HI_LO_c_HI_22_port);
   HI_LO_c_reg_HI_21_inst : HS65_LH_DFPRQX9 port map( D => n515, CP => clk, RN 
                           => n1748, Q => HI_LO_c_HI_21_port);
   HI_LO_c_reg_HI_20_inst : HS65_LH_DFPRQX9 port map( D => n514, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_20_port);
   HI_LO_c_reg_HI_19_inst : HS65_LH_DFPRQX9 port map( D => n513, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_19_port);
   HI_LO_c_reg_HI_18_inst : HS65_LH_DFPRQX9 port map( D => n512, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_18_port);
   HI_LO_c_reg_HI_17_inst : HS65_LH_DFPRQX9 port map( D => n511, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_17_port);
   HI_LO_c_reg_HI_16_inst : HS65_LH_DFPRQX9 port map( D => n510, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_16_port);
   HI_LO_c_reg_HI_15_inst : HS65_LH_DFPRQX9 port map( D => n509, CP => clk, RN 
                           => n1747, Q => HI_LO_c_HI_15_port);
   HI_LO_c_reg_HI_14_inst : HS65_LH_DFPRQX9 port map( D => n508, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_14_port);
   HI_LO_c_reg_HI_13_inst : HS65_LH_DFPRQX9 port map( D => n507, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_13_port);
   HI_LO_c_reg_HI_12_inst : HS65_LH_DFPRQX9 port map( D => n506, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_12_port);
   HI_LO_c_reg_HI_11_inst : HS65_LH_DFPRQX9 port map( D => n505, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_11_port);
   HI_LO_c_reg_HI_10_inst : HS65_LH_DFPRQX9 port map( D => n504, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_10_port);
   HI_LO_c_reg_HI_9_inst : HS65_LH_DFPRQX9 port map( D => n503, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_9_port);
   HI_LO_c_reg_HI_8_inst : HS65_LH_DFPRQX9 port map( D => n502, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_8_port);
   HI_LO_c_reg_HI_7_inst : HS65_LH_DFPRQX9 port map( D => n501, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_7_port);
   HI_LO_c_reg_HI_6_inst : HS65_LH_DFPRQX9 port map( D => n500, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_6_port);
   HI_LO_c_reg_HI_5_inst : HS65_LH_DFPRQX9 port map( D => n499, CP => clk, RN 
                           => n1745, Q => HI_LO_c_HI_5_port);
   HI_LO_c_reg_HI_4_inst : HS65_LH_DFPRQX9 port map( D => n498, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_4_port);
   HI_LO_c_reg_HI_3_inst : HS65_LH_DFPRQX9 port map( D => n497, CP => clk, RN 
                           => n1746, Q => HI_LO_c_HI_3_port);
   HI_LO_c_reg_HI_2_inst : HS65_LH_DFPRQX9 port map( D => n496, CP => clk, RN 
                           => n1745, Q => HI_LO_c_HI_2_port);
   HI_LO_c_reg_HI_1_inst : HS65_LH_DFPRQX9 port map( D => n495, CP => clk, RN 
                           => n1745, Q => HI_LO_c_HI_1_port);
   HI_LO_c_reg_HI_0_inst : HS65_LH_DFPRQX9 port map( D => n494, CP => clk, RN 
                           => n1745, Q => HI_LO_c_HI_0_port);
   HI_LO_c_reg_LO_31_inst : HS65_LH_DFPRQX9 port map( D => n493, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_31_port);
   HI_LO_c_reg_LO_30_inst : HS65_LH_DFPRQX9 port map( D => n492, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_30_port);
   HI_LO_c_reg_LO_29_inst : HS65_LH_DFPRQX9 port map( D => n491, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_29_port);
   HI_LO_c_reg_LO_28_inst : HS65_LH_DFPRQX9 port map( D => n490, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_28_port);
   HI_LO_c_reg_LO_27_inst : HS65_LH_DFPRQX9 port map( D => n489, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_27_port);
   HI_LO_c_reg_LO_26_inst : HS65_LH_DFPRQX9 port map( D => n488, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_26_port);
   HI_LO_c_reg_LO_25_inst : HS65_LH_DFPRQX9 port map( D => n487, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_25_port);
   HI_LO_c_reg_LO_24_inst : HS65_LH_DFPRQX9 port map( D => n486, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_24_port);
   HI_LO_c_reg_LO_23_inst : HS65_LH_DFPRQX9 port map( D => n485, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_23_port);
   HI_LO_c_reg_LO_22_inst : HS65_LH_DFPRQX9 port map( D => n484, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_22_port);
   HI_LO_c_reg_LO_21_inst : HS65_LH_DFPRQX9 port map( D => n483, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_21_port);
   HI_LO_c_reg_LO_20_inst : HS65_LH_DFPRQX9 port map( D => n482, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_20_port);
   HI_LO_c_reg_LO_19_inst : HS65_LH_DFPRQX9 port map( D => n481, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_19_port);
   HI_LO_c_reg_LO_18_inst : HS65_LH_DFPRQX9 port map( D => n480, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_18_port);
   HI_LO_c_reg_LO_17_inst : HS65_LH_DFPRQX9 port map( D => n479, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_17_port);
   HI_LO_c_reg_LO_16_inst : HS65_LH_DFPRQX9 port map( D => n478, CP => clk, RN 
                           => n1744, Q => HI_LO_c_LO_16_port);
   HI_LO_c_reg_LO_15_inst : HS65_LH_DFPRQX9 port map( D => n477, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_15_port);
   HI_LO_c_reg_LO_14_inst : HS65_LH_DFPRQX9 port map( D => n476, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_14_port);
   HI_LO_c_reg_LO_13_inst : HS65_LH_DFPRQX9 port map( D => n475, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_13_port);
   HI_LO_c_reg_LO_12_inst : HS65_LH_DFPRQX9 port map( D => n474, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_12_port);
   HI_LO_c_reg_LO_11_inst : HS65_LH_DFPRQX9 port map( D => n473, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_11_port);
   HI_LO_c_reg_LO_10_inst : HS65_LH_DFPRQX9 port map( D => n472, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_10_port);
   HI_LO_c_reg_LO_9_inst : HS65_LH_DFPRQX9 port map( D => n471, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_9_port);
   HI_LO_c_reg_LO_8_inst : HS65_LH_DFPRQX9 port map( D => n470, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_8_port);
   HI_LO_c_reg_LO_7_inst : HS65_LH_DFPRQX9 port map( D => n469, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_7_port);
   HI_LO_c_reg_LO_6_inst : HS65_LH_DFPRQX9 port map( D => n468, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_6_port);
   HI_LO_c_reg_LO_5_inst : HS65_LH_DFPRQX9 port map( D => n467, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_5_port);
   HI_LO_c_reg_LO_4_inst : HS65_LH_DFPRQX9 port map( D => n466, CP => clk, RN 
                           => n1743, Q => HI_LO_c_LO_4_port);
   HI_LO_c_reg_LO_3_inst : HS65_LH_DFPRQX9 port map( D => n465, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_3_port);
   HI_LO_c_reg_LO_2_inst : HS65_LH_DFPRQX9 port map( D => n464, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_2_port);
   HI_LO_c_reg_LO_1_inst : HS65_LH_DFPRQX9 port map( D => n463, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_1_port);
   HI_LO_c_reg_LO_0_inst : HS65_LH_DFPRQX9 port map( D => n462, CP => clk, RN 
                           => n1745, Q => HI_LO_c_LO_0_port);
   n6 <= '0';
   n7 <= '0';
   n8 <= '0';
   n9 <= '1';
   n10 <= '0';
   lt_136 : alu_DW_cmp_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => n1731,
                           A(1) => alu_i(43), A(0) => alu_i(42), B(31) => 
                           alu_i(41), B(30) => alu_i(40), B(29) => alu_i(39), 
                           B(28) => n1727, B(27) => n1726, B(26) => n1725, 
                           B(25) => n1724, B(24) => n1723, B(23) => alu_i(33), 
                           B(22) => alu_i(32), B(21) => n1720, B(20) => n1719, 
                           B(19) => n1718, B(18) => n1717, B(17) => n1716, 
                           B(16) => n1715, B(15) => n1714, B(14) => n1713, 
                           B(13) => n1712, B(12) => n1711, B(11) => n1710, 
                           B(10) => n1709, B(9) => n1708, B(8) => n1707, B(7) 
                           => n1706, B(6) => n1705, B(5) => n1704, B(4) => 
                           n1703, B(3) => alu_i(13), B(2) => alu_i(12), B(1) =>
                           alu_i(11), B(0) => alu_i(10), TC => n9, GE_LT => n9,
                           GE_GT_EQ => n10, GE_LT_GT_LE => N647, EQ_NE => 
                           n_1014);
   sub_68 : alu_DW01_sub_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => n1731,
                           A(1) => alu_i(43), A(0) => alu_i(42), B(31) => 
                           alu_i(41), B(30) => alu_i(40), B(29) => alu_i(39), 
                           B(28) => n1727, B(27) => n1726, B(26) => n1725, 
                           B(25) => n1724, B(24) => n1723, B(23) => alu_i(33), 
                           B(22) => alu_i(32), B(21) => n1720, B(20) => n1719, 
                           B(19) => n1718, B(18) => n1717, B(17) => n1716, 
                           B(16) => n1715, B(15) => n1714, B(14) => n1713, 
                           B(13) => n1712, B(12) => n1711, B(11) => n1710, 
                           B(10) => n1709, B(9) => n1708, B(8) => n1707, B(7) 
                           => n1706, B(6) => n1705, B(5) => n1704, B(4) => 
                           n1703, B(3) => alu_i(13), B(2) => alu_i(12), B(1) =>
                           alu_i(11), B(0) => alu_i(10), CI => n6, DIFF(31) => 
                           N161, DIFF(30) => N160, DIFF(29) => N159, DIFF(28) 
                           => N158, DIFF(27) => N157, DIFF(26) => N156, 
                           DIFF(25) => N155, DIFF(24) => N154, DIFF(23) => N153
                           , DIFF(22) => N152, DIFF(21) => N151, DIFF(20) => 
                           N150, DIFF(19) => N149, DIFF(18) => N148, DIFF(17) 
                           => N147, DIFF(16) => N146, DIFF(15) => N145, 
                           DIFF(14) => N144, DIFF(13) => N143, DIFF(12) => N142
                           , DIFF(11) => N141, DIFF(10) => N140, DIFF(9) => 
                           N139, DIFF(8) => N138, DIFF(7) => N137, DIFF(6) => 
                           N136, DIFF(5) => N135, DIFF(4) => N134, DIFF(3) => 
                           N133, DIFF(2) => N132, DIFF(1) => N131, DIFF(0) => 
                           N130, CO => n_1015);
   r325 : alu_DW01_cmp6_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => n1731,
                           A(1) => alu_i(43), A(0) => alu_i(42), B(31) => 
                           alu_i(41), B(30) => alu_i(40), B(29) => alu_i(39), 
                           B(28) => n1727, B(27) => n1726, B(26) => n1725, 
                           B(25) => n1724, B(24) => n1723, B(23) => alu_i(33), 
                           B(22) => alu_i(32), B(21) => n1720, B(20) => n1719, 
                           B(19) => n1718, B(18) => n1717, B(17) => n1716, 
                           B(16) => n1715, B(15) => n1714, B(14) => n1713, 
                           B(13) => n1712, B(12) => n1711, B(11) => n1710, 
                           B(10) => n1709, B(9) => n1708, B(8) => n1707, B(7) 
                           => n1706, B(6) => n1705, B(5) => n1704, B(4) => 
                           n1703, B(3) => alu_i(13), B(2) => alu_i(12), B(1) =>
                           alu_i(11), B(0) => alu_i(10), TC => n7, LT => N648, 
                           GT => n_1016, EQ => N713, LE => n_1017, GE => n_1018
                           , NE => N714);
   r321 : alu_DW01_add_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => n1731,
                           A(1) => alu_i(43), A(0) => alu_i(42), B(31) => 
                           alu_i(41), B(30) => alu_i(40), B(29) => alu_i(39), 
                           B(28) => n1727, B(27) => n1726, B(26) => n1725, 
                           B(25) => n1724, B(24) => n1723, B(23) => alu_i(33), 
                           B(22) => alu_i(32), B(21) => n1720, B(20) => n1719, 
                           B(19) => n1718, B(18) => n1717, B(17) => n1716, 
                           B(16) => n1715, B(15) => n1714, B(14) => n1713, 
                           B(13) => n1712, B(12) => n1711, B(11) => n1710, 
                           B(10) => n1709, B(9) => n1708, B(8) => n1707, B(7) 
                           => n1706, B(6) => n1705, B(5) => n1704, B(4) => 
                           n1703, B(3) => alu_i(13), B(2) => alu_i(12), B(1) =>
                           alu_i(11), B(0) => alu_i(10), CI => n8, SUM(31) => 
                           N129, SUM(30) => N128, SUM(29) => N127, SUM(28) => 
                           N126, SUM(27) => N125, SUM(26) => N124, SUM(25) => 
                           N123, SUM(24) => N122, SUM(23) => N121, SUM(22) => 
                           N120, SUM(21) => N119, SUM(20) => N118, SUM(19) => 
                           N117, SUM(18) => N116, SUM(17) => N115, SUM(16) => 
                           N114, SUM(15) => N113, SUM(14) => N112, SUM(13) => 
                           N111, SUM(12) => N110, SUM(11) => N109, SUM(10) => 
                           N108, SUM(9) => N107, SUM(8) => N106, SUM(7) => N105
                           , SUM(6) => N104, SUM(5) => N103, SUM(4) => N102, 
                           SUM(3) => N101, SUM(2) => N100, SUM(1) => N99, 
                           SUM(0) => N98, CO => n_1019);
   mult_71 : alu_DW_mult_uns_0 port map( a(31) => alu_i(73), a(30) => alu_i(72)
                           , a(29) => alu_i(71), a(28) => alu_i(70), a(27) => 
                           alu_i(69), a(26) => alu_i(68), a(25) => alu_i(67), 
                           a(24) => alu_i(66), a(23) => alu_i(65), a(22) => 
                           alu_i(64), a(21) => alu_i(63), a(20) => alu_i(62), 
                           a(19) => alu_i(61), a(18) => alu_i(60), a(17) => 
                           alu_i(59), a(16) => alu_i(58), a(15) => alu_i(57), 
                           a(14) => alu_i(56), a(13) => alu_i(55), a(12) => 
                           alu_i(54), a(11) => alu_i(53), a(10) => alu_i(52), 
                           a(9) => alu_i(51), a(8) => alu_i(50), a(7) => 
                           alu_i(49), a(6) => alu_i(48), a(5) => alu_i(47), 
                           a(4) => alu_i(46), a(3) => alu_i(45), a(2) => n1731,
                           a(1) => alu_i(43), a(0) => alu_i(42), b(31) => 
                           alu_i(41), b(30) => alu_i(40), b(29) => alu_i(39), 
                           b(28) => n1727, b(27) => n1726, b(26) => n1725, 
                           b(25) => n1724, b(24) => n1723, b(23) => alu_i(33), 
                           b(22) => alu_i(32), b(21) => n1720, b(20) => n1719, 
                           b(19) => n1718, b(18) => n1717, b(17) => n1716, 
                           b(16) => n1715, b(15) => n1714, b(14) => n1713, 
                           b(13) => n1712, b(12) => n1711, b(11) => n1710, 
                           b(10) => n1709, b(9) => n1708, b(8) => n1707, b(7) 
                           => n1706, b(6) => n1705, b(5) => n1704, b(4) => 
                           n1703, b(3) => alu_i(13), b(2) => alu_i(12), b(1) =>
                           alu_i(11), b(0) => alu_i(10), product(63) => N225, 
                           product(62) => N224, product(61) => N223, 
                           product(60) => N222, product(59) => N221, 
                           product(58) => N220, product(57) => N219, 
                           product(56) => N218, product(55) => N217, 
                           product(54) => N216, product(53) => N215, 
                           product(52) => N214, product(51) => N213, 
                           product(50) => N212, product(49) => N211, 
                           product(48) => N210, product(47) => N209, 
                           product(46) => N208, product(45) => N207, 
                           product(44) => N206, product(43) => N205, 
                           product(42) => N204, product(41) => N203, 
                           product(40) => N202, product(39) => N201, 
                           product(38) => N200, product(37) => N199, 
                           product(36) => N198, product(35) => N197, 
                           product(34) => N196, product(33) => N195, 
                           product(32) => N194, product(31) => N193, 
                           product(30) => N192, product(29) => N191, 
                           product(28) => N190, product(27) => N189, 
                           product(26) => N188, product(25) => N187, 
                           product(24) => N186, product(23) => N185, 
                           product(22) => N184, product(21) => N183, 
                           product(20) => N182, product(19) => N181, 
                           product(18) => N180, product(17) => N179, 
                           product(16) => N178, product(15) => N177, 
                           product(14) => N176, product(13) => N175, 
                           product(12) => N174, product(11) => N173, 
                           product(10) => N172, product(9) => N171, product(8) 
                           => N170, product(7) => N169, product(6) => N168, 
                           product(5) => N167, product(4) => N166, product(3) 
                           => N165, product(2) => N164, product(1) => N163, 
                           product(0) => N162);
   U7 : HS65_LH_IVX9 port map( A => n421, Z => n1641);
   U8 : HS65_LH_IVX9 port map( A => n317, Z => n1642);
   U9 : HS65_LH_NAND4ABX3 port map( A => n87, B => n88, C => n89, D => n90, Z 
                           => n86);
   U10 : HS65_LH_BFX9 port map( A => alu_i(29), Z => n1718);
   U11 : HS65_LH_BFX9 port map( A => alu_i(37), Z => n1726);
   U12 : HS65_LH_BFX9 port map( A => alu_i(36), Z => n1725);
   U13 : HS65_LH_BFX9 port map( A => alu_i(20), Z => n1709);
   U14 : HS65_LH_BFX9 port map( A => alu_i(22), Z => n1711);
   U15 : HS65_LH_BFX9 port map( A => alu_i(23), Z => n1712);
   U16 : HS65_LH_BFX9 port map( A => alu_i(24), Z => n1713);
   U17 : HS65_LH_BFX9 port map( A => alu_i(26), Z => n1715);
   U18 : HS65_LH_BFX9 port map( A => alu_i(27), Z => n1716);
   U19 : HS65_LH_BFX9 port map( A => alu_i(28), Z => n1717);
   U20 : HS65_LH_BFX9 port map( A => alu_i(30), Z => n1719);
   U21 : HS65_LH_BFX9 port map( A => alu_i(31), Z => n1720);
   U22 : HS65_LH_BFX9 port map( A => alu_i(34), Z => n1723);
   U23 : HS65_LH_BFX9 port map( A => alu_i(35), Z => n1724);
   U24 : HS65_LH_BFX9 port map( A => alu_i(21), Z => n1710);
   U25 : HS65_LH_BFX9 port map( A => alu_i(38), Z => n1727);
   U26 : HS65_LH_BFX9 port map( A => alu_i(25), Z => n1714);
   U27 : HS65_LH_BFX9 port map( A => alu_i(14), Z => n1703);
   U28 : HS65_LH_BFX9 port map( A => alu_i(16), Z => n1705);
   U29 : HS65_LH_BFX9 port map( A => alu_i(17), Z => n1706);
   U30 : HS65_LH_BFX9 port map( A => alu_i(15), Z => n1704);
   U31 : HS65_LH_BFX9 port map( A => alu_i(18), Z => n1707);
   U32 : HS65_LH_BFX9 port map( A => alu_i(19), Z => n1708);
   U33 : HS65_LH_IVX9 port map( A => n1686, Z => n1685);
   U34 : HS65_LH_IVX9 port map( A => n1686, Z => n1684);
   U35 : HS65_LH_IVX9 port map( A => n1694, Z => n1689);
   U36 : HS65_LH_IVX9 port map( A => n1694, Z => n1690);
   U37 : HS65_LH_IVX9 port map( A => n1694, Z => n1691);
   U38 : HS65_LH_IVX9 port map( A => n1693, Z => n1692);
   U39 : HS65_LH_AOI12X2 port map( A => n1651, B => n1642, C => n1682, Z => 
                           n235);
   U40 : HS65_LH_AOI12X2 port map( A => n1651, B => n1641, C => n1682, Z => 
                           n206_port);
   U41 : HS65_LH_IVX9 port map( A => n421, Z => n1751);
   U42 : HS65_LH_IVX9 port map( A => n317, Z => n1749);
   U43 : HS65_LH_IVX9 port map( A => n1682, Z => n1680);
   U44 : HS65_LH_IVX9 port map( A => n1682, Z => n1681);
   U45 : HS65_LH_BFX9 port map( A => n1687, Z => n1694);
   U46 : HS65_LH_BFX9 port map( A => n1687, Z => n1693);
   U47 : HS65_LH_BFX9 port map( A => n1793, Z => n1663);
   U48 : HS65_LH_BFX9 port map( A => n1793, Z => n1662);
   U49 : HS65_LH_BFX9 port map( A => n1795, Z => n1665);
   U50 : HS65_LH_BFX9 port map( A => n1792, Z => n1660);
   U51 : HS65_LH_BFX9 port map( A => n1792, Z => n1661);
   U52 : HS65_LH_IVX9 port map( A => n1683, Z => n1686);
   U53 : HS65_LH_BFX9 port map( A => n1687, Z => n1695);
   U54 : HS65_LH_BFX9 port map( A => n1688, Z => n1696);
   U55 : HS65_LH_BFX9 port map( A => n1688, Z => n1697);
   U56 : HS65_LH_BFX9 port map( A => n1795, Z => n1666);
   U57 : HS65_LH_BFX9 port map( A => n1793, Z => n1664);
   U58 : HS65_LH_BFX9 port map( A => n1688, Z => n1698);
   U59 : HS65_LH_IVX9 port map( A => n94, Z => n1793);
   U60 : HS65_LH_IVX9 port map( A => n96, Z => n1792);
   U61 : HS65_LH_IVX9 port map( A => n91, Z => n1795);
   U62 : HS65_LH_AND2X4 port map( A => n379, B => n1799, Z => n211_port);
   U63 : HS65_LH_NAND2X7 port map( A => n1752, B => n1756, Z => n421);
   U64 : HS65_LH_NOR2AX3 port map( A => n1670, B => n421, Z => n204_port);
   U65 : HS65_LH_NAND2X7 port map( A => n1750, B => n1756, Z => n317);
   U66 : HS65_LH_NOR4ABX2 port map( A => n91, B => n92, C => n1672, D => n93, Z
                           => n90);
   U67 : HS65_LH_NAND3X5 port map( A => n94, B => n1679, C => n96, Z => n93);
   U68 : HS65_LH_BFX9 port map( A => n92, Z => n1683);
   U69 : HS65_LH_NAND2X7 port map( A => n97, B => n1799, Z => n92);
   U70 : HS65_LH_IVX9 port map( A => n1672, Z => n1671);
   U71 : HS65_LH_IVX9 port map( A => n119_port, Z => n1672);
   U72 : HS65_LH_BFX9 port map( A => n98_port, Z => n1677);
   U73 : HS65_LH_BFX9 port map( A => n1768, Z => n1651);
   U74 : HS65_LH_IVX9 port map( A => n1679, Z => n1682);
   U75 : HS65_LH_BFX9 port map( A => n1768, Z => n1652);
   U76 : HS65_LH_IVX9 port map( A => n101_port, Z => n1798);
   U77 : HS65_LH_BFX9 port map( A => n98_port, Z => n1678);
   U78 : HS65_LH_BFX9 port map( A => n86, Z => n1687);
   U79 : HS65_LH_BFX9 port map( A => n86, Z => n1688);
   U80 : HS65_LH_BFX9 port map( A => n1768, Z => n1653);
   U81 : HS65_LH_BFX9 port map( A => n1654, Z => n1656);
   U82 : HS65_LH_BFX9 port map( A => n1655, Z => n1658);
   U83 : HS65_LH_BFX9 port map( A => n1654, Z => n1657);
   U84 : HS65_LH_BFX9 port map( A => n1655, Z => n1659);
   U85 : HS65_LH_CB4I6X9 port map( A => n1799, B => n99_port, C => n1794, D => 
                           n1676, Z => n88);
   U86 : HS65_LH_AOI13X5 port map( A => n101_port, B => n102_port, C => 
                           n103_port, D => n1796, Z => n87);
   U87 : HS65_LH_AOI12X2 port map( A => n97, B => n1798, C => n1677, Z => n89);
   U88 : HS65_LH_NAND3X5 port map( A => n432, B => n1801, C => n433, Z => 
                           n119_port);
   U89 : HS65_LH_IVX9 port map( A => n396, Z => n1768);
   U90 : HS65_LH_NOR2X6 port map( A => n1801, B => n1797, Z => n97);
   U91 : HS65_LH_AO32X4 port map( A => n104_port, B => n1801, C => n432, D => 
                           n1798, E => n379, Z => n98_port);
   U92 : HS65_LH_AOI222X2 port map( A => n1751, B => n194_port, C => n111_port,
                           D => n130_port, E => n1643, F => n131_port, Z => 
                           n185_port);
   U93 : HS65_LH_AOI222X2 port map( A => n109_port, B => n110_port, C => 
                           n111_port, D => n112_port, E => n1644, F => 
                           n114_port, Z => n108_port);
   U94 : HS65_LH_AOI222X2 port map( A => n275, B => n182_port, C => n214_port, 
                           D => n181_port, E => n211_port, F => alu_i(11), Z =>
                           n368);
   U95 : HS65_LH_AOI222X2 port map( A => n275, B => n160_port, C => n214_port, 
                           D => n161_port, E => n211_port, F => alu_i(12), Z =>
                           n361);
   U96 : HS65_LH_AOI222X2 port map( A => n275, B => n144_port, C => n214_port, 
                           D => n142_port, E => n211_port, F => alu_i(13), Z =>
                           n354);
   U97 : HS65_LH_AOI222X2 port map( A => n1754, B => n241, C => n1643, D => 
                           n166_port, E => alu_i(13), F => n200_port, Z => n240
                           );
   U98 : HS65_LH_AOI222X2 port map( A => n111_port, B => n114_port, C => n1751,
                           D => n177_port, E => n122_port, F => n112_port, Z =>
                           n176_port);
   U99 : HS65_LH_AOI212X4 port map( A => n120_port, B => n168_port, C => n1751,
                           D => n171_port, E => n420, Z => n415);
   U100 : HS65_LH_AO22X9 port map( A => n160_port, B => n212_port, C => 
                           n172_port, D => n111_port, Z => n420);
   U101 : HS65_LH_AOI212X4 port map( A => n273, B => n142_port, C => n212_port,
                           D => n215_port, E => n274, Z => n268);
   U102 : HS65_LH_AO22X9 port map( A => n213_port, B => n145_port, C => 
                           n216_port, D => n1749, Z => n274);
   U103 : HS65_LH_AOI212X4 port map( A => n145_port, B => n160_port, C => n1749
                           , D => n161_port, E => n162_port, Z => n159_port);
   U104 : HS65_LH_AO22X9 port map( A => n163_port, B => n120_port, C => 
                           n164_port, D => n109_port, Z => n162_port);
   U105 : HS65_LH_AOI212X4 port map( A => n120_port, B => n141_port, C => n1749
                           , D => n142_port, E => n143_port, Z => n140_port);
   U106 : HS65_LH_AO22X9 port map( A => n144_port, B => n1645, C => n146_port, 
                           D => n113_port, Z => n143_port);
   U107 : HS65_LH_IVX9 port map( A => n434, Z => n1752);
   U108 : HS65_LH_IVX9 port map( A => n190_port, Z => n1750);
   U109 : HS65_LH_AND2X4 port map( A => n364, B => n1750, Z => n214_port);
   U110 : HS65_LH_MX41X7 port map( D0 => alu_i(13), S0 => n1652, D1 => 
                           alu_i(12), S1 => n1649, D2 => n1656, S2 => alu_i(11)
                           , D3 => n1668, S3 => alu_i(10), Z => n144_port);
   U111 : HS65_LH_NAND3X5 port map( A => n1794, B => n1801, C => n104_port, Z 
                           => n96);
   U112 : HS65_LH_AND2X4 port map( A => n364, B => n1752, Z => n122_port);
   U113 : HS65_LH_NOR2X6 port map( A => n1801, B => n427, Z => n379);
   U114 : HS65_LH_NAND3X5 port map( A => n433, B => n1801, C => n1794, Z => n94
                           );
   U115 : HS65_LH_NOR2X6 port map( A => n433, B => n99_port, Z => n101_port);
   U116 : HS65_LH_IVX9 port map( A => n307, Z => n1756);
   U117 : HS65_LH_IVX9 port map( A => n102_port, Z => n1799);
   U118 : HS65_LH_MX41X7 port map( D0 => n1757, S0 => n164_port, D1 => n364, S1
                           => n168_port, D2 => n1756, S2 => n172_port, D3 => 
                           n1759, S3 => n163_port, Z => n241);
   U119 : HS65_LH_MX41X7 port map( D0 => n1757, S0 => n136_port, D1 => n1759, 
                           S1 => n132_port, D2 => n364, S2 => n129_port, D3 => 
                           n1756, S3 => n128_port, Z => n375);
   U120 : HS65_LH_MX41X7 port map( D0 => n1756, S0 => n297, D1 => n1757, S1 => 
                           n296, D2 => n1759, S2 => n181_port, D3 => n364, S3 
                           => n182_port, Z => n254);
   U121 : HS65_LH_NAND2X7 port map( A => n104_port, B => n379, Z => n91);
   U122 : HS65_LH_MX41X7 port map( D0 => n364, S0 => n144_port, D1 => n1757, S1
                           => n276, D2 => n1759, S2 => n142_port, D3 => n1756, 
                           S3 => n277, Z => n224_port);
   U123 : HS65_LH_MX41X7 port map( D0 => n364, S0 => n121_port, D1 => n1757, S1
                           => n123_port, D2 => n1759, S2 => n110_port, D3 => 
                           n1756, S3 => n112_port, Z => n350);
   U124 : HS65_LH_MX41X7 port map( D0 => n1757, S0 => n288, D1 => n364, S1 => 
                           n160_port, D2 => n1759, S2 => n161_port, D3 => n1756
                           , S3 => n283, Z => n236);
   U125 : HS65_LH_OAI21X3 port map( A => alu_i(39), B => n1685, C => n1680, Z 
                           => n253);
   U126 : HS65_LH_OAI21X3 port map( A => alu_i(40), B => n1685, C => n1680, Z 
                           => n234);
   U127 : HS65_LH_OAI21X3 port map( A => alu_i(41), B => n1685, C => n1680, Z 
                           => n219_port);
   U128 : HS65_LH_AO222X4 port map( A => n123_port, B => n1756, C => n110_port,
                           D => n1757, E => n121_port, F => n1759, Z => 
                           n178_port);
   U129 : HS65_LH_AO222X4 port map( A => n181_port, B => n1757, C => n182_port,
                           D => n1759, E => n296, F => n1756, Z => n116_port);
   U130 : HS65_LH_IVX9 port map( A => n427, Z => n1794);
   U131 : HS65_LH_BFX9 port map( A => n95, Z => n1679);
   U132 : HS65_LH_NAND2X7 port map( A => n97, B => n104_port, Z => n95);
   U133 : HS65_LH_IVX9 port map( A => n432, Z => n1797);
   U134 : HS65_LH_BFX9 port map( A => n1673, Z => n1674);
   U135 : HS65_LH_IVX9 port map( A => n343, Z => n1762);
   U136 : HS65_LH_BFX9 port map( A => n1673, Z => n1675);
   U137 : HS65_LH_BFX9 port map( A => n1770, Z => n1655);
   U138 : HS65_LH_BFX9 port map( A => n1770, Z => n1654);
   U139 : HS65_LH_BFX9 port map( A => n1667, Z => n1669);
   U140 : HS65_LH_BFX9 port map( A => n1667, Z => n1668);
   U141 : HS65_LH_BFX9 port map( A => n1667, Z => n1670);
   U142 : HS65_LH_BFX9 port map( A => n1767, Z => n1647);
   U143 : HS65_LH_AO22X9 port map( A => n163_port, B => n109_port, C => 
                           n161_port, D => n1646, Z => n419);
   U144 : HS65_LH_BFX9 port map( A => n1767, Z => n1649);
   U145 : HS65_LH_BFX9 port map( A => n1767, Z => n1650);
   U146 : HS65_LH_BFX9 port map( A => n1767, Z => n1648);
   U147 : HS65_LH_AO22X9 port map( A => n248, B => n1749, C => n178_port, D => 
                           n1752, Z => n334);
   U148 : HS65_LH_AO22X9 port map( A => n261, B => n1749, C => n133_port, D => 
                           n1755, Z => n304);
   U149 : HS65_LH_AO22X9 port map( A => n250, B => n1749, C => n116_port, D => 
                           n1755, Z => n295);
   U150 : HS65_LH_AO12X9 port map( A => n1651, B => n275, C => n211_port, Z => 
                           n377);
   U151 : HS65_LH_BFX9 port map( A => n1673, Z => n1676);
   U152 : HS65_LH_OAI222X2 port map( A => n221_port, B => n1700, C => n1699, D 
                           => n220_port, E => n396, F => n1701, Z => n160_port)
                           ;
   U153 : HS65_LH_IVX9 port map( A => n221_port, Z => n1767);
   U154 : HS65_LH_OAI222X2 port map( A => n221_port, B => n1729, C => n220_port
                           , D => n1730, E => n396, F => n1728, Z => n121_port)
                           ;
   U155 : HS65_LH_NAND3X5 port map( A => n97, B => n1753, C => n99_port, Z => 
                           n190_port);
   U156 : HS65_LH_NOR2X6 port map( A => n434, B => n193_port, Z => n111_port);
   U157 : HS65_LH_OAI22X6 port map( A => n396, B => n1729, C => n221_port, D =>
                           n1730, Z => n168_port);
   U158 : HS65_LH_OAI22X6 port map( A => n396, B => n1700, C => n221_port, D =>
                           n1699, Z => n182_port);
   U159 : HS65_LH_NAND3X5 port map( A => n433, B => n1753, C => n97, Z => n434)
                           ;
   U160 : HS65_LH_NOR2X6 port map( A => n190_port, B => n193_port, Z => 
                           n212_port);
   U161 : HS65_LH_NOR2AX3 port map( A => alu_i(5), B => n1800, Z => n433);
   U162 : HS65_LH_NOR2X6 port map( A => n434, B => n306, Z => n1643);
   U163 : HS65_LH_NOR2X6 port map( A => n434, B => n306, Z => n113_port);
   U164 : HS65_LH_NOR2X6 port map( A => n434, B => n306, Z => n1644);
   U165 : HS65_LH_OAI222X2 port map( A => n1762, B => n306, C => n1758, D => 
                           n189_port, E => n1764, F => n307, Z => n265);
   U166 : HS65_LH_IVX9 port map( A => n310, Z => n1764);
   U167 : HS65_LH_OAI21X3 port map( A => n221_port, B => n421, C => n96, Z => 
                           n200_port);
   U168 : HS65_LH_NOR2X6 port map( A => n1761, B => n1758, Z => n364);
   U169 : HS65_LH_NOR2X6 port map( A => n192_port, B => n306, Z => n120_port);
   U170 : HS65_LH_OAI32X5 port map( A => n427, B => alu_i(7), C => n428, D => 
                           n429, E => n1791, Z => n426);
   U171 : HS65_LH_AOI12X2 port map( A => n1686, B => n1699, C => n1682, Z => 
                           n429);
   U172 : HS65_LH_AOI22X6 port map( A => N648, B => n99_port, C => N647, D => 
                           n1799, Z => n428);
   U173 : HS65_LH_NOR2X6 port map( A => n305, B => n307, Z => n275);
   U174 : HS65_LH_NOR2X6 port map( A => n190_port, B => n306, Z => n145_port);
   U175 : HS65_LH_NOR2X6 port map( A => alu_i(5), B => alu_i(6), Z => n104_port
                           );
   U176 : HS65_LH_NOR2X6 port map( A => n190_port, B => n306, Z => n1646);
   U177 : HS65_LH_OAI212X5 port map( A => n1763, B => n306, C => n1762, D => 
                           n307, E => n308, Z => n133_port);
   U178 : HS65_LH_IVX9 port map( A => n309, Z => n1763);
   U179 : HS65_LH_NAND3X5 port map( A => n1651, B => alu_i(10), C => n1759, Z 
                           => n308);
   U180 : HS65_LH_NOR2X6 port map( A => n190_port, B => n306, Z => n1645);
   U181 : HS65_LH_NOR2X6 port map( A => n305, B => n306, Z => n273);
   U182 : HS65_LH_AOI222X2 port map( A => n211_port, B => n1711, C => n212_port
                           , D => n259, E => n214_port, F => n260, Z => n258);
   U183 : HS65_LH_AOI222X2 port map( A => n211_port, B => n1712, C => n212_port
                           , D => n248, E => n214_port, F => n249, Z => n247);
   U184 : HS65_LH_AOI222X2 port map( A => n211_port, B => n1713, C => n212_port
                           , D => n229, E => n214_port, F => n230, Z => n228);
   U185 : HS65_LH_AOI222X2 port map( A => n1754, B => n199_port, C => n1644, D 
                           => n148_port, E => n1703, F => n200_port, Z => 
                           n198_port);
   U186 : HS65_LH_NOR2X6 port map( A => n192_port, B => n307, Z => n109_port);
   U187 : HS65_LH_NAND2X7 port map( A => n1771, B => n1769, Z => n396);
   U188 : HS65_LH_NOR2X6 port map( A => n1800, B => alu_i(5), Z => n99_port);
   U189 : HS65_LH_AOI212X4 port map( A => n273, B => n144_port, C => n1646, D 
                           => n215_port, E => n315, Z => n314);
   U190 : HS65_LH_OAI212X5 port map( A => n316, B => n1722, C => n1766, D => 
                           n317, E => n318, Z => n315);
   U191 : HS65_LH_IVX9 port map( A => n213_port, Z => n1766);
   U192 : HS65_LH_CBI4I1X5 port map( A => n1686, B => n1722, C => n1682, D => 
                           alu_i(65), Z => n318);
   U193 : HS65_LH_AOI212X4 port map( A => n211_port, B => n1703, C => n212_port
                           , D => n310, E => n342, Z => n337);
   U194 : HS65_LH_AO22X9 port map( A => n343, B => n214_port, C => n260, D => 
                           n145_port, Z => n342);
   U195 : HS65_LH_AOI212X4 port map( A => n273, B => n161_port, C => n212_port,
                           D => n230, E => n282, Z => n281);
   U196 : HS65_LH_AO22X9 port map( A => n1709, B => n211_port, C => n283, D => 
                           n214_port, Z => n282);
   U197 : HS65_LH_NOR2X6 port map( A => n1730, B => n396, Z => n150_port);
   U198 : HS65_LH_AOI212X4 port map( A => alu_i(65), B => n1672, C => n1686, D 
                           => n1738, E => n1682, Z => n316);
   U199 : HS65_LH_IVX9 port map( A => alu_i(7), Z => n1801);
   U200 : HS65_LH_NAND2X7 port map( A => n1758, B => n1761, Z => n307);
   U201 : HS65_LH_OAI212X5 port map( A => alu_i(62), B => n92, C => n119_port, 
                           D => n1737, E => n1681, Z => n339);
   U202 : HS65_LH_OAI212X5 port map( A => alu_i(53), B => n1684, C => n119_port
                           , D => n1734, E => n95, Z => n410);
   U203 : HS65_LH_MX41X7 port map( D0 => n1706, S0 => n1652, D1 => n1705, S1 =>
                           n1649, D2 => n1704, S2 => n1658, D3 => n1703, S3 => 
                           n1669, Z => n142_port);
   U204 : HS65_LH_MX41X7 port map( D0 => n1705, S0 => n1653, D1 => n1704, S1 =>
                           n1650, D2 => n1703, S2 => n1658, D3 => alu_i(13), S3
                           => n1670, Z => n161_port);
   U205 : HS65_LH_MX41X7 port map( D0 => n1727, S0 => n1653, D1 => alu_i(39), 
                           S1 => n1650, D2 => alu_i(40), S2 => n1659, D3 => 
                           alu_i(41), S3 => n1670, Z => n129_port);
   U206 : HS65_LH_OAI212X5 port map( A => n220_port, B => n1728, C => n221_port
                           , D => n1729, E => n222_port, Z => n218_port);
   U207 : HS65_LH_AOI12X2 port map( A => n1727, B => n1668, C => n150_port, Z 
                           => n222_port);
   U208 : HS65_LH_OAI212X5 port map( A => alu_i(71), B => n1683, C => n1671, D 
                           => n1740, E => n235, Z => n251);
   U209 : HS65_LH_OAI212X5 port map( A => alu_i(11), B => n92, C => n119_port, 
                           D => n1700, E => n1681, Z => n348);
   U210 : HS65_LH_OAI212X5 port map( A => alu_i(12), B => n1683, C => n1671, D 
                           => n1701, E => n1680, Z => n242);
   U211 : HS65_LH_OAI212X5 port map( A => alu_i(13), B => n92, C => n119_port, 
                           D => n1702, E => n1680, Z => n202_port);
   U212 : HS65_LH_OAI212X5 port map( A => alu_i(47), B => n1684, C => n1671, D 
                           => n1732, E => n1680, Z => n179_port);
   U213 : HS65_LH_OAI212X5 port map( A => alu_i(50), B => n1684, C => n1671, D 
                           => n1733, E => n1680, Z => n134_port);
   U214 : HS65_LH_OAI212X5 port map( A => alu_i(56), B => n1684, C => n119_port
                           , D => n1735, E => n1679, Z => n390);
   U215 : HS65_LH_OAI212X5 port map( A => alu_i(59), B => n1684, C => n119_port
                           , D => n1736, E => n1681, Z => n369);
   U216 : HS65_LH_MX41X7 port map( D0 => n1723, S0 => n1653, D1 => n1724, S1 =>
                           n1767, D2 => n1725, S2 => n1659, D3 => n1726, S3 => 
                           n1670, Z => n132_port);
   U217 : HS65_LH_IVX9 port map( A => n192_port, Z => n1754);
   U218 : HS65_LH_IVX9 port map( A => n305, Z => n1755);
   U219 : HS65_LH_NOR3X4 port map( A => n104_port, B => alu_i(8), C => alu_i(7)
                           , Z => n103_port);
   U220 : HS65_LH_MX41X7 port map( D0 => n1725, S0 => n1653, D1 => n1726, S1 =>
                           n1650, D2 => n1727, S2 => n1658, D3 => alu_i(39), S3
                           => n1670, Z => n163_port);
   U221 : HS65_LH_NOR2X6 port map( A => n421, B => n220_port, Z => n203_port);
   U222 : HS65_LH_MX41X7 port map( D0 => n1711, S0 => n1653, D1 => n1712, S1 =>
                           n1650, D2 => n1713, S2 => n1659, D3 => n1714, S3 => 
                           n1670, Z => n130_port);
   U223 : HS65_LH_MX41X7 port map( D0 => n1724, S0 => n1652, D1 => n1725, S1 =>
                           n1649, D2 => n1726, S2 => n1657, D3 => n1727, S3 => 
                           n1669, Z => n110_port);
   U224 : HS65_LH_MX41X7 port map( D0 => alu_i(32), S0 => n1653, D1 => 
                           alu_i(33), S1 => n1650, D2 => n1723, S2 => n1659, D3
                           => n1724, S3 => n1670, Z => n164_port);
   U225 : HS65_LH_MX41X7 port map( D0 => n1719, S0 => n1651, D1 => n1720, S1 =>
                           n1647, D2 => alu_i(32), S2 => n1656, D3 => alu_i(33)
                           , S3 => n1668, Z => n136_port);
   U226 : HS65_LH_MX41X7 port map( D0 => n1715, S0 => n1653, D1 => n1716, S1 =>
                           n1650, D2 => n1717, S2 => n1659, D3 => n1718, S3 => 
                           n1670, Z => n128_port);
   U227 : HS65_LH_MX41X7 port map( D0 => n1716, S0 => n1652, D1 => n1717, S1 =>
                           n1649, D2 => n1718, S2 => n1657, D3 => n1719, S3 => 
                           n1669, Z => n112_port);
   U228 : HS65_LH_MX41X7 port map( D0 => n1704, S0 => n1652, D1 => n1703, S1 =>
                           n1648, D2 => alu_i(13), S2 => n1657, D3 => alu_i(12)
                           , S3 => n1669, Z => n181_port);
   U229 : HS65_LH_MX41X7 port map( D0 => n1712, S0 => n1652, D1 => n1713, S1 =>
                           n1649, D2 => n1714, S2 => n1658, D3 => n1715, S3 => 
                           n1669, Z => n114_port);
   U230 : HS65_LH_MX41X7 port map( D0 => n1717, S0 => n1652, D1 => n1716, S1 =>
                           n1648, D2 => n1715, S2 => n1657, D3 => n1714, S3 => 
                           n1669, Z => n230);
   U231 : HS65_LH_MX41X7 port map( D0 => n1718, S0 => n1651, D1 => n1717, S1 =>
                           n1648, D2 => n1716, S2 => n1656, D3 => n1715, S3 => 
                           n1669, Z => n215_port);
   U232 : HS65_LH_NOR2X6 port map( A => n192_port, B => n193_port, Z => 
                           n151_port);
   U233 : HS65_LH_NOR2X6 port map( A => alu_i(8), B => alu_i(9), Z => n432);
   U234 : HS65_LH_MX41X7 port map( D0 => n1726, S0 => n1652, D1 => n1727, S1 =>
                           n1649, D2 => alu_i(39), S2 => n1658, D3 => alu_i(40)
                           , S3 => n1669, Z => n141_port);
   U235 : HS65_LH_MX41X7 port map( D0 => n1709, S0 => n1653, D1 => n1647, S1 =>
                           n1708, D2 => n1707, S2 => n1658, D3 => n1706, S3 => 
                           n1670, Z => n288);
   U236 : HS65_LH_MX41X7 port map( D0 => n1710, S0 => n1652, D1 => n1709, S1 =>
                           n1649, D2 => n1656, S2 => n1708, D3 => n1707, S3 => 
                           n1669, Z => n276);
   U237 : HS65_LH_MX41X7 port map( D0 => n1718, S0 => n1653, D1 => n1719, S1 =>
                           n1650, D2 => n1720, S2 => n1658, D3 => alu_i(32), S3
                           => n1670, Z => n153_port);
   U238 : HS65_LH_IVX9 port map( A => n306, Z => n1757);
   U239 : HS65_LH_MX41X7 port map( D0 => n1715, S0 => n1652, D1 => n1714, S1 =>
                           n1648, D2 => n1713, S2 => n1657, D3 => n1712, S3 => 
                           n1669, Z => n260);
   U240 : HS65_LH_MX41X7 port map( D0 => alu_i(33), S0 => n1652, D1 => n1723, 
                           S1 => n1650, D2 => n1724, S2 => n1658, D3 => n1725, 
                           S3 => n1670, Z => n155_port);
   U241 : HS65_LH_MX41X7 port map( D0 => n1707, S0 => n1653, D1 => n1647, S1 =>
                           n1708, D2 => n1709, S2 => n1659, D3 => n1710, S3 => 
                           n1670, Z => n131_port);
   U242 : HS65_LH_MX41X7 port map( D0 => n1711, S0 => n1652, D1 => n1710, S1 =>
                           n1649, D2 => n1709, S2 => n1658, D3 => n1668, S3 => 
                           n1708, Z => n310);
   U243 : HS65_LH_MX41X7 port map( D0 => n1716, S0 => n1651, D1 => n1715, S1 =>
                           n1648, D2 => n1714, S2 => n1657, D3 => n1713, S3 => 
                           n1669, Z => n249);
   U244 : HS65_LH_MX41X7 port map( D0 => n1713, S0 => n1652, D1 => n1712, S1 =>
                           n1648, D2 => n1711, S2 => n1657, D3 => n1710, S3 => 
                           n1669, Z => n283);
   U245 : HS65_LH_MX41X7 port map( D0 => n1714, S0 => n1652, D1 => n1713, S1 =>
                           n1648, D2 => n1712, S2 => n1657, D3 => n1711, S3 => 
                           n1669, Z => n277);
   U246 : HS65_LH_MX41X7 port map( D0 => alu_i(33), S0 => n1651, D1 => 
                           alu_i(32), S1 => n1647, D2 => n1720, S2 => n1656, D3
                           => n1719, S3 => n1668, Z => n213_port);
   U247 : HS65_LH_IVX9 port map( A => n193_port, Z => n1759);
   U248 : HS65_LH_MX41X7 port map( D0 => n1719, S0 => n1651, D1 => n1718, S1 =>
                           n1648, D2 => n1717, S2 => n1657, D3 => n1716, S3 => 
                           n1669, Z => n259);
   U249 : HS65_LH_MX41X7 port map( D0 => alu_i(32), S0 => n1651, D1 => n1720, 
                           S1 => n1647, D2 => n1719, S2 => n1657, D3 => n1718, 
                           S3 => n1668, Z => n229);
   U250 : HS65_LH_IVX9 port map( A => n220_port, Z => n1770);
   U251 : HS65_LH_NAND2X7 port map( A => alu_i(8), B => n1796, Z => n427);
   U252 : HS65_LH_MX41X7 port map( D0 => n1720, S0 => n1651, D1 => n1719, S1 =>
                           n1648, D2 => n1718, S2 => n1656, D3 => n1717, S3 => 
                           n1668, Z => n248);
   U253 : HS65_LH_MX41X7 port map( D0 => n1651, S0 => n1708, D1 => n1707, S1 =>
                           n1648, D2 => n1706, S2 => n1657, D3 => n1705, S3 => 
                           n1669, Z => n296);
   U254 : HS65_LH_MX41X7 port map( D0 => n1704, S0 => n1651, D1 => n1705, S1 =>
                           n1648, D2 => n1706, S2 => n1657, D3 => n1707, S3 => 
                           n1668, Z => n177_port);
   U255 : HS65_LH_MX41X7 port map( D0 => n1714, S0 => n1653, D1 => n1715, S1 =>
                           n1650, D2 => n1716, S2 => n1658, D3 => n1717, S3 => 
                           n1670, Z => n154_port);
   U256 : HS65_LH_MX41X7 port map( D0 => n1713, S0 => n1653, D1 => n1714, S1 =>
                           n1650, D2 => n1715, S2 => n1659, D3 => n1716, S3 => 
                           n1670, Z => n170_port);
   U257 : HS65_LH_MX41X7 port map( D0 => n1717, S0 => n1653, D1 => n1718, S1 =>
                           n1650, D2 => n1719, S2 => n1658, D3 => n1720, S3 => 
                           n1670, Z => n172_port);
   U258 : HS65_LH_MX41X7 port map( D0 => n1720, S0 => n1652, D1 => alu_i(32), 
                           S1 => n1648, D2 => alu_i(33), S2 => n1657, D3 => 
                           n1723, S3 => n1669, Z => n123_port);
   U259 : HS65_LH_MX41X7 port map( D0 => n1703, S0 => n1652, D1 => alu_i(13), 
                           S1 => n1649, D2 => n1656, S2 => alu_i(12), D3 => 
                           n1668, S3 => alu_i(11), Z => n309);
   U260 : HS65_LH_MX41X7 port map( D0 => n1651, S0 => n1708, D1 => n1709, S1 =>
                           n1648, D2 => n1710, S2 => n1656, D3 => n1711, S3 => 
                           n1668, Z => n115_port);
   U261 : HS65_LH_MX41X7 port map( D0 => n1712, S0 => n1652, D1 => n1711, S1 =>
                           n1649, D2 => n1710, S2 => n1657, D3 => n1709, S3 => 
                           n1669, Z => n297);
   U262 : HS65_LH_NAND2X7 port map( A => alu_i(5), B => n1800, Z => n102_port);
   U263 : HS65_LH_MX41X7 port map( D0 => n1707, S0 => n1652, D1 => n1706, S1 =>
                           n1649, D2 => n1705, S2 => n1658, D3 => n1704, S3 => 
                           n1669, Z => n343);
   U264 : HS65_LH_MX41X7 port map( D0 => n1709, S0 => n1653, D1 => n1710, S1 =>
                           n1650, D2 => n1711, S2 => n1658, D3 => n1712, S3 => 
                           n1670, Z => n171_port);
   U265 : HS65_LH_IVX9 port map( A => alu_i(6), Z => n1800);
   U266 : HS65_LH_MX41X7 port map( D0 => n1710, S0 => n1652, D1 => n1711, S1 =>
                           n1649, D2 => n1712, S2 => n1658, D3 => n1713, S3 => 
                           n1670, Z => n146_port);
   U267 : HS65_LH_MX41X7 port map( D0 => n1703, S0 => n1653, D1 => n1704, S1 =>
                           n1650, D2 => n1705, S2 => n1659, D3 => n1706, S3 => 
                           n1670, Z => n194_port);
   U268 : HS65_LH_MX41X7 port map( D0 => n1706, S0 => n1652, D1 => n1707, S1 =>
                           n1649, D2 => n1656, S2 => n1708, D3 => n1709, S3 => 
                           n1669, Z => n148_port);
   U269 : HS65_LH_MX41X7 port map( D0 => n1705, S0 => n1651, D1 => n1706, S1 =>
                           n1647, D2 => n1707, S2 => n1656, D3 => n1668, S3 => 
                           n1708, Z => n166_port);
   U270 : HS65_LH_OAI21X3 port map( A => n1720, B => n1685, C => n1680, Z => 
                           n332);
   U271 : HS65_LH_OAI21X3 port map( A => n1723, B => n1685, C => n1680, Z => 
                           n302);
   U272 : HS65_LH_OAI21X3 port map( A => n1724, B => n1685, C => n1680, Z => 
                           n293);
   U273 : HS65_LH_OAI21X3 port map( A => n1726, B => n1685, C => n1680, Z => 
                           n270);
   U274 : HS65_LH_OAI21X3 port map( A => n1709, B => n1683, C => n95, Z => n417
                           );
   U275 : HS65_LH_IVX9 port map( A => alu_i(9), Z => n1796);
   U276 : HS65_LH_MX41X7 port map( D0 => n1726, S0 => n1651, D1 => n1725, S1 =>
                           n1647, D2 => n1724, S2 => n1656, D3 => n1723, S3 => 
                           n1668, Z => n216_port);
   U277 : HS65_LH_MX41X7 port map( D0 => n1724, S0 => n1651, D1 => n1723, S1 =>
                           n1647, D2 => alu_i(33), S2 => n1656, D3 => alu_i(32)
                           , S3 => n1668, Z => n250);
   U278 : HS65_LH_MX41X7 port map( D0 => n1723, S0 => n1651, D1 => alu_i(33), 
                           S1 => n1647, D2 => alu_i(32), S2 => n1656, D3 => 
                           n1720, S3 => n1668, Z => n261);
   U279 : HS65_LH_OAI21X3 port map( A => n1731, B => n1685, C => n206_port, Z 
                           => n243);
   U280 : HS65_LH_OAI21X3 port map( A => n1705, B => n1685, C => n1679, Z => 
                           n169_port);
   U281 : HS65_LH_OAI21X3 port map( A => n1707, B => n1685, C => n95, Z => 
                           n135_port);
   U282 : HS65_LH_OAI21X3 port map( A => n1713, B => n1685, C => n1679, Z => 
                           n391);
   U283 : HS65_LH_OAI21X3 port map( A => n1714, B => n1685, C => n95, Z => n385
                           );
   U284 : HS65_LH_OAI21X3 port map( A => n1715, B => n1685, C => n1679, Z => 
                           n378);
   U285 : HS65_LH_OAI21X3 port map( A => n1716, B => n1685, C => n95, Z => n370
                           );
   U286 : HS65_LH_OAI21X3 port map( A => n1717, B => n1685, C => n1679, Z => 
                           n363);
   U287 : HS65_LH_OAI21X3 port map( A => n1718, B => n1685, C => n95, Z => n356
                           );
   U288 : HS65_LH_OAI21X3 port map( A => n1727, B => n1685, C => n1680, Z => 
                           n264);
   U289 : HS65_LH_MX41X7 port map( D0 => n1725, S0 => n1651, D1 => n1724, S1 =>
                           n1647, D2 => n1723, S2 => n1656, D3 => alu_i(33), S3
                           => n1668, Z => n231);
   U290 : HS65_LH_OAI21X3 port map( A => n1704, B => n1683, C => n1679, Z => 
                           n180_port);
   U291 : HS65_LH_OAI21X3 port map( A => n1706, B => n92, C => n95, Z => 
                           n152_port);
   U292 : HS65_LH_OAI21X3 port map( A => n1708, B => n1683, C => n1679, Z => 
                           n118_port);
   U293 : HS65_LH_NOR3X4 port map( A => n1796, B => alu_i(8), C => n435, Z => 
                           alu_o(32));
   U294 : HS65_LH_AOI33X5 port map( A => n104_port, B => alu_i(7), C => N714, D
                           => n433, E => n1801, F => N713, Z => n435);
   U295 : HS65_LH_OAI21X3 port map( A => n1711, B => n92, C => n95, Z => n404);
   U296 : HS65_LH_OAI21X3 port map( A => n1712, B => n1683, C => n1679, Z => 
                           n398);
   U297 : HS65_LH_AO33X9 port map( A => n1760, B => n1758, C => n1752, D => 
                           n1755, E => n144_port, F => n1759, Z => n272);
   U298 : HS65_LH_AO222X4 port map( A => n1659, B => n1725, C => n1668, D => 
                           n1724, E => n1647, F => n1726, Z => n263);
   U299 : HS65_LH_AO222X4 port map( A => n1659, B => n1726, C => n1668, D => 
                           n1725, E => n1647, F => n1727, Z => n252);
   U300 : HS65_LH_AO222X4 port map( A => n1659, B => n1727, C => n1668, D => 
                           n1726, E => n1647, F => alu_i(39), Z => n233);
   U301 : HS65_LH_AO312X9 port map( A => n1759, B => n160_port, C => n1755, D 
                           => n1725, E => n286, F => n287, Z => n285);
   U302 : HS65_LH_CBI4I6X5 port map( A => n1725, B => n1684, C => n1679, D => 
                           n1739, Z => n287);
   U303 : HS65_LH_OAI212X5 port map( A => alu_i(68), B => n1683, C => n1671, D 
                           => n1739, E => n1681, Z => n286);
   U304 : HS65_LH_BFX9 port map( A => n100_port, Z => n1673);
   U305 : HS65_LH_NOR3X4 port map( A => n1797, B => alu_i(7), C => n102_port, Z
                           => n100_port);
   U306 : HS65_LH_BFX9 port map( A => n201_port, Z => n1667);
   U307 : HS65_LH_NOR2X6 port map( A => n1769, B => n1771, Z => n201_port);
   U308 : HS65_LH_IVX9 port map( A => n357, Z => n1760);
   U309 : HS65_LH_AO22X9 port map( A => n1705, B => n211_port, C => n288, D => 
                           n214_port, Z => n327);
   U310 : HS65_LH_AO22X9 port map( A => n1706, B => n211_port, C => n276, D => 
                           n214_port, Z => n319);
   U311 : HS65_LH_BFX9 port map( A => n1741, Z => n1743);
   U312 : HS65_LH_BFX9 port map( A => n1741, Z => n1744);
   U313 : HS65_LH_BFX9 port map( A => n1741, Z => n1745);
   U314 : HS65_LH_BFX9 port map( A => n1742, Z => n1746);
   U315 : HS65_LH_BFX9 port map( A => n1742, Z => n1747);
   U316 : HS65_LH_BFX9 port map( A => n1742, Z => n1748);
   U317 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_0_port, B => n1693, C => 
                           N162, D => n1689, Z => n462);
   U318 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_1_port, B => n1696, C => 
                           N195, D => n1691, Z => n495);
   U319 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_2_port, B => n1696, C => 
                           N196, D => n1691, Z => n496);
   U320 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_3_port, B => n1696, C => 
                           N197, D => n1691, Z => n497);
   U321 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_5_port, B => n1696, C => 
                           N199, D => n1692, Z => n499);
   U322 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_9_port, B => n1696, C => 
                           N203, D => n1692, Z => n503);
   U323 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_11_port, B => n1697, C => 
                           N205, D => n1692, Z => n505);
   U324 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_13_port, B => n1697, C => 
                           N207, D => n1692, Z => n507);
   U325 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_14_port, B => n1697, C => 
                           N208, D => n1692, Z => n508);
   U326 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_15_port, B => n1697, C => 
                           N209, D => n1692, Z => n509);
   U327 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_16_port, B => n1697, C => 
                           N210, D => n1689, Z => n510);
   U328 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_17_port, B => n1697, C => 
                           N211, D => n1690, Z => n511);
   U329 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_18_port, B => n1697, C => 
                           N212, D => n1691, Z => n512);
   U330 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_19_port, B => n1697, C => 
                           N213, D => n1692, Z => n513);
   U331 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_21_port, B => n1697, C => 
                           N215, D => n1689, Z => n515);
   U332 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_24_port, B => n1697, C => 
                           N218, D => n1690, Z => n518);
   U333 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_25_port, B => n1697, C => 
                           N219, D => n1691, Z => n519);
   U334 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_28_port, B => n1697, C => 
                           N222, D => n1689, Z => n522);
   U335 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_29_port, B => n1697, C => 
                           N223, D => n1690, Z => n523);
   U336 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_30_port, B => n1698, C => 
                           N224, D => n1691, Z => n524);
   U337 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_31_port, B => n1698, C => 
                           N225, D => n1692, Z => n525);
   U338 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_12_port, B => n1695, C => 
                           N174, D => n1690, Z => n474);
   U339 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_16_port, B => n1695, C => 
                           N178, D => n1690, Z => n478);
   U340 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_8_port, B => n1696, C => 
                           N202, D => n1692, Z => n502);
   U341 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_8_port, B => n1695, C => 
                           N170, D => n1689, Z => n470);
   U342 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_13_port, B => n1695, C => 
                           N175, D => n1690, Z => n475);
   U343 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_14_port, B => n1695, C => 
                           N176, D => n1690, Z => n476);
   U344 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_15_port, B => n1695, C => 
                           N177, D => n1690, Z => n477);
   U345 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_6_port, B => n1696, C => 
                           N200, D => n1692, Z => n500);
   U346 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_7_port, B => n1696, C => 
                           N201, D => n1692, Z => n501);
   U347 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_26_port, B => n1697, C => 
                           N220, D => n1692, Z => n520);
   U348 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_20_port, B => n1695, C => 
                           N182, D => n1690, Z => n482);
   U349 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_24_port, B => n1696, C => 
                           N186, D => n1691, Z => n486);
   U350 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_31_port, B => n1696, C => 
                           N193, D => n1691, Z => n493);
   U351 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_4_port, B => n1695, C => 
                           N166, D => n1689, Z => n466);
   U352 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_5_port, B => n1695, C => 
                           N167, D => n1689, Z => n467);
   U353 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_9_port, B => n1695, C => 
                           N171, D => n1689, Z => n471);
   U354 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_11_port, B => n1695, C => 
                           N173, D => n1689, Z => n473);
   U355 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_17_port, B => n1695, C => 
                           N179, D => n1690, Z => n479);
   U356 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_18_port, B => n1695, C => 
                           N180, D => n1690, Z => n480);
   U357 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_19_port, B => n1695, C => 
                           N181, D => n1690, Z => n481);
   U358 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_21_port, B => n1695, C => 
                           N183, D => n1690, Z => n483);
   U359 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_25_port, B => n1696, C => 
                           N187, D => n1691, Z => n487);
   U360 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_29_port, B => n1696, C => 
                           N191, D => n1691, Z => n491);
   U361 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_30_port, B => n1696, C => 
                           N192, D => n1691, Z => n492);
   U362 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_1_port, B => n1694, C => 
                           N163, D => n1689, Z => n463);
   U363 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_2_port, B => n1695, C => 
                           N164, D => n1689, Z => n464);
   U364 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_3_port, B => n1695, C => 
                           N165, D => n1689, Z => n465);
   U365 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_6_port, B => n1695, C => 
                           N168, D => n1689, Z => n468);
   U366 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_7_port, B => n1695, C => 
                           N169, D => n1689, Z => n469);
   U367 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_10_port, B => n1695, C => 
                           N172, D => n1689, Z => n472);
   U368 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_22_port, B => n1696, C => 
                           N184, D => n1690, Z => n484);
   U369 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_23_port, B => n1696, C => 
                           N185, D => n1690, Z => n485);
   U370 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_26_port, B => n1696, C => 
                           N188, D => n1691, Z => n488);
   U371 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_27_port, B => n1696, C => 
                           N189, D => n1691, Z => n489);
   U372 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_0_port, B => n1696, C => 
                           N194, D => n1691, Z => n494);
   U373 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_4_port, B => n1696, C => 
                           N198, D => n1692, Z => n498);
   U374 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_10_port, B => n1697, C => 
                           N204, D => n1692, Z => n504);
   U375 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_20_port, B => n1697, C => 
                           N214, D => n1689, Z => n514);
   U376 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_22_port, B => n1697, C => 
                           N216, D => n1690, Z => n516);
   U377 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_23_port, B => n1697, C => 
                           N217, D => n1691, Z => n517);
   U378 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_27_port, B => n1697, C => 
                           N221, D => n1692, Z => n521);
   U379 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_28_port, B => n1696, C => 
                           N190, D => n1691, Z => n490);
   U380 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_12_port, B => n1697, C => 
                           N206, D => n1692, Z => n506);
   U381 : HS65_LH_NAND2X7 port map( A => alu_i(2), B => n1758, Z => n306);
   U382 : HS65_LH_NAND3X5 port map( A => n97, B => n433, C => alu_i(4), Z => 
                           n192_port);
   U383 : HS65_LH_OAI32X5 port map( A => n189_port, B => alu_i(3), C => 
                           n190_port, D => n191_port, E => n1790, Z => 
                           n188_port);
   U384 : HS65_LH_OA12X9 port map( A => n92, B => n1703, C => n95, Z => 
                           n191_port);
   U385 : HS65_LH_OAI32X5 port map( A => n357, B => alu_i(3), C => n192_port, D
                           => n412, E => n1734, Z => n411);
   U386 : HS65_LH_OA12X9 port map( A => n1683, B => n1710, C => n1679, Z => 
                           n412);
   U387 : HS65_LH_OAI32X5 port map( A => n305, B => alu_i(3), C => n189_port, D
                           => n341, E => n1737, Z => n340);
   U388 : HS65_LH_OA12X9 port map( A => n92, B => n1719, C => n95, Z => n341);
   U389 : HS65_LH_NAND3X5 port map( A => n99_port, B => n97, C => alu_i(4), Z 
                           => n305);
   U390 : HS65_LH_AOI222X2 port map( A => n122_port, B => n132_port, C => n1665
                           , D => HI_LO_c_LO_12_port, E => n113_port, F => 
                           n128_port, Z => n402);
   U391 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_31_port, C => 
                           N129, D => n1677, E => N161, F => n1675, Z => 
                           n209_port);
   U392 : HS65_LH_AOI222X2 port map( A => n1643, B => n130_port, C => n1663, D 
                           => HI_LO_c_HI_8_port, E => n1751, F => n131_port, Z 
                           => n126_port);
   U393 : HS65_LH_AOI222X2 port map( A => N114, B => n1677, C => n1665, D => 
                           HI_LO_c_LO_16_port, E => n1752, F => n375, Z => n374
                           );
   U394 : HS65_LH_AOI222X2 port map( A => N113, B => n1677, C => n113_port, D 
                           => n153_port, E => n1665, F => HI_LO_c_LO_15_port, Z
                           => n383);
   U395 : HS65_LH_AOI222X2 port map( A => N111, B => n1677, C => n109_port, D 
                           => n121_port, E => n1665, F => HI_LO_c_LO_13_port, Z
                           => n395);
   U396 : HS65_LH_AOI222X2 port map( A => n1665, B => HI_LO_c_LO_0_port, C => 
                           alu_i(10), D => n430, E => alu_i(11), F => n200_port
                           , Z => n424);
   U397 : HS65_LH_OAI212X5 port map( A => n396, B => n421, C => alu_i(42), D =>
                           n1683, E => n431, Z => n430);
   U398 : HS65_LH_OA12X9 port map( A => n1791, B => n119_port, C => n235, Z => 
                           n431);
   U399 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_1_port, C => 
                           N99, D => n1677, E => N131, F => n1675, Z => n346);
   U400 : HS65_LH_AOI222X2 port map( A => N112, B => n1677, C => n111_port, D 
                           => n164_port, E => n1665, F => HI_LO_c_LO_14_port, Z
                           => n389);
   U401 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_11_port, C => 
                           N141, D => n1675, E => n1660, F => n1711, Z => n408)
                           ;
   U402 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_21_port, C => 
                           N151, D => n1674, E => n1660, F => alu_i(32), Z => 
                           n330);
   U403 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_24_port, C => 
                           N154, D => n1674, E => n1661, F => n1724, Z => n300)
                           ;
   U404 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_25_port, C => 
                           N155, D => n1674, E => n1661, F => n1725, Z => n291)
                           ;
   U405 : HS65_LH_AOI212X4 port map( A => n273, B => n160_port, C => n1645, D 
                           => n230, E => n324, Z => n323);
   U406 : HS65_LH_OAI212X5 port map( A => n325, B => n1721, C => n1765, D => 
                           n317, E => n326, Z => n324);
   U407 : HS65_LH_IVX9 port map( A => n229, Z => n1765);
   U408 : HS65_LH_CBI4I1X5 port map( A => n1686, B => n1721, C => n1682, D => 
                           alu_i(64), Z => n326);
   U409 : HS65_LH_NAND2X7 port map( A => alu_i(3), B => n1761, Z => n193_port);
   U410 : HS65_LH_OAI22X6 port map( A => alu_i(2), B => n141_port, C => 
                           n150_port, D => n1761, Z => n357);
   U411 : HS65_LH_AOI212X4 port map( A => alu_i(64), B => n1672, C => n1686, D 
                           => n1778, E => n1682, Z => n325);
   U412 : HS65_LH_IVX9 port map( A => alu_i(64), Z => n1778);
   U413 : HS65_LH_NAND2X7 port map( A => alu_i(0), B => n1769, Z => n221_port);
   U414 : HS65_LH_OAI21X3 port map( A => alu_i(2), B => n309, C => n405, Z => 
                           n189_port);
   U415 : HS65_LH_OAI21X3 port map( A => n1699, B => n396, C => alu_i(2), Z => 
                           n405);
   U416 : HS65_LH_OAI212X5 port map( A => alu_i(63), B => n92, C => n119_port, 
                           D => n1779, E => n1681, Z => n333);
   U417 : HS65_LH_IVX9 port map( A => alu_i(63), Z => n1779);
   U418 : HS65_LH_OAI212X5 port map( A => alu_i(66), B => n1683, C => n119_port
                           , D => n1777, E => n1681, Z => n303);
   U419 : HS65_LH_IVX9 port map( A => alu_i(66), Z => n1777);
   U420 : HS65_LH_OAI212X5 port map( A => alu_i(67), B => n92, C => n1671, D =>
                           n1776, E => n1681, Z => n294);
   U421 : HS65_LH_IVX9 port map( A => alu_i(67), Z => n1776);
   U422 : HS65_LH_OAI212X5 port map( A => alu_i(69), B => n1683, C => n1671, D 
                           => n1775, E => n1681, Z => n271);
   U423 : HS65_LH_IVX9 port map( A => alu_i(69), Z => n1775);
   U424 : HS65_LH_OAI212X5 port map( A => alu_i(46), B => n1684, C => n1671, D 
                           => n1790, E => n1681, Z => n187_port);
   U425 : HS65_LH_OAI212X5 port map( A => alu_i(52), B => n1684, C => n119_port
                           , D => n1786, E => n1680, Z => n418);
   U426 : HS65_LH_IVX9 port map( A => alu_i(52), Z => n1786);
   U427 : HS65_LH_OAI212X5 port map( A => alu_i(70), B => n92, C => n1671, D =>
                           n1774, E => n235, Z => n262);
   U428 : HS65_LH_IVX9 port map( A => alu_i(70), Z => n1774);
   U429 : HS65_LH_OAI212X5 port map( A => alu_i(72), B => n92, C => n1671, D =>
                           n1773, E => n235, Z => n232);
   U430 : HS65_LH_IVX9 port map( A => alu_i(72), Z => n1773);
   U431 : HS65_LH_OAI212X5 port map( A => alu_i(73), B => n1683, C => n1671, D 
                           => n1772, E => n223_port, Z => n217_port);
   U432 : HS65_LH_IVX9 port map( A => alu_i(73), Z => n1772);
   U433 : HS65_LH_NOR2X6 port map( A => n1682, B => n1661, Z => n223_port);
   U434 : HS65_LH_OAI212X5 port map( A => alu_i(48), B => n1684, C => n1671, D 
                           => n1789, E => n1680, Z => n167_port);
   U435 : HS65_LH_IVX9 port map( A => alu_i(48), Z => n1789);
   U436 : HS65_LH_OAI212X5 port map( A => alu_i(49), B => n1684, C => n1671, D 
                           => n1788, E => n1680, Z => n149_port);
   U437 : HS65_LH_IVX9 port map( A => alu_i(49), Z => n1788);
   U438 : HS65_LH_OAI212X5 port map( A => alu_i(58), B => n1684, C => n119_port
                           , D => n1782, E => n1681, Z => n376);
   U439 : HS65_LH_IVX9 port map( A => alu_i(58), Z => n1782);
   U440 : HS65_LH_OAI212X5 port map( A => alu_i(51), B => n1684, C => n1787, D 
                           => n119_port, E => n1681, Z => n117_port);
   U441 : HS65_LH_IVX9 port map( A => alu_i(51), Z => n1787);
   U442 : HS65_LH_OAI212X5 port map( A => alu_i(54), B => n1684, C => n119_port
                           , D => n1785, E => n95, Z => n403);
   U443 : HS65_LH_IVX9 port map( A => alu_i(54), Z => n1785);
   U444 : HS65_LH_OAI212X5 port map( A => alu_i(55), B => n1684, C => n1671, D 
                           => n1784, E => n1681, Z => n397);
   U445 : HS65_LH_IVX9 port map( A => alu_i(55), Z => n1784);
   U446 : HS65_LH_OAI212X5 port map( A => alu_i(57), B => n1684, C => n119_port
                           , D => n1783, E => n1681, Z => n384);
   U447 : HS65_LH_IVX9 port map( A => alu_i(57), Z => n1783);
   U448 : HS65_LH_OAI212X5 port map( A => alu_i(60), B => n1684, C => n1671, D 
                           => n1781, E => n1681, Z => n362);
   U449 : HS65_LH_IVX9 port map( A => alu_i(60), Z => n1781);
   U450 : HS65_LH_OAI212X5 port map( A => alu_i(61), B => n1684, C => n119_port
                           , D => n1780, E => n1681, Z => n355);
   U451 : HS65_LH_IVX9 port map( A => alu_i(61), Z => n1780);
   U452 : HS65_LH_NAND2X7 port map( A => alu_i(1), B => n1771, Z => n220_port);
   U453 : HS65_LH_IVX9 port map( A => alu_i(3), Z => n1758);
   U454 : HS65_LH_IVX9 port map( A => alu_i(10), Z => n1699);
   U455 : HS65_LH_IVX9 port map( A => alu_i(41), Z => n1730);
   U456 : HS65_LH_IVX9 port map( A => alu_i(11), Z => n1700);
   U457 : HS65_LH_IVX9 port map( A => alu_i(40), Z => n1729);
   U458 : HS65_LH_IVX9 port map( A => alu_i(32), Z => n1721);
   U459 : HS65_LH_IVX9 port map( A => alu_i(33), Z => n1722);
   U460 : HS65_LH_IVX9 port map( A => alu_i(39), Z => n1728);
   U461 : HS65_LH_IVX9 port map( A => alu_i(12), Z => n1701);
   U462 : HS65_LH_IVX9 port map( A => alu_i(13), Z => n1702);
   U463 : HS65_LH_AO222X4 port map( A => n155_port, B => n1757, C => alu_i(3), 
                           D => n1760, E => n153_port, F => n1756, Z => 
                           n199_port);
   U464 : HS65_LH_IVX9 port map( A => alu_i(2), Z => n1761);
   U465 : HS65_LH_OAI21X3 port map( A => alu_i(43), B => n1685, C => n206_port,
                           Z => n349);
   U466 : HS65_LH_OAI21X3 port map( A => alu_i(45), B => n92, C => n206_port, Z
                           => n205_port);
   U467 : HS65_LH_NAND4ABX3 port map( A => n399, B => n400, C => n401, D => 
                           n402, Z => alu_o(12));
   U468 : HS65_LH_MX41X7 port map( D0 => n109_port, S0 => n129_port, D1 => 
                           n1750, S1 => n265, D2 => n1711, S2 => n403, D3 => 
                           alu_i(54), S3 => n404, Z => n400);
   U469 : HS65_LH_AO222X4 port map( A => HI_LO_c_HI_12_port, B => n1664, C => 
                           n1712, D => n1661, E => n130_port, F => n1751, Z => 
                           n399);
   U470 : HS65_LH_AOI222X2 port map( A => N142, B => n1674, C => n111_port, D 
                           => n136_port, E => N110, F => n1677, Z => n401);
   U471 : HS65_LH_NAND4ABX3 port map( A => n105_port, B => n106_port, C => 
                           n107_port, D => n108_port, Z => alu_o(9));
   U472 : HS65_LH_MX41X7 port map( D0 => n1751, S0 => n115_port, D1 => n1750, 
                           S1 => n116_port, D2 => n1708, S2 => n117_port, D3 =>
                           alu_i(51), S3 => n118_port, Z => n106_port);
   U473 : HS65_LH_MX41X7 port map( D0 => N107, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_9_port, D2 => n120_port, S2 => n121_port,
                           D3 => n122_port, S3 => n123_port, Z => n105_port);
   U474 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_9_port, C => 
                           N139, D => n1674, E => n1660, F => n1709, Z => 
                           n107_port);
   U475 : HS65_LH_NAND4ABX3 port map( A => n365, B => n366, C => n367, D => 
                           n368, Z => alu_o(17));
   U476 : HS65_LH_MX41X7 port map( D0 => n1749, S0 => n249, D1 => n1752, S1 => 
                           n350, D2 => n1716, S2 => n369, D3 => alu_i(59), S3 
                           => n370, Z => n366);
   U477 : HS65_LH_MX41X7 port map( D0 => N115, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_17_port, D2 => n1645, S2 => n297, D3 => 
                           n212_port, S3 => n296, Z => n365);
   U478 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_17_port, C => 
                           N147, D => n1674, E => n1660, F => n1717, Z => n367)
                           ;
   U479 : HS65_LH_NAND4ABX3 port map( A => n358, B => n359, C => n360, D => 
                           n361, Z => alu_o(18));
   U480 : HS65_LH_MX41X7 port map( D0 => n1749, S0 => n230, D1 => n1752, S1 => 
                           n241, D2 => n1717, S2 => n362, D3 => alu_i(60), S3 
                           => n363, Z => n359);
   U481 : HS65_LH_MX41X7 port map( D0 => N116, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_18_port, D2 => n212_port, S2 => n288, D3 
                           => n1646, S3 => n283, Z => n358);
   U482 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_18_port, C => 
                           N148, D => n1674, E => n1660, F => n1718, Z => n360)
                           ;
   U483 : HS65_LH_NAND4ABX3 port map( A => n351, B => n352, C => n353, D => 
                           n354, Z => alu_o(19));
   U484 : HS65_LH_MX41X7 port map( D0 => n1749, S0 => n215_port, D1 => n1752, 
                           S1 => n199_port, D2 => n1718, S2 => n355, D3 => 
                           alu_i(61), S3 => n356, Z => n352);
   U485 : HS65_LH_MX41X7 port map( D0 => N117, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_19_port, D2 => n212_port, S2 => n276, D3 
                           => n145_port, S3 => n277, Z => n351);
   U486 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_19_port, C => 
                           N149, D => n1674, E => n1660, F => n1719, Z => n353)
                           ;
   U487 : HS65_LH_NAND4ABX3 port map( A => n371, B => n372, C => n373, D => 
                           n374, Z => alu_o(16));
   U488 : HS65_LH_MX41X7 port map( D0 => n1749, S0 => n260, D1 => n1715, S1 => 
                           n376, D2 => alu_i(10), S2 => n377, D3 => alu_i(58), 
                           S3 => n378, Z => n371);
   U489 : HS65_LH_AO222X4 port map( A => n343, B => n212_port, C => n309, D => 
                           n214_port, E => n310, F => n1646, Z => n372);
   U490 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_16_port, C => 
                           N146, D => n1675, E => n1660, F => n1716, Z => n373)
                           ;
   U491 : HS65_LH_NAND4ABX3 port map( A => n255, B => n256, C => n257, D => 
                           n258, Z => alu_o(28));
   U492 : HS65_LH_MX41X7 port map( D0 => n1645, S0 => n261, D1 => n1727, S1 => 
                           n262, D2 => n1749, S2 => n263, D3 => alu_i(70), S3 
                           => n264, Z => n256);
   U493 : HS65_LH_MX41X7 port map( D0 => N126, S0 => n1678, D1 => n1751, S1 => 
                           n129_port, D2 => n1665, S2 => HI_LO_c_LO_28_port, D3
                           => n1755, S3 => n265, Z => n255);
   U494 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_28_port, C => 
                           N158, D => n1674, E => n1661, F => alu_i(39), Z => 
                           n257);
   U495 : HS65_LH_NAND4ABX3 port map( A => n244, B => n245, C => n246, D => 
                           n247, Z => alu_o(29));
   U496 : HS65_LH_MX41X7 port map( D0 => n1646, S0 => n250, D1 => alu_i(39), S1
                           => n251, D2 => n1749, S2 => n252, D3 => alu_i(71), 
                           S3 => n253, Z => n245);
   U497 : HS65_LH_MX41X7 port map( D0 => N127, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_29_port, D2 => n1751, S2 => n121_port, D3
                           => n1755, S3 => n254, Z => n244);
   U498 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_29_port, C => 
                           N159, D => n1674, E => n1660, F => alu_i(40), Z => 
                           n246);
   U499 : HS65_LH_NAND4ABX3 port map( A => n225_port, B => n226, C => n227, D 
                           => n228, Z => alu_o(30));
   U500 : HS65_LH_MX41X7 port map( D0 => n145_port, S0 => n231, D1 => alu_i(40)
                           , S1 => n232, D2 => n1749, S2 => n233, D3 => 
                           alu_i(72), S3 => n234, Z => n226);
   U501 : HS65_LH_MX41X7 port map( D0 => N128, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_30_port, D2 => n1751, S2 => n168_port, D3
                           => n1755, S3 => n236, Z => n225_port);
   U502 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_30_port, C => 
                           N160, D => n1674, E => n1660, F => alu_i(41), Z => 
                           n227);
   U503 : HS65_LH_NAND4ABX3 port map( A => n207_port, B => n208_port, C => 
                           n209_port, D => n210_port, Z => alu_o(31));
   U504 : HS65_LH_MX41X7 port map( D0 => n1645, S0 => n216_port, D1 => 
                           alu_i(41), S1 => n217_port, D2 => n1749, S2 => 
                           n218_port, D3 => alu_i(73), S3 => n219_port, Z => 
                           n208_port);
   U505 : HS65_LH_AO222X4 port map( A => n1641, B => n150_port, C => n224_port,
                           D => n1755, E => HI_LO_c_LO_31_port, F => n1666, Z 
                           => n207_port);
   U506 : HS65_LH_AOI222X2 port map( A => n211_port, B => n1714, C => n212_port
                           , D => n213_port, E => n214_port, F => n215_port, Z 
                           => n210_port);
   U507 : HS65_LH_NAND4ABX3 port map( A => n237, B => n238, C => n239, D => 
                           n240, Z => alu_o(2));
   U508 : HS65_LH_MX41X7 port map( D0 => n1731, S0 => n242, D1 => n203_port, S1
                           => n1703, D2 => n204_port, S2 => n1704, D3 => 
                           alu_i(12), S3 => n243, Z => n238);
   U509 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_2_port, D1 => 
                           n122_port, S1 => n170_port, D2 => n111_port, S2 => 
                           n171_port, D3 => n1749, S3 => n160_port, Z => n237);
   U510 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_2_port, C => 
                           N100, D => n1677, E => N132, F => n1675, Z => n239);
   U511 : HS65_LH_NAND4ABX3 port map( A => n380, B => n381, C => n382, D => 
                           n383, Z => alu_o(15));
   U512 : HS65_LH_MX41X7 port map( D0 => n150_port, S0 => n109_port, D1 => 
                           n1750, S1 => n224_port, D2 => n1714, S2 => n384, D3 
                           => alu_i(57), S3 => n385, Z => n380);
   U513 : HS65_LH_AO222X4 port map( A => n155_port, B => n111_port, C => 
                           n141_port, D => n122_port, E => n154_port, F => 
                           n1751, Z => n381);
   U514 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_15_port, C => 
                           N145, D => n1674, E => n1660, F => n1715, Z => n382)
                           ;
   U515 : HS65_LH_NAND4ABX3 port map( A => n195_port, B => n196_port, C => 
                           n197_port, D => n198_port, Z => alu_o(3));
   U516 : HS65_LH_MX41X7 port map( D0 => alu_i(45), S0 => n202_port, D1 => 
                           n203_port, S1 => n1704, D2 => n204_port, S2 => n1705
                           , D3 => alu_i(13), S3 => n205_port, Z => n196_port);
   U517 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_3_port, D1 => 
                           n122_port, S1 => n154_port, D2 => n1749, S2 => 
                           n144_port, D3 => n111_port, S3 => n146_port, Z => 
                           n195_port);
   U518 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_3_port, C => 
                           N101, D => n1677, E => N133, F => n1675, Z => 
                           n197_port);
   U519 : HS65_LH_NAND4ABX3 port map( A => n124_port, B => n125_port, C => 
                           n126_port, D => n127_port, Z => alu_o(8));
   U520 : HS65_LH_MX41X7 port map( D0 => n109_port, S0 => n132_port, D1 => 
                           n1750, S1 => n133_port, D2 => n1707, S2 => n134_port
                           , D3 => alu_i(50), S3 => n135_port, Z => n125_port);
   U521 : HS65_LH_MX41X7 port map( D0 => n1661, S0 => n1708, D1 => N138, S1 => 
                           n1675, D2 => N106, S2 => n1678, D3 => n122_port, S3 
                           => n136_port, Z => n124_port);
   U522 : HS65_LH_AOI222X2 port map( A => n111_port, B => n128_port, C => 
                           n120_port, D => n129_port, E => n1665, F => 
                           HI_LO_c_LO_8_port, Z => n127_port);
   U523 : HS65_LH_NAND4ABX3 port map( A => n173_port, B => n174_port, C => 
                           n175_port, D => n176_port, Z => alu_o(5));
   U524 : HS65_LH_MX41X7 port map( D0 => n1643, S0 => n115_port, D1 => n1754, 
                           S1 => n178_port, D2 => n1704, S2 => n179_port, D3 =>
                           alu_i(47), S3 => n180_port, Z => n174_port);
   U525 : HS65_LH_MX41X7 port map( D0 => N103, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_5_port, D2 => n1749, S2 => n181_port, D3 
                           => n145_port, S3 => n182_port, Z => n173_port);
   U526 : HS65_LH_AOI222X2 port map( A => n1662, B => HI_LO_c_HI_5_port, C => 
                           N135, D => n1674, E => n1660, F => n1705, Z => 
                           n175_port);
   U527 : HS65_LH_NAND4ABX3 port map( A => n392, B => n393, C => n394, D => 
                           n395, Z => alu_o(13));
   U528 : HS65_LH_MX41X7 port map( D0 => n1751, S0 => n114_port, D1 => n1643, 
                           S1 => n112_port, D2 => n1712, S2 => n397, D3 => 
                           alu_i(55), S3 => n398, Z => n392);
   U529 : HS65_LH_AO222X4 port map( A => n110_port, B => n122_port, C => n254, 
                           D => n1750, E => n123_port, F => n111_port, Z => 
                           n393);
   U530 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_13_port, C => 
                           N143, D => n1675, E => n1660, F => n1713, Z => n394)
                           ;
   U531 : HS65_LH_NAND4ABX3 port map( A => n344, B => n345, C => n346, D => 
                           n347, Z => alu_o(1));
   U532 : HS65_LH_MX41X7 port map( D0 => alu_i(43), S0 => n348, D1 => n203_port
                           , S1 => alu_i(13), D2 => n204_port, S2 => n1703, D3 
                           => alu_i(11), S3 => n349, Z => n345);
   U533 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_1_port, D1 => 
                           n1749, S1 => n182_port, D2 => n122_port, S2 => 
                           n114_port, D3 => n1754, S3 => n350, Z => n344);
   U534 : HS65_LH_AOI222X2 port map( A => n113_port, B => n177_port, C => 
                           n111_port, D => n115_port, E => alu_i(12), F => 
                           n200_port, Z => n347);
   U535 : HS65_LH_NAND4ABX3 port map( A => n386, B => n387, C => n388, D => 
                           n389, Z => alu_o(14));
   U536 : HS65_LH_MX41X7 port map( D0 => n109_port, S0 => n168_port, D1 => 
                           n1750, S1 => n236, D2 => n1713, S2 => n390, D3 => 
                           alu_i(56), S3 => n391, Z => n386);
   U537 : HS65_LH_AO222X4 port map( A => n172_port, B => n1644, C => n163_port,
                           D => n122_port, E => n170_port, F => n1641, Z => 
                           n387);
   U538 : HS65_LH_AOI222X2 port map( A => n1663, B => HI_LO_c_HI_14_port, C => 
                           N144, D => n1675, E => n1660, F => n1714, Z => n388)
                           ;
   U539 : HS65_LH_NAND4ABX3 port map( A => n406, B => n407, C => n408, D => 
                           n409, Z => alu_o(11));
   U540 : HS65_LH_MX41X7 port map( D0 => n122_port, S0 => n155_port, D1 => 
                           n212_port, S1 => n144_port, D2 => n1751, S2 => 
                           n146_port, D3 => n1749, S3 => n276, Z => n407);
   U541 : HS65_LH_MX41X7 port map( D0 => N109, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_11_port, D2 => n111_port, S2 => n153_port
                           , D3 => n1644, S3 => n154_port, Z => n406);
   U542 : HS65_LH_AOI212X4 port map( A => n1710, B => n410, C => n145_port, D 
                           => n142_port, E => n411, Z => n409);
   U543 : HS65_LH_NAND4ABX3 port map( A => n311, B => n312, C => n313, D => 
                           n314, Z => alu_o(23));
   U544 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_23_port, D1 =>
                           n1661, S1 => n1723, D2 => N153, S2 => n1675, D3 => 
                           N121, S3 => n1678, Z => n312);
   U545 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_23_port, D1 =>
                           n1751, S1 => n155_port, D2 => n1644, S2 => n141_port
                           , D3 => n150_port, S3 => n111_port, Z => n311);
   U546 : HS65_LH_AOI212X4 port map( A => n275, B => n142_port, C => n212_port,
                           D => n277, E => n319, Z => n313);
   U547 : HS65_LH_NAND4ABX3 port map( A => n320, B => n321, C => n322, D => 
                           n323, Z => alu_o(22));
   U548 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_22_port, D1 =>
                           n1661, S1 => alu_i(33), D2 => N152, S2 => n1675, D3 
                           => N120, S3 => n1678, Z => n321);
   U549 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_22_port, D1 =>
                           n1751, S1 => n164_port, D2 => n111_port, S2 => 
                           n168_port, D3 => n113_port, S3 => n163_port, Z => 
                           n320);
   U550 : HS65_LH_AOI212X4 port map( A => n275, B => n161_port, C => n212_port,
                           D => n283, E => n327, Z => n322);
   U551 : HS65_LH_NAND4ABX3 port map( A => n278, B => n279, C => n280, D => 
                           n281, Z => alu_o(26));
   U552 : HS65_LH_AO212X4 port map( A => n231, B => n1642, C => n229, D => 
                           n1645, E => n285, Z => n279);
   U553 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_26_port, D1 =>
                           n113_port, S1 => n168_port, D2 => n1751, S2 => 
                           n163_port, D3 => n275, S3 => n288, Z => n278);
   U554 : HS65_LH_AOI212X4 port map( A => N124, B => n1677, C => N156, D => 
                           n1675, E => n284, Z => n280);
   U555 : HS65_LH_NAND4ABX3 port map( A => n156_port, B => n157_port, C => 
                           n158_port, D => n159_port, Z => alu_o(6));
   U556 : HS65_LH_MX41X7 port map( D0 => n1751, S0 => n166_port, D1 => n1705, 
                           S1 => n167_port, D2 => n151_port, S2 => n168_port, 
                           D3 => alu_i(48), S3 => n169_port, Z => n157_port);
   U557 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_6_port, D1 => 
                           n111_port, S1 => n170_port, D2 => n1644, S2 => 
                           n171_port, D3 => n122_port, S3 => n172_port, Z => 
                           n156_port);
   U558 : HS65_LH_AOI212X4 port map( A => N104, B => n1677, C => N136, D => 
                           n1675, E => n165_port, Z => n158_port);
   U559 : HS65_LH_NAND4ABX3 port map( A => n137_port, B => n138_port, C => 
                           n139_port, D => n140_port, Z => alu_o(7));
   U560 : HS65_LH_MX41X7 port map( D0 => n1751, S0 => n148_port, D1 => n1706, 
                           S1 => n149_port, D2 => n150_port, S2 => n151_port, 
                           D3 => alu_i(49), S3 => n152_port, Z => n138_port);
   U561 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_7_port, D1 => 
                           n122_port, S1 => n153_port, D2 => n111_port, S2 => 
                           n154_port, D3 => n109_port, S3 => n155_port, Z => 
                           n137_port);
   U562 : HS65_LH_AOI212X4 port map( A => N105, B => n1677, C => N137, D => 
                           n1675, E => n147_port, Z => n139_port);
   U563 : HS65_LH_NAND4ABX3 port map( A => n335, B => n336, C => n337, D => 
                           n338, Z => alu_o(20));
   U564 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_20_port, D1 =>
                           n1661, S1 => n1720, D2 => N150, S2 => n1676, D3 => 
                           N118, S3 => n1678, Z => n336);
   U565 : HS65_LH_MX41X7 port map( D0 => n1751, S0 => n136_port, D1 => n1644, 
                           S1 => n132_port, D2 => n111_port, S2 => n129_port, 
                           D3 => n1666, S3 => HI_LO_c_LO_20_port, Z => n335);
   U566 : HS65_LH_AOI212X4 port map( A => n1719, B => n339, C => n1749, D => 
                           n259, E => n340, Z => n338);
   U567 : HS65_LH_NAND4ABX3 port map( A => n422, B => n423, C => n424, D => 
                           n425, Z => alu_o(0));
   U568 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_0_port, D1 => 
                           N130, S1 => n1675, D2 => N98, S2 => n1678, D3 => 
                           n1754, S3 => n375, Z => n422);
   U569 : HS65_LH_AO222X4 port map( A => n194_port, B => n1644, C => n131_port,
                           D => n111_port, E => n130_port, F => n122_port, Z =>
                           n423);
   U570 : HS65_LH_AOI212X4 port map( A => n204_port, B => alu_i(13), C => 
                           n203_port, D => alu_i(12), E => n426, Z => n425);
   U571 : HS65_LH_NAND4ABX3 port map( A => n266, B => n267, C => n268, D => 
                           n269, Z => alu_o(27));
   U572 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_27_port, D1 =>
                           n1661, S1 => n1727, D2 => N157, S2 => n1675, D3 => 
                           N125, S3 => n1678, Z => n267);
   U573 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_27_port, D1 =>
                           n275, S1 => n276, D2 => n211_port, S2 => n1710, D3 
                           => n214_port, S3 => n277, Z => n266);
   U574 : HS65_LH_AOI212X4 port map( A => alu_i(69), B => n270, C => n1726, D 
                           => n271, E => n272, Z => n269);
   U575 : HS65_LH_NAND4ABX3 port map( A => n289, B => n290, C => n291, D => 
                           n292, Z => alu_o(25));
   U576 : HS65_LH_MX41X7 port map( D0 => N123, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_25_port, D2 => n1643, S2 => n121_port, D3
                           => n1751, S3 => n110_port, Z => n289);
   U577 : HS65_LH_MX41X7 port map( D0 => n211_port, S0 => n1708, D1 => 
                           n214_port, S1 => n297, D2 => n212_port, S2 => n249, 
                           D3 => n1646, S3 => n248, Z => n290);
   U578 : HS65_LH_AOI212X4 port map( A => alu_i(67), B => n293, C => n1724, D 
                           => n294, E => n295, Z => n292);
   U579 : HS65_LH_NAND4ABX3 port map( A => n183_port, B => n184_port, C => 
                           n185_port, D => n186_port, Z => alu_o(4));
   U580 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_4_port, D1 => 
                           n1661, S1 => n1704, D2 => N134, S2 => n1676, D3 => 
                           N102, S3 => n1678, Z => n183_port);
   U581 : HS65_LH_MX41X7 port map( D0 => n122_port, S0 => n128_port, D1 => 
                           n1665, S1 => HI_LO_c_LO_4_port, D2 => n120_port, S2 
                           => n132_port, D3 => n109_port, S3 => n136_port, Z =>
                           n184_port);
   U582 : HS65_LH_AOI212X4 port map( A => n151_port, B => n129_port, C => n1703
                           , D => n187_port, E => n188_port, Z => n186_port);
   U583 : HS65_LH_NAND4ABX3 port map( A => n298, B => n299, C => n300, D => 
                           n301, Z => alu_o(24));
   U584 : HS65_LH_MX41X7 port map( D0 => N122, S0 => n1678, D1 => n1751, S1 => 
                           n132_port, D2 => n113_port, S2 => n129_port, D3 => 
                           n1666, S3 => HI_LO_c_LO_24_port, Z => n298);
   U585 : HS65_LH_MX41X7 port map( D0 => n211_port, S0 => n1707, D1 => 
                           n214_port, S1 => n310, D2 => n212_port, S2 => n260, 
                           D3 => n1645, S3 => n259, Z => n299);
   U586 : HS65_LH_AOI212X4 port map( A => alu_i(66), B => n302, C => n1723, D 
                           => n303, E => n304, Z => n301);
   U587 : HS65_LH_NAND4ABX3 port map( A => n328, B => n329, C => n330, D => 
                           n331, Z => alu_o(21));
   U588 : HS65_LH_MX41X7 port map( D0 => n211_port, S0 => n1704, D1 => 
                           n214_port, S1 => n296, D2 => n1646, S2 => n249, D3 
                           => n273, S3 => n182_port, Z => n329);
   U589 : HS65_LH_MX41X7 port map( D0 => N119, S0 => n1678, D1 => n1665, S1 => 
                           HI_LO_c_LO_21_port, D2 => n212_port, S2 => n297, D3 
                           => n275, S3 => n181_port, Z => n328);
   U590 : HS65_LH_AOI212X4 port map( A => alu_i(63), B => n332, C => n1720, D 
                           => n333, E => n334, Z => n331);
   U591 : HS65_LH_NAND4ABX3 port map( A => n413, B => n414, C => n415, D => 
                           n416, Z => alu_o(10));
   U592 : HS65_LH_MX41X7 port map( D0 => n1663, S0 => HI_LO_c_HI_10_port, D1 =>
                           n1661, S1 => n1710, D2 => N140, S2 => n1676, D3 => 
                           N108, S3 => n1677, Z => n414);
   U593 : HS65_LH_MX41X7 port map( D0 => n1666, S0 => HI_LO_c_LO_10_port, D1 =>
                           n122_port, S1 => n164_port, D2 => n1643, S2 => 
                           n170_port, D3 => n1642, S3 => n288, Z => n413);
   U594 : HS65_LH_AOI212X4 port map( A => alu_i(52), B => n417, C => n1709, D 
                           => n418, E => n419, Z => n416);
   U595 : HS65_LH_IVX9 port map( A => alu_i(1), Z => n1769);
   U596 : HS65_LH_IVX9 port map( A => alu_i(0), Z => n1771);
   U597 : HS65_LH_IVX9 port map( A => alu_i(68), Z => n1739);
   U598 : HS65_LH_IVX9 port map( A => alu_i(53), Z => n1734);
   U599 : HS65_LH_IVX9 port map( A => alu_i(62), Z => n1737);
   U600 : HS65_LH_IVX9 port map( A => alu_i(47), Z => n1732);
   U601 : HS65_LH_IVX9 port map( A => alu_i(50), Z => n1733);
   U602 : HS65_LH_IVX9 port map( A => alu_i(56), Z => n1735);
   U603 : HS65_LH_IVX9 port map( A => alu_i(59), Z => n1736);
   U604 : HS65_LH_IVX9 port map( A => alu_i(71), Z => n1740);
   U605 : HS65_LH_IVX9 port map( A => alu_i(65), Z => n1738);
   U606 : HS65_LH_BFX9 port map( A => rst_n, Z => n1741);
   U607 : HS65_LH_BFX9 port map( A => rst_n, Z => n1742);
   U608 : HS65_LH_BFX9 port map( A => alu_i(44), Z => n1731);
   U609 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_26_port, B => n1664, C => 
                           n1726, D => n1661, Z => n284);
   U610 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_6_port, B => n1664, C => 
                           n1706, D => n1661, Z => n165_port);
   U611 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_7_port, B => n1664, C => 
                           n1707, D => n1661, Z => n147_port);
   U612 : HS65_LH_IVX9 port map( A => alu_i(4), Z => n1753);
   U613 : HS65_LH_IVX9 port map( A => alu_i(46), Z => n1790);
   U614 : HS65_LH_IVX9 port map( A => alu_i(42), Z => n1791);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity exe_top is

   port( clk, rst_n : in std_logic;  exe_top_i : in std_logic_vector (134 
         downto 0);  exe_top_o : out std_logic_vector (81 downto 0));

end exe_top;

architecture SYN_Behavioral of exe_top is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component exe_top_DW01_add_0
      port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (11 downto 0);  CO : out std_logic);
   end component;
   
   component alu_ctrl
      port( alu_ctrl_i : in std_logic_vector (9 downto 0);  alu_ctrl_o : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component alu
      port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 
            0);  alu_o : out std_logic_vector (32 downto 0));
   end component;
   
   signal exe_top_o_BRANCH_port, exe_top_o_BRANCH_PC_11_port, 
      exe_top_o_BRANCH_PC_10_port, exe_top_o_BRANCH_PC_9_port, 
      exe_top_o_BRANCH_PC_8_port, exe_top_o_BRANCH_PC_7_port, 
      exe_top_o_BRANCH_PC_6_port, exe_top_o_BRANCH_PC_5_port, 
      exe_top_o_BRANCH_PC_4_port, exe_top_o_BRANCH_PC_3_port, 
      exe_top_o_BRANCH_PC_2_port, exe_top_o_BRANCH_PC_1_port, 
      exe_top_o_BRANCH_PC_0_port, exe_top_o_RESULT_31_port, 
      exe_top_o_RESULT_30_port, exe_top_o_RESULT_29_port, 
      exe_top_o_RESULT_28_port, exe_top_o_RESULT_27_port, 
      exe_top_o_RESULT_26_port, exe_top_o_RESULT_25_port, 
      exe_top_o_RESULT_24_port, exe_top_o_RESULT_23_port, 
      exe_top_o_RESULT_22_port, exe_top_o_RESULT_21_port, 
      exe_top_o_RESULT_20_port, exe_top_o_RESULT_19_port, 
      exe_top_o_RESULT_18_port, exe_top_o_RESULT_17_port, 
      exe_top_o_RESULT_16_port, exe_top_o_RESULT_15_port, 
      exe_top_o_RESULT_14_port, exe_top_o_RESULT_13_port, 
      exe_top_o_RESULT_12_port, exe_top_o_RESULT_11_port, 
      exe_top_o_RESULT_10_port, exe_top_o_RESULT_9_port, 
      exe_top_o_RESULT_8_port, exe_top_o_RESULT_7_port, exe_top_o_RESULT_6_port
      , exe_top_o_RESULT_5_port, exe_top_o_RESULT_4_port, 
      exe_top_o_RESULT_3_port, exe_top_o_RESULT_2_port, exe_top_o_RESULT_1_port
      , exe_top_o_RESULT_0_port, exe_top_o_WRITE_REG_4_port, 
      exe_top_o_WRITE_REG_3_port, exe_top_o_WRITE_REG_2_port, 
      exe_top_o_WRITE_REG_1_port, exe_top_o_WRITE_REG_0_port, src_b_31_port, 
      src_b_30_port, src_b_29_port, src_b_28_port, src_b_27_port, src_b_26_port
      , src_b_25_port, src_b_24_port, src_b_23_port, src_b_22_port, 
      src_b_21_port, src_b_20_port, src_b_19_port, src_b_18_port, src_b_17_port
      , src_b_16_port, src_b_15_port, src_b_14_port, src_b_13_port, 
      src_b_12_port, src_b_11_port, src_b_10_port, src_b_9_port, src_b_8_port, 
      src_b_7_port, src_b_6_port, src_b_5_port, src_b_4_port, src_b_3_port, 
      src_b_2_port, src_b_1_port, src_b_0_port, op_aluCtrl_alu_4_port, 
      op_aluCtrl_alu_3_port, op_aluCtrl_alu_2_port, op_aluCtrl_alu_1_port, 
      op_aluCtrl_alu_0_port, n3, n6, n7, n8, n_1020 : std_logic;

begin
   exe_top_o <= ( exe_top_o_BRANCH_port, exe_top_o_BRANCH_PC_11_port, 
      exe_top_o_BRANCH_PC_10_port, exe_top_o_BRANCH_PC_9_port, 
      exe_top_o_BRANCH_PC_8_port, exe_top_o_BRANCH_PC_7_port, 
      exe_top_o_BRANCH_PC_6_port, exe_top_o_BRANCH_PC_5_port, 
      exe_top_o_BRANCH_PC_4_port, exe_top_o_BRANCH_PC_3_port, 
      exe_top_o_BRANCH_PC_2_port, exe_top_o_BRANCH_PC_1_port, 
      exe_top_o_BRANCH_PC_0_port, exe_top_o_RESULT_31_port, 
      exe_top_o_RESULT_30_port, exe_top_o_RESULT_29_port, 
      exe_top_o_RESULT_28_port, exe_top_o_RESULT_27_port, 
      exe_top_o_RESULT_26_port, exe_top_o_RESULT_25_port, 
      exe_top_o_RESULT_24_port, exe_top_o_RESULT_23_port, 
      exe_top_o_RESULT_22_port, exe_top_o_RESULT_21_port, 
      exe_top_o_RESULT_20_port, exe_top_o_RESULT_19_port, 
      exe_top_o_RESULT_18_port, exe_top_o_RESULT_17_port, 
      exe_top_o_RESULT_16_port, exe_top_o_RESULT_15_port, 
      exe_top_o_RESULT_14_port, exe_top_o_RESULT_13_port, 
      exe_top_o_RESULT_12_port, exe_top_o_RESULT_11_port, 
      exe_top_o_RESULT_10_port, exe_top_o_RESULT_9_port, 
      exe_top_o_RESULT_8_port, exe_top_o_RESULT_7_port, exe_top_o_RESULT_6_port
      , exe_top_o_RESULT_5_port, exe_top_o_RESULT_4_port, 
      exe_top_o_RESULT_3_port, exe_top_o_RESULT_2_port, exe_top_o_RESULT_1_port
      , exe_top_o_RESULT_0_port, exe_top_o_WRITE_REG_4_port, 
      exe_top_o_WRITE_REG_3_port, exe_top_o_WRITE_REG_2_port, 
      exe_top_o_WRITE_REG_1_port, exe_top_o_WRITE_REG_0_port, exe_top_i(97), 
      exe_top_i(96), exe_top_i(95), exe_top_i(94), exe_top_i(93), exe_top_i(92)
      , exe_top_i(91), exe_top_i(90), exe_top_i(89), exe_top_i(88), 
      exe_top_i(87), exe_top_i(86), exe_top_i(85), exe_top_i(84), exe_top_i(83)
      , exe_top_i(82), exe_top_i(81), exe_top_i(80), exe_top_i(79), 
      exe_top_i(78), exe_top_i(77), exe_top_i(76), exe_top_i(75), exe_top_i(74)
      , exe_top_i(73), exe_top_i(72), exe_top_i(71), exe_top_i(70), 
      exe_top_i(69), exe_top_i(68), exe_top_i(67), exe_top_i(66) );
   
   n3 <= '0';
   alu_inst : alu port map( clk => clk, rst_n => rst_n, alu_i(73) => 
                           exe_top_i(129), alu_i(72) => exe_top_i(128), 
                           alu_i(71) => exe_top_i(127), alu_i(70) => 
                           exe_top_i(126), alu_i(69) => exe_top_i(125), 
                           alu_i(68) => exe_top_i(124), alu_i(67) => 
                           exe_top_i(123), alu_i(66) => exe_top_i(122), 
                           alu_i(65) => exe_top_i(121), alu_i(64) => 
                           exe_top_i(120), alu_i(63) => exe_top_i(119), 
                           alu_i(62) => exe_top_i(118), alu_i(61) => 
                           exe_top_i(117), alu_i(60) => exe_top_i(116), 
                           alu_i(59) => exe_top_i(115), alu_i(58) => 
                           exe_top_i(114), alu_i(57) => exe_top_i(113), 
                           alu_i(56) => exe_top_i(112), alu_i(55) => 
                           exe_top_i(111), alu_i(54) => exe_top_i(110), 
                           alu_i(53) => exe_top_i(109), alu_i(52) => 
                           exe_top_i(108), alu_i(51) => exe_top_i(107), 
                           alu_i(50) => exe_top_i(106), alu_i(49) => 
                           exe_top_i(105), alu_i(48) => exe_top_i(104), 
                           alu_i(47) => exe_top_i(103), alu_i(46) => 
                           exe_top_i(102), alu_i(45) => exe_top_i(101), 
                           alu_i(44) => exe_top_i(100), alu_i(43) => 
                           exe_top_i(99), alu_i(42) => exe_top_i(98), alu_i(41)
                           => src_b_31_port, alu_i(40) => src_b_30_port, 
                           alu_i(39) => src_b_29_port, alu_i(38) => 
                           src_b_28_port, alu_i(37) => src_b_27_port, alu_i(36)
                           => src_b_26_port, alu_i(35) => src_b_25_port, 
                           alu_i(34) => src_b_24_port, alu_i(33) => 
                           src_b_23_port, alu_i(32) => src_b_22_port, alu_i(31)
                           => src_b_21_port, alu_i(30) => src_b_20_port, 
                           alu_i(29) => src_b_19_port, alu_i(28) => 
                           src_b_18_port, alu_i(27) => src_b_17_port, alu_i(26)
                           => src_b_16_port, alu_i(25) => src_b_15_port, 
                           alu_i(24) => src_b_14_port, alu_i(23) => 
                           src_b_13_port, alu_i(22) => src_b_12_port, alu_i(21)
                           => src_b_11_port, alu_i(20) => src_b_10_port, 
                           alu_i(19) => src_b_9_port, alu_i(18) => src_b_8_port
                           , alu_i(17) => src_b_7_port, alu_i(16) => 
                           src_b_6_port, alu_i(15) => src_b_5_port, alu_i(14) 
                           => src_b_4_port, alu_i(13) => src_b_3_port, 
                           alu_i(12) => src_b_2_port, alu_i(11) => src_b_1_port
                           , alu_i(10) => src_b_0_port, alu_i(9) => 
                           op_aluCtrl_alu_4_port, alu_i(8) => 
                           op_aluCtrl_alu_3_port, alu_i(7) => 
                           op_aluCtrl_alu_2_port, alu_i(6) => 
                           op_aluCtrl_alu_1_port, alu_i(5) => 
                           op_aluCtrl_alu_0_port, alu_i(4) => exe_top_i(134), 
                           alu_i(3) => exe_top_i(133), alu_i(2) => 
                           exe_top_i(132), alu_i(1) => exe_top_i(131), alu_i(0)
                           => exe_top_i(130), alu_o(32) => 
                           exe_top_o_BRANCH_port, alu_o(31) => 
                           exe_top_o_RESULT_31_port, alu_o(30) => 
                           exe_top_o_RESULT_30_port, alu_o(29) => 
                           exe_top_o_RESULT_29_port, alu_o(28) => 
                           exe_top_o_RESULT_28_port, alu_o(27) => 
                           exe_top_o_RESULT_27_port, alu_o(26) => 
                           exe_top_o_RESULT_26_port, alu_o(25) => 
                           exe_top_o_RESULT_25_port, alu_o(24) => 
                           exe_top_o_RESULT_24_port, alu_o(23) => 
                           exe_top_o_RESULT_23_port, alu_o(22) => 
                           exe_top_o_RESULT_22_port, alu_o(21) => 
                           exe_top_o_RESULT_21_port, alu_o(20) => 
                           exe_top_o_RESULT_20_port, alu_o(19) => 
                           exe_top_o_RESULT_19_port, alu_o(18) => 
                           exe_top_o_RESULT_18_port, alu_o(17) => 
                           exe_top_o_RESULT_17_port, alu_o(16) => 
                           exe_top_o_RESULT_16_port, alu_o(15) => 
                           exe_top_o_RESULT_15_port, alu_o(14) => 
                           exe_top_o_RESULT_14_port, alu_o(13) => 
                           exe_top_o_RESULT_13_port, alu_o(12) => 
                           exe_top_o_RESULT_12_port, alu_o(11) => 
                           exe_top_o_RESULT_11_port, alu_o(10) => 
                           exe_top_o_RESULT_10_port, alu_o(9) => 
                           exe_top_o_RESULT_9_port, alu_o(8) => 
                           exe_top_o_RESULT_8_port, alu_o(7) => 
                           exe_top_o_RESULT_7_port, alu_o(6) => 
                           exe_top_o_RESULT_6_port, alu_o(5) => 
                           exe_top_o_RESULT_5_port, alu_o(4) => 
                           exe_top_o_RESULT_4_port, alu_o(3) => 
                           exe_top_o_RESULT_3_port, alu_o(2) => 
                           exe_top_o_RESULT_2_port, alu_o(1) => 
                           exe_top_o_RESULT_1_port, alu_o(0) => 
                           exe_top_o_RESULT_0_port);
   alu_ctrl_inst : alu_ctrl port map( alu_ctrl_i(9) => exe_top_i(32), 
                           alu_ctrl_i(8) => exe_top_i(31), alu_ctrl_i(7) => 
                           exe_top_i(30), alu_ctrl_i(6) => exe_top_i(29), 
                           alu_ctrl_i(5) => exe_top_i(28), alu_ctrl_i(4) => 
                           exe_top_i(27), alu_ctrl_i(3) => exe_top_i(26), 
                           alu_ctrl_i(2) => exe_top_i(25), alu_ctrl_i(1) => 
                           exe_top_i(24), alu_ctrl_i(0) => exe_top_i(23), 
                           alu_ctrl_o(4) => op_aluCtrl_alu_4_port, 
                           alu_ctrl_o(3) => op_aluCtrl_alu_3_port, 
                           alu_ctrl_o(2) => op_aluCtrl_alu_2_port, 
                           alu_ctrl_o(1) => op_aluCtrl_alu_1_port, 
                           alu_ctrl_o(0) => op_aluCtrl_alu_0_port);
   add_43 : exe_top_DW01_add_0 port map( A(11) => exe_top_i(22), A(10) => 
                           exe_top_i(21), A(9) => exe_top_i(20), A(8) => 
                           exe_top_i(19), A(7) => exe_top_i(18), A(6) => 
                           exe_top_i(17), A(5) => exe_top_i(16), A(4) => 
                           exe_top_i(15), A(3) => exe_top_i(14), A(2) => 
                           exe_top_i(13), A(1) => exe_top_i(12), A(0) => 
                           exe_top_i(11), B(11) => exe_top_i(44), B(10) => 
                           exe_top_i(43), B(9) => exe_top_i(42), B(8) => 
                           exe_top_i(41), B(7) => exe_top_i(40), B(6) => 
                           exe_top_i(39), B(5) => exe_top_i(38), B(4) => 
                           exe_top_i(37), B(3) => exe_top_i(36), B(2) => 
                           exe_top_i(35), B(1) => exe_top_i(34), B(0) => 
                           exe_top_i(33), CI => n3, SUM(11) => 
                           exe_top_o_BRANCH_PC_11_port, SUM(10) => 
                           exe_top_o_BRANCH_PC_10_port, SUM(9) => 
                           exe_top_o_BRANCH_PC_9_port, SUM(8) => 
                           exe_top_o_BRANCH_PC_8_port, SUM(7) => 
                           exe_top_o_BRANCH_PC_7_port, SUM(6) => 
                           exe_top_o_BRANCH_PC_6_port, SUM(5) => 
                           exe_top_o_BRANCH_PC_5_port, SUM(4) => 
                           exe_top_o_BRANCH_PC_4_port, SUM(3) => 
                           exe_top_o_BRANCH_PC_3_port, SUM(2) => 
                           exe_top_o_BRANCH_PC_2_port, SUM(1) => 
                           exe_top_o_BRANCH_PC_1_port, SUM(0) => 
                           exe_top_o_BRANCH_PC_0_port, CO => n_1020);
   U42 : HS65_LH_AO22X9 port map( A => exe_top_i(52), B => exe_top_i(65), C => 
                           exe_top_i(85), D => n6, Z => src_b_19_port);
   U43 : HS65_LH_AO22X9 port map( A => exe_top_i(60), B => exe_top_i(65), C => 
                           exe_top_i(93), D => n7, Z => src_b_27_port);
   U44 : HS65_LH_AO22X9 port map( A => exe_top_i(58), B => exe_top_i(65), C => 
                           exe_top_i(91), D => n7, Z => src_b_25_port);
   U45 : HS65_LH_AO22X9 port map( A => exe_top_i(45), B => exe_top_i(65), C => 
                           exe_top_i(78), D => n6, Z => src_b_12_port);
   U46 : HS65_LH_AO22X9 port map( A => exe_top_i(48), B => exe_top_i(65), C => 
                           exe_top_i(81), D => n6, Z => src_b_15_port);
   U47 : HS65_LH_AO22X9 port map( A => exe_top_i(46), B => exe_top_i(65), C => 
                           exe_top_i(79), D => n6, Z => src_b_13_port);
   U48 : HS65_LH_AO22X9 port map( A => exe_top_i(37), B => exe_top_i(65), C => 
                           exe_top_i(70), D => n6, Z => src_b_4_port);
   U49 : HS65_LH_AO22X9 port map( A => exe_top_i(51), B => exe_top_i(65), C => 
                           exe_top_i(84), D => n6, Z => src_b_18_port);
   U50 : HS65_LH_AO22X9 port map( A => exe_top_i(38), B => exe_top_i(65), C => 
                           exe_top_i(71), D => n7, Z => src_b_5_port);
   U51 : HS65_LH_AO22X9 port map( A => exe_top_i(59), B => exe_top_i(65), C => 
                           exe_top_i(92), D => n7, Z => src_b_26_port);
   U52 : HS65_LH_AO22X9 port map( A => exe_top_i(50), B => exe_top_i(65), C => 
                           exe_top_i(83), D => n6, Z => src_b_17_port);
   U53 : HS65_LH_AO22X9 port map( A => exe_top_i(57), B => exe_top_i(65), C => 
                           exe_top_i(90), D => n7, Z => src_b_24_port);
   U54 : HS65_LH_AO22X9 port map( A => exe_top_i(53), B => exe_top_i(65), C => 
                           exe_top_i(86), D => n7, Z => src_b_20_port);
   U55 : HS65_LH_AO22X9 port map( A => exe_top_i(40), B => exe_top_i(65), C => 
                           exe_top_i(73), D => n6, Z => src_b_7_port);
   U56 : HS65_LH_AO22X9 port map( A => exe_top_i(44), B => exe_top_i(65), C => 
                           exe_top_i(77), D => n6, Z => src_b_11_port);
   U57 : HS65_LH_AO22X9 port map( A => exe_top_i(54), B => exe_top_i(65), C => 
                           exe_top_i(87), D => n7, Z => src_b_21_port);
   U58 : HS65_LH_AO22X9 port map( A => exe_top_i(42), B => exe_top_i(65), C => 
                           exe_top_i(75), D => n7, Z => src_b_9_port);
   U59 : HS65_LH_AO22X9 port map( A => exe_top_i(61), B => exe_top_i(65), C => 
                           exe_top_i(94), D => n7, Z => src_b_28_port);
   U60 : HS65_LH_AO22X9 port map( A => exe_top_i(33), B => exe_top_i(65), C => 
                           exe_top_i(66), D => n6, Z => src_b_0_port);
   U61 : HS65_LH_AO22X9 port map( A => exe_top_i(64), B => exe_top_i(65), C => 
                           exe_top_i(97), D => n6, Z => src_b_31_port);
   U62 : HS65_LH_AO22X9 port map( A => exe_top_i(34), B => exe_top_i(65), C => 
                           exe_top_i(67), D => n6, Z => src_b_1_port);
   U63 : HS65_LH_AO22X9 port map( A => exe_top_i(63), B => exe_top_i(65), C => 
                           exe_top_i(96), D => n7, Z => src_b_30_port);
   U64 : HS65_LH_AO22X9 port map( A => exe_top_i(55), B => exe_top_i(65), C => 
                           exe_top_i(88), D => n7, Z => src_b_22_port);
   U65 : HS65_LH_AO22X9 port map( A => exe_top_i(56), B => exe_top_i(65), C => 
                           exe_top_i(89), D => n7, Z => src_b_23_port);
   U66 : HS65_LH_AO22X9 port map( A => exe_top_i(62), B => exe_top_i(65), C => 
                           exe_top_i(95), D => n7, Z => src_b_29_port);
   U67 : HS65_LH_AO22X9 port map( A => exe_top_i(35), B => exe_top_i(65), C => 
                           exe_top_i(68), D => n7, Z => src_b_2_port);
   U68 : HS65_LH_AO22X9 port map( A => exe_top_i(36), B => exe_top_i(65), C => 
                           exe_top_i(69), D => n7, Z => src_b_3_port);
   U69 : HS65_LH_AO22X9 port map( A => exe_top_i(47), B => exe_top_i(65), C => 
                           exe_top_i(80), D => n6, Z => src_b_14_port);
   U70 : HS65_LH_AO22X9 port map( A => exe_top_i(39), B => exe_top_i(65), C => 
                           exe_top_i(72), D => n6, Z => src_b_6_port);
   U71 : HS65_LH_AO22X9 port map( A => exe_top_i(43), B => exe_top_i(65), C => 
                           exe_top_i(76), D => n6, Z => src_b_10_port);
   U72 : HS65_LH_AO22X9 port map( A => exe_top_i(41), B => exe_top_i(65), C => 
                           exe_top_i(74), D => n7, Z => src_b_8_port);
   U73 : HS65_LH_AO22X9 port map( A => exe_top_i(49), B => exe_top_i(65), C => 
                           exe_top_i(82), D => n6, Z => src_b_16_port);
   U74 : HS65_LH_IVX9 port map( A => exe_top_i(10), Z => n8);
   U75 : HS65_LH_AO22X9 port map( A => exe_top_i(5), B => n8, C => exe_top_i(0)
                           , D => exe_top_i(10), Z => 
                           exe_top_o_WRITE_REG_0_port);
   U76 : HS65_LH_AO22X9 port map( A => exe_top_i(6), B => n8, C => exe_top_i(1)
                           , D => exe_top_i(10), Z => 
                           exe_top_o_WRITE_REG_1_port);
   U77 : HS65_LH_AO22X9 port map( A => exe_top_i(7), B => n8, C => exe_top_i(2)
                           , D => exe_top_i(10), Z => 
                           exe_top_o_WRITE_REG_2_port);
   U78 : HS65_LH_AO22X9 port map( A => exe_top_i(8), B => n8, C => exe_top_i(3)
                           , D => exe_top_i(10), Z => 
                           exe_top_o_WRITE_REG_3_port);
   U79 : HS65_LH_AO22X9 port map( A => exe_top_i(9), B => n8, C => 
                           exe_top_i(10), D => exe_top_i(4), Z => 
                           exe_top_o_WRITE_REG_4_port);
   U80 : HS65_LH_IVX9 port map( A => exe_top_i(65), Z => n6);
   U81 : HS65_LH_IVX9 port map( A => exe_top_i(65), Z => n7);

end SYN_Behavioral;
