
module controller ( .ctrl_i({\ctrl_i[OPCODE][5] , \ctrl_i[OPCODE][4] , 
        \ctrl_i[OPCODE][3] , \ctrl_i[OPCODE][2] , \ctrl_i[OPCODE][1] , 
        \ctrl_i[OPCODE][0] }), .ctrl_o({\ctrl_o[REGDST] , \ctrl_o[ALUSRC_B] , 
        \ctrl_o[MEMTOREG] , \ctrl_o[REGWRITE] , \ctrl_o[MEMWEN_N] , 
        \ctrl_o[BRANCH] , \ctrl_o[CALU_OP][3] , \ctrl_o[CALU_OP][2] , 
        \ctrl_o[CALU_OP][1] , \ctrl_o[CALU_OP][0] }) );
  input \ctrl_i[OPCODE][5] , \ctrl_i[OPCODE][4] , \ctrl_i[OPCODE][3] ,
         \ctrl_i[OPCODE][2] , \ctrl_i[OPCODE][1] , \ctrl_i[OPCODE][0] ;
  output \ctrl_o[REGDST] , \ctrl_o[ALUSRC_B] , \ctrl_o[MEMTOREG] ,
         \ctrl_o[REGWRITE] , \ctrl_o[MEMWEN_N] , \ctrl_o[BRANCH] ,
         \ctrl_o[CALU_OP][3] , \ctrl_o[CALU_OP][2] , \ctrl_o[CALU_OP][1] ,
         \ctrl_o[CALU_OP][0] ;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n3, n4, n5, n6, n7, n8, n24;

  HS65_LH_IVX9 U3 ( .A(1'b1), .Z(\ctrl_o[CALU_OP][3] ) );
  HS65_LH_OAI31X5 U5 ( .A(n22), .B(n14), .C(n15), .D(n8), .Z(n21) );
  HS65_LH_NOR2X6 U6 ( .A(n24), .B(n4), .Z(n22) );
  HS65_LH_NAND2X7 U7 ( .A(n17), .B(n8), .Z(n10) );
  HS65_LH_NAND2X7 U8 ( .A(n19), .B(n16), .Z(n11) );
  HS65_LH_IVX9 U9 ( .A(n19), .Z(n4) );
  HS65_LH_NOR4ABX2 U10 ( .A(n16), .B(n5), .C(n7), .D(\ctrl_i[OPCODE][2] ), .Z(
        n15) );
  HS65_LH_NOR3AX2 U11 ( .A(n23), .B(\ctrl_i[OPCODE][1] ), .C(
        \ctrl_i[OPCODE][2] ), .Z(n14) );
  HS65_LH_NOR3X4 U12 ( .A(n7), .B(\ctrl_i[OPCODE][2] ), .C(n5), .Z(n19) );
  HS65_LH_NAND3X5 U13 ( .A(n23), .B(\ctrl_i[OPCODE][1] ), .C(
        \ctrl_i[OPCODE][2] ), .Z(n12) );
  HS65_LH_NOR4ABX2 U14 ( .A(n16), .B(n5), .C(\ctrl_i[OPCODE][1] ), .D(
        \ctrl_i[OPCODE][2] ), .Z(n13) );
  HS65_LH_NOR3X4 U15 ( .A(n24), .B(\ctrl_i[OPCODE][3] ), .C(n4), .Z(n17) );
  HS65_LH_NAND3X5 U16 ( .A(n16), .B(n7), .C(\ctrl_i[OPCODE][2] ), .Z(n20) );
  HS65_LH_NOR3AX2 U17 ( .A(\ctrl_i[OPCODE][3] ), .B(n5), .C(
        \ctrl_i[OPCODE][5] ), .Z(n23) );
  HS65_LH_NOR2X6 U18 ( .A(\ctrl_i[OPCODE][5] ), .B(\ctrl_i[OPCODE][3] ), .Z(
        n16) );
  HS65_LH_IVX9 U19 ( .A(\ctrl_i[OPCODE][4] ), .Z(n8) );
  HS65_LH_OAI21X3 U20 ( .A(\ctrl_i[OPCODE][4] ), .B(n11), .C(n6), .Z(
        \ctrl_o[CALU_OP][2] ) );
  HS65_LH_IVX9 U21 ( .A(\ctrl_i[OPCODE][1] ), .Z(n7) );
  HS65_LH_IVX9 U22 ( .A(\ctrl_i[OPCODE][5] ), .Z(n24) );
  HS65_LH_IVX9 U23 ( .A(\ctrl_o[BRANCH] ), .Z(n6) );
  HS65_LH_NOR2X6 U24 ( .A(n20), .B(\ctrl_i[OPCODE][4] ), .Z(\ctrl_o[BRANCH] )
         );
  HS65_LH_IVX9 U25 ( .A(\ctrl_i[OPCODE][0] ), .Z(n5) );
  HS65_LH_OAI21X3 U26 ( .A(\ctrl_i[OPCODE][4] ), .B(n12), .C(n21), .Z(
        \ctrl_o[ALUSRC_B] ) );
  HS65_LH_OAI31X5 U27 ( .A(n20), .B(\ctrl_i[OPCODE][4] ), .C(n5), .D(n21), .Z(
        \ctrl_o[CALU_OP][0] ) );
  HS65_LH_OAI21X3 U28 ( .A(\ctrl_i[OPCODE][4] ), .B(n9), .C(n10), .Z(
        \ctrl_o[REGWRITE] ) );
  HS65_LH_NOR4ABX2 U29 ( .A(n11), .B(n12), .C(n13), .D(n14), .Z(n9) );
  HS65_LH_NAND4ABX3 U30 ( .A(n17), .B(\ctrl_i[OPCODE][2] ), .C(n8), .D(n18), 
        .Z(\ctrl_o[MEMWEN_N] ) );
  HS65_LH_NOR3X4 U31 ( .A(n5), .B(n24), .C(n7), .Z(n18) );
  HS65_LH_CBI4I1X5 U32 ( .A(n3), .B(n12), .C(\ctrl_i[OPCODE][4] ), .D(n6), .Z(
        \ctrl_o[CALU_OP][1] ) );
  HS65_LH_IVX9 U33 ( .A(n15), .Z(n3) );
  HS65_LH_CB4I6X9 U34 ( .A(n13), .B(n15), .C(n8), .D(\ctrl_o[CALU_OP][2] ), 
        .Z(\ctrl_o[REGDST] ) );
  HS65_LH_IVX9 U35 ( .A(n10), .Z(\ctrl_o[MEMTOREG] ) );
endmodule


module pc ( clk, rst_n, halt_i, npc_i, pc_o );
  input [11:0] npc_i;
  output [11:0] pc_o;
  input clk, rst_n, halt_i;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n1;

  HS65_LH_DFPSQX9 \pc_c_reg[11]  ( .D(n13), .CP(clk), .SN(rst_n), .Q(pc_o[11])
         );
  HS65_LH_DFPSQX9 \pc_c_reg[10]  ( .D(n12), .CP(clk), .SN(rst_n), .Q(pc_o[10])
         );
  HS65_LH_DFPSQX9 \pc_c_reg[9]  ( .D(n11), .CP(clk), .SN(rst_n), .Q(pc_o[9])
         );
  HS65_LH_DFPSQX9 \pc_c_reg[8]  ( .D(n10), .CP(clk), .SN(rst_n), .Q(pc_o[8])
         );
  HS65_LH_DFPSQX9 \pc_c_reg[7]  ( .D(n9), .CP(clk), .SN(rst_n), .Q(pc_o[7]) );
  HS65_LH_DFPSQX9 \pc_c_reg[6]  ( .D(n8), .CP(clk), .SN(rst_n), .Q(pc_o[6]) );
  HS65_LH_DFPSQX9 \pc_c_reg[5]  ( .D(n7), .CP(clk), .SN(rst_n), .Q(pc_o[5]) );
  HS65_LH_DFPSQX9 \pc_c_reg[4]  ( .D(n6), .CP(clk), .SN(rst_n), .Q(pc_o[4]) );
  HS65_LH_DFPSQX9 \pc_c_reg[3]  ( .D(n5), .CP(clk), .SN(rst_n), .Q(pc_o[3]) );
  HS65_LH_DFPSQX9 \pc_c_reg[2]  ( .D(n4), .CP(clk), .SN(rst_n), .Q(pc_o[2]) );
  HS65_LH_DFPSQX9 \pc_c_reg[1]  ( .D(n3), .CP(clk), .SN(rst_n), .Q(pc_o[1]) );
  HS65_LH_DFPSQX9 \pc_c_reg[0]  ( .D(n2), .CP(clk), .SN(rst_n), .Q(pc_o[0]) );
  HS65_LH_AO22X9 U2 ( .A(pc_o[9]), .B(halt_i), .C(npc_i[9]), .D(n1), .Z(n11)
         );
  HS65_LH_AO22X9 U3 ( .A(pc_o[0]), .B(halt_i), .C(npc_i[0]), .D(n1), .Z(n2) );
  HS65_LH_AO22X9 U4 ( .A(pc_o[1]), .B(halt_i), .C(npc_i[1]), .D(n1), .Z(n3) );
  HS65_LH_AO22X9 U5 ( .A(pc_o[2]), .B(halt_i), .C(npc_i[2]), .D(n1), .Z(n4) );
  HS65_LH_AO22X9 U6 ( .A(pc_o[3]), .B(halt_i), .C(npc_i[3]), .D(n1), .Z(n5) );
  HS65_LH_AO22X9 U7 ( .A(pc_o[4]), .B(halt_i), .C(npc_i[4]), .D(n1), .Z(n6) );
  HS65_LH_AO22X9 U8 ( .A(pc_o[5]), .B(halt_i), .C(npc_i[5]), .D(n1), .Z(n7) );
  HS65_LH_AO22X9 U9 ( .A(pc_o[6]), .B(halt_i), .C(npc_i[6]), .D(n1), .Z(n8) );
  HS65_LH_AO22X9 U10 ( .A(pc_o[7]), .B(halt_i), .C(npc_i[7]), .D(n1), .Z(n9)
         );
  HS65_LH_AO22X9 U11 ( .A(pc_o[8]), .B(halt_i), .C(npc_i[8]), .D(n1), .Z(n10)
         );
  HS65_LH_AO22X9 U12 ( .A(pc_o[10]), .B(halt_i), .C(npc_i[10]), .D(n1), .Z(n12) );
  HS65_LH_AO22X9 U13 ( .A(pc_o[11]), .B(halt_i), .C(npc_i[11]), .D(n1), .Z(n13) );
  HS65_LH_IVX9 U14 ( .A(halt_i), .Z(n1) );
endmodule


module if_top_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HS65_LH_HA1X4 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .CO(carry[11]), .S0(
        SUM[10]) );
  HS65_LH_HA1X4 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .CO(carry[10]), .S0(SUM[9])
         );
  HS65_LH_HA1X4 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .CO(carry[9]), .S0(SUM[8])
         );
  HS65_LH_HA1X4 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .CO(carry[8]), .S0(SUM[7])
         );
  HS65_LH_HA1X4 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .CO(carry[7]), .S0(SUM[6])
         );
  HS65_LH_HA1X4 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .CO(carry[6]), .S0(SUM[5])
         );
  HS65_LH_HA1X4 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .CO(carry[5]), .S0(SUM[4])
         );
  HS65_LH_HA1X4 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .CO(carry[4]), .S0(SUM[3])
         );
  HS65_LH_HA1X4 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .CO(carry[3]), .S0(SUM[2])
         );
  HS65_LH_HA1X4 U1_1_1 ( .A0(A[1]), .B0(A[0]), .CO(carry[2]), .S0(SUM[1]) );
  HS65_LHS_XOR2X3 U1 ( .A(carry[11]), .B(A[11]), .Z(SUM[11]) );
  HS65_LH_CNIVX3 U2 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module if_top ( clk, rst_n, .if_top_i({\if_top_i[HALT_I] , 
        \if_top_i[BRANCH_PC][11] , \if_top_i[BRANCH_PC][10] , 
        \if_top_i[BRANCH_PC][9] , \if_top_i[BRANCH_PC][8] , 
        \if_top_i[BRANCH_PC][7] , \if_top_i[BRANCH_PC][6] , 
        \if_top_i[BRANCH_PC][5] , \if_top_i[BRANCH_PC][4] , 
        \if_top_i[BRANCH_PC][3] , \if_top_i[BRANCH_PC][2] , 
        \if_top_i[BRANCH_PC][1] , \if_top_i[BRANCH_PC][0] , \if_top_i[PCSRC] }
        ), .if_top_o({\if_top_o[IMEM_ADDR][11] , \if_top_o[IMEM_ADDR][10] , 
        \if_top_o[IMEM_ADDR][9] , \if_top_o[IMEM_ADDR][8] , 
        \if_top_o[IMEM_ADDR][7] , \if_top_o[IMEM_ADDR][6] , 
        \if_top_o[IMEM_ADDR][5] , \if_top_o[IMEM_ADDR][4] , 
        \if_top_o[IMEM_ADDR][3] , \if_top_o[IMEM_ADDR][2] , 
        \if_top_o[IMEM_ADDR][1] , \if_top_o[IMEM_ADDR][0] , 
        \if_top_o[PC_PLUS1][11] , \if_top_o[PC_PLUS1][10] , 
        \if_top_o[PC_PLUS1][9] , \if_top_o[PC_PLUS1][8] , 
        \if_top_o[PC_PLUS1][7] , \if_top_o[PC_PLUS1][6] , 
        \if_top_o[PC_PLUS1][5] , \if_top_o[PC_PLUS1][4] , 
        \if_top_o[PC_PLUS1][3] , \if_top_o[PC_PLUS1][2] , 
        \if_top_o[PC_PLUS1][1] , \if_top_o[PC_PLUS1][0] }) );
  input clk, rst_n, \if_top_i[HALT_I] , \if_top_i[BRANCH_PC][11] ,
         \if_top_i[BRANCH_PC][10] , \if_top_i[BRANCH_PC][9] ,
         \if_top_i[BRANCH_PC][8] , \if_top_i[BRANCH_PC][7] ,
         \if_top_i[BRANCH_PC][6] , \if_top_i[BRANCH_PC][5] ,
         \if_top_i[BRANCH_PC][4] , \if_top_i[BRANCH_PC][3] ,
         \if_top_i[BRANCH_PC][2] , \if_top_i[BRANCH_PC][1] ,
         \if_top_i[BRANCH_PC][0] , \if_top_i[PCSRC] ;
  output \if_top_o[IMEM_ADDR][11] , \if_top_o[IMEM_ADDR][10] ,
         \if_top_o[IMEM_ADDR][9] , \if_top_o[IMEM_ADDR][8] ,
         \if_top_o[IMEM_ADDR][7] , \if_top_o[IMEM_ADDR][6] ,
         \if_top_o[IMEM_ADDR][5] , \if_top_o[IMEM_ADDR][4] ,
         \if_top_o[IMEM_ADDR][3] , \if_top_o[IMEM_ADDR][2] ,
         \if_top_o[IMEM_ADDR][1] , \if_top_o[IMEM_ADDR][0] ,
         \if_top_o[PC_PLUS1][11] , \if_top_o[PC_PLUS1][10] ,
         \if_top_o[PC_PLUS1][9] , \if_top_o[PC_PLUS1][8] ,
         \if_top_o[PC_PLUS1][7] , \if_top_o[PC_PLUS1][6] ,
         \if_top_o[PC_PLUS1][5] , \if_top_o[PC_PLUS1][4] ,
         \if_top_o[PC_PLUS1][3] , \if_top_o[PC_PLUS1][2] ,
         \if_top_o[PC_PLUS1][1] , \if_top_o[PC_PLUS1][0] ;
  wire   n1;
  wire   [11:0] s_npc;

  pc pc_inst ( .clk(clk), .rst_n(rst_n), .halt_i(\if_top_i[HALT_I] ), .npc_i(
        s_npc), .pc_o({\if_top_o[IMEM_ADDR][11] , \if_top_o[IMEM_ADDR][10] , 
        \if_top_o[IMEM_ADDR][9] , \if_top_o[IMEM_ADDR][8] , 
        \if_top_o[IMEM_ADDR][7] , \if_top_o[IMEM_ADDR][6] , 
        \if_top_o[IMEM_ADDR][5] , \if_top_o[IMEM_ADDR][4] , 
        \if_top_o[IMEM_ADDR][3] , \if_top_o[IMEM_ADDR][2] , 
        \if_top_o[IMEM_ADDR][1] , \if_top_o[IMEM_ADDR][0] }) );
  if_top_DW01_inc_0 add_37 ( .A({\if_top_o[IMEM_ADDR][11] , 
        \if_top_o[IMEM_ADDR][10] , \if_top_o[IMEM_ADDR][9] , 
        \if_top_o[IMEM_ADDR][8] , \if_top_o[IMEM_ADDR][7] , 
        \if_top_o[IMEM_ADDR][6] , \if_top_o[IMEM_ADDR][5] , 
        \if_top_o[IMEM_ADDR][4] , \if_top_o[IMEM_ADDR][3] , 
        \if_top_o[IMEM_ADDR][2] , \if_top_o[IMEM_ADDR][1] , 
        \if_top_o[IMEM_ADDR][0] }), .SUM({\if_top_o[PC_PLUS1][11] , 
        \if_top_o[PC_PLUS1][10] , \if_top_o[PC_PLUS1][9] , 
        \if_top_o[PC_PLUS1][8] , \if_top_o[PC_PLUS1][7] , 
        \if_top_o[PC_PLUS1][6] , \if_top_o[PC_PLUS1][5] , 
        \if_top_o[PC_PLUS1][4] , \if_top_o[PC_PLUS1][3] , 
        \if_top_o[PC_PLUS1][2] , \if_top_o[PC_PLUS1][1] , 
        \if_top_o[PC_PLUS1][0] }) );
  HS65_LH_IVX9 U2 ( .A(\if_top_i[PCSRC] ), .Z(n1) );
  HS65_LH_AO22X9 U3 ( .A(\if_top_o[PC_PLUS1][9] ), .B(n1), .C(
        \if_top_i[PCSRC] ), .D(\if_top_i[BRANCH_PC][9] ), .Z(s_npc[9]) );
  HS65_LH_AO22X9 U4 ( .A(\if_top_o[PC_PLUS1][0] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][0] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[0]) );
  HS65_LH_AO22X9 U5 ( .A(\if_top_o[PC_PLUS1][1] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][1] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[1]) );
  HS65_LH_AO22X9 U6 ( .A(\if_top_o[PC_PLUS1][2] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][2] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[2]) );
  HS65_LH_AO22X9 U7 ( .A(\if_top_o[PC_PLUS1][3] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][3] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[3]) );
  HS65_LH_AO22X9 U8 ( .A(\if_top_o[PC_PLUS1][4] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][4] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[4]) );
  HS65_LH_AO22X9 U9 ( .A(\if_top_o[PC_PLUS1][5] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][5] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[5]) );
  HS65_LH_AO22X9 U10 ( .A(\if_top_o[PC_PLUS1][6] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][6] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[6]) );
  HS65_LH_AO22X9 U11 ( .A(\if_top_o[PC_PLUS1][7] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][7] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[7]) );
  HS65_LH_AO22X9 U12 ( .A(\if_top_o[PC_PLUS1][8] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][8] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[8]) );
  HS65_LH_AO22X9 U13 ( .A(\if_top_o[PC_PLUS1][10] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][10] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[10]) );
  HS65_LH_AO22X9 U14 ( .A(\if_top_o[PC_PLUS1][11] ), .B(n1), .C(
        \if_top_i[BRANCH_PC][11] ), .D(\if_top_i[PCSRC] ), .Z(s_npc[11]) );
endmodule


module if_id ( clk, rst_n, halt_i, .IF_ID_i({\IF_ID_i[PC_PLUS1][11] , 
        \IF_ID_i[PC_PLUS1][10] , \IF_ID_i[PC_PLUS1][9] , 
        \IF_ID_i[PC_PLUS1][8] , \IF_ID_i[PC_PLUS1][7] , \IF_ID_i[PC_PLUS1][6] , 
        \IF_ID_i[PC_PLUS1][5] , \IF_ID_i[PC_PLUS1][4] , \IF_ID_i[PC_PLUS1][3] , 
        \IF_ID_i[PC_PLUS1][2] , \IF_ID_i[PC_PLUS1][1] , \IF_ID_i[PC_PLUS1][0] 
        }), .IF_ID_o({\IF_ID_o[PC_PLUS1][11] , \IF_ID_o[PC_PLUS1][10] , 
        \IF_ID_o[PC_PLUS1][9] , \IF_ID_o[PC_PLUS1][8] , \IF_ID_o[PC_PLUS1][7] , 
        \IF_ID_o[PC_PLUS1][6] , \IF_ID_o[PC_PLUS1][5] , \IF_ID_o[PC_PLUS1][4] , 
        \IF_ID_o[PC_PLUS1][3] , \IF_ID_o[PC_PLUS1][2] , \IF_ID_o[PC_PLUS1][1] , 
        \IF_ID_o[PC_PLUS1][0] }) );
  input clk, rst_n, halt_i, \IF_ID_i[PC_PLUS1][11] , \IF_ID_i[PC_PLUS1][10] ,
         \IF_ID_i[PC_PLUS1][9] , \IF_ID_i[PC_PLUS1][8] ,
         \IF_ID_i[PC_PLUS1][7] , \IF_ID_i[PC_PLUS1][6] ,
         \IF_ID_i[PC_PLUS1][5] , \IF_ID_i[PC_PLUS1][4] ,
         \IF_ID_i[PC_PLUS1][3] , \IF_ID_i[PC_PLUS1][2] ,
         \IF_ID_i[PC_PLUS1][1] , \IF_ID_i[PC_PLUS1][0] ;
  output \IF_ID_o[PC_PLUS1][11] , \IF_ID_o[PC_PLUS1][10] ,
         \IF_ID_o[PC_PLUS1][9] , \IF_ID_o[PC_PLUS1][8] ,
         \IF_ID_o[PC_PLUS1][7] , \IF_ID_o[PC_PLUS1][6] ,
         \IF_ID_o[PC_PLUS1][5] , \IF_ID_o[PC_PLUS1][4] ,
         \IF_ID_o[PC_PLUS1][3] , \IF_ID_o[PC_PLUS1][2] ,
         \IF_ID_o[PC_PLUS1][1] , \IF_ID_o[PC_PLUS1][0] ;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n1;

  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][11]  ( .D(n13), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][11] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][10]  ( .D(n12), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][10] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][9]  ( .D(n11), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][9] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][8]  ( .D(n10), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][8] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][7]  ( .D(n9), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][7] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][6]  ( .D(n8), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][6] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][5]  ( .D(n7), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][5] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][4]  ( .D(n6), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][4] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][3]  ( .D(n5), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][3] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][2]  ( .D(n4), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][2] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][1]  ( .D(n3), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][1] ) );
  HS65_LH_DFPRQX9 \if_id_c_reg[PC_PLUS1][0]  ( .D(n2), .CP(clk), .RN(rst_n), 
        .Q(\IF_ID_o[PC_PLUS1][0] ) );
  HS65_LH_AO22X9 U2 ( .A(\IF_ID_o[PC_PLUS1][11] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][11] ), .D(n1), .Z(n13) );
  HS65_LH_AO22X9 U3 ( .A(\IF_ID_o[PC_PLUS1][7] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][7] ), .D(n1), .Z(n9) );
  HS65_LH_AO22X9 U4 ( .A(\IF_ID_o[PC_PLUS1][8] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][8] ), .D(n1), .Z(n10) );
  HS65_LH_AO22X9 U5 ( .A(\IF_ID_o[PC_PLUS1][9] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][9] ), .D(n1), .Z(n11) );
  HS65_LH_AO22X9 U6 ( .A(\IF_ID_o[PC_PLUS1][10] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][10] ), .D(n1), .Z(n12) );
  HS65_LH_AO22X9 U7 ( .A(halt_i), .B(\IF_ID_o[PC_PLUS1][0] ), .C(
        \IF_ID_i[PC_PLUS1][0] ), .D(n1), .Z(n2) );
  HS65_LH_AO22X9 U8 ( .A(\IF_ID_o[PC_PLUS1][1] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][1] ), .D(n1), .Z(n3) );
  HS65_LH_AO22X9 U9 ( .A(\IF_ID_o[PC_PLUS1][2] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][2] ), .D(n1), .Z(n4) );
  HS65_LH_AO22X9 U10 ( .A(\IF_ID_o[PC_PLUS1][3] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][3] ), .D(n1), .Z(n5) );
  HS65_LH_AO22X9 U11 ( .A(\IF_ID_o[PC_PLUS1][4] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][4] ), .D(n1), .Z(n6) );
  HS65_LH_AO22X9 U12 ( .A(\IF_ID_o[PC_PLUS1][5] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][5] ), .D(n1), .Z(n7) );
  HS65_LH_AO22X9 U13 ( .A(\IF_ID_o[PC_PLUS1][6] ), .B(halt_i), .C(
        \IF_ID_i[PC_PLUS1][6] ), .D(n1), .Z(n8) );
  HS65_LH_IVX9 U14 ( .A(halt_i), .Z(n1) );
endmodule


module regfile ( clk, rst_n, .regfile_i({\regfile_i[ADRREAD0][4] , 
        \regfile_i[ADRREAD0][3] , \regfile_i[ADRREAD0][2] , 
        \regfile_i[ADRREAD0][1] , \regfile_i[ADRREAD0][0] , 
        \regfile_i[ADRREAD1][4] , \regfile_i[ADRREAD1][3] , 
        \regfile_i[ADRREAD1][2] , \regfile_i[ADRREAD1][1] , 
        \regfile_i[ADRREAD1][0] , \regfile_i[ADRWRITE][4] , 
        \regfile_i[ADRWRITE][3] , \regfile_i[ADRWRITE][2] , 
        \regfile_i[ADRWRITE][1] , \regfile_i[ADRWRITE][0] , 
        \regfile_i[WRITE_DATA][31] , \regfile_i[WRITE_DATA][30] , 
        \regfile_i[WRITE_DATA][29] , \regfile_i[WRITE_DATA][28] , 
        \regfile_i[WRITE_DATA][27] , \regfile_i[WRITE_DATA][26] , 
        \regfile_i[WRITE_DATA][25] , \regfile_i[WRITE_DATA][24] , 
        \regfile_i[WRITE_DATA][23] , \regfile_i[WRITE_DATA][22] , 
        \regfile_i[WRITE_DATA][21] , \regfile_i[WRITE_DATA][20] , 
        \regfile_i[WRITE_DATA][19] , \regfile_i[WRITE_DATA][18] , 
        \regfile_i[WRITE_DATA][17] , \regfile_i[WRITE_DATA][16] , 
        \regfile_i[WRITE_DATA][15] , \regfile_i[WRITE_DATA][14] , 
        \regfile_i[WRITE_DATA][13] , \regfile_i[WRITE_DATA][12] , 
        \regfile_i[WRITE_DATA][11] , \regfile_i[WRITE_DATA][10] , 
        \regfile_i[WRITE_DATA][9] , \regfile_i[WRITE_DATA][8] , 
        \regfile_i[WRITE_DATA][7] , \regfile_i[WRITE_DATA][6] , 
        \regfile_i[WRITE_DATA][5] , \regfile_i[WRITE_DATA][4] , 
        \regfile_i[WRITE_DATA][3] , \regfile_i[WRITE_DATA][2] , 
        \regfile_i[WRITE_DATA][1] , \regfile_i[WRITE_DATA][0] , 
        \regfile_i[FORWARD_A] , \regfile_i[FORWARD_B] , \regfile_i[WR_EN] }), 
    .regfile_o({\regfile_o[READ_DATA0][31] , \regfile_o[READ_DATA0][30] , 
        \regfile_o[READ_DATA0][29] , \regfile_o[READ_DATA0][28] , 
        \regfile_o[READ_DATA0][27] , \regfile_o[READ_DATA0][26] , 
        \regfile_o[READ_DATA0][25] , \regfile_o[READ_DATA0][24] , 
        \regfile_o[READ_DATA0][23] , \regfile_o[READ_DATA0][22] , 
        \regfile_o[READ_DATA0][21] , \regfile_o[READ_DATA0][20] , 
        \regfile_o[READ_DATA0][19] , \regfile_o[READ_DATA0][18] , 
        \regfile_o[READ_DATA0][17] , \regfile_o[READ_DATA0][16] , 
        \regfile_o[READ_DATA0][15] , \regfile_o[READ_DATA0][14] , 
        \regfile_o[READ_DATA0][13] , \regfile_o[READ_DATA0][12] , 
        \regfile_o[READ_DATA0][11] , \regfile_o[READ_DATA0][10] , 
        \regfile_o[READ_DATA0][9] , \regfile_o[READ_DATA0][8] , 
        \regfile_o[READ_DATA0][7] , \regfile_o[READ_DATA0][6] , 
        \regfile_o[READ_DATA0][5] , \regfile_o[READ_DATA0][4] , 
        \regfile_o[READ_DATA0][3] , \regfile_o[READ_DATA0][2] , 
        \regfile_o[READ_DATA0][1] , \regfile_o[READ_DATA0][0] , 
        \regfile_o[READ_DATA1][31] , \regfile_o[READ_DATA1][30] , 
        \regfile_o[READ_DATA1][29] , \regfile_o[READ_DATA1][28] , 
        \regfile_o[READ_DATA1][27] , \regfile_o[READ_DATA1][26] , 
        \regfile_o[READ_DATA1][25] , \regfile_o[READ_DATA1][24] , 
        \regfile_o[READ_DATA1][23] , \regfile_o[READ_DATA1][22] , 
        \regfile_o[READ_DATA1][21] , \regfile_o[READ_DATA1][20] , 
        \regfile_o[READ_DATA1][19] , \regfile_o[READ_DATA1][18] , 
        \regfile_o[READ_DATA1][17] , \regfile_o[READ_DATA1][16] , 
        \regfile_o[READ_DATA1][15] , \regfile_o[READ_DATA1][14] , 
        \regfile_o[READ_DATA1][13] , \regfile_o[READ_DATA1][12] , 
        \regfile_o[READ_DATA1][11] , \regfile_o[READ_DATA1][10] , 
        \regfile_o[READ_DATA1][9] , \regfile_o[READ_DATA1][8] , 
        \regfile_o[READ_DATA1][7] , \regfile_o[READ_DATA1][6] , 
        \regfile_o[READ_DATA1][5] , \regfile_o[READ_DATA1][4] , 
        \regfile_o[READ_DATA1][3] , \regfile_o[READ_DATA1][2] , 
        \regfile_o[READ_DATA1][1] , \regfile_o[READ_DATA1][0] }) );
  input clk, rst_n, \regfile_i[ADRREAD0][4] , \regfile_i[ADRREAD0][3] ,
         \regfile_i[ADRREAD0][2] , \regfile_i[ADRREAD0][1] ,
         \regfile_i[ADRREAD0][0] , \regfile_i[ADRREAD1][4] ,
         \regfile_i[ADRREAD1][3] , \regfile_i[ADRREAD1][2] ,
         \regfile_i[ADRREAD1][1] , \regfile_i[ADRREAD1][0] ,
         \regfile_i[ADRWRITE][4] , \regfile_i[ADRWRITE][3] ,
         \regfile_i[ADRWRITE][2] , \regfile_i[ADRWRITE][1] ,
         \regfile_i[ADRWRITE][0] , \regfile_i[WRITE_DATA][31] ,
         \regfile_i[WRITE_DATA][30] , \regfile_i[WRITE_DATA][29] ,
         \regfile_i[WRITE_DATA][28] , \regfile_i[WRITE_DATA][27] ,
         \regfile_i[WRITE_DATA][26] , \regfile_i[WRITE_DATA][25] ,
         \regfile_i[WRITE_DATA][24] , \regfile_i[WRITE_DATA][23] ,
         \regfile_i[WRITE_DATA][22] , \regfile_i[WRITE_DATA][21] ,
         \regfile_i[WRITE_DATA][20] , \regfile_i[WRITE_DATA][19] ,
         \regfile_i[WRITE_DATA][18] , \regfile_i[WRITE_DATA][17] ,
         \regfile_i[WRITE_DATA][16] , \regfile_i[WRITE_DATA][15] ,
         \regfile_i[WRITE_DATA][14] , \regfile_i[WRITE_DATA][13] ,
         \regfile_i[WRITE_DATA][12] , \regfile_i[WRITE_DATA][11] ,
         \regfile_i[WRITE_DATA][10] , \regfile_i[WRITE_DATA][9] ,
         \regfile_i[WRITE_DATA][8] , \regfile_i[WRITE_DATA][7] ,
         \regfile_i[WRITE_DATA][6] , \regfile_i[WRITE_DATA][5] ,
         \regfile_i[WRITE_DATA][4] , \regfile_i[WRITE_DATA][3] ,
         \regfile_i[WRITE_DATA][2] , \regfile_i[WRITE_DATA][1] ,
         \regfile_i[WRITE_DATA][0] , \regfile_i[FORWARD_A] ,
         \regfile_i[FORWARD_B] , \regfile_i[WR_EN] ;
  output \regfile_o[READ_DATA0][31] , \regfile_o[READ_DATA0][30] ,
         \regfile_o[READ_DATA0][29] , \regfile_o[READ_DATA0][28] ,
         \regfile_o[READ_DATA0][27] , \regfile_o[READ_DATA0][26] ,
         \regfile_o[READ_DATA0][25] , \regfile_o[READ_DATA0][24] ,
         \regfile_o[READ_DATA0][23] , \regfile_o[READ_DATA0][22] ,
         \regfile_o[READ_DATA0][21] , \regfile_o[READ_DATA0][20] ,
         \regfile_o[READ_DATA0][19] , \regfile_o[READ_DATA0][18] ,
         \regfile_o[READ_DATA0][17] , \regfile_o[READ_DATA0][16] ,
         \regfile_o[READ_DATA0][15] , \regfile_o[READ_DATA0][14] ,
         \regfile_o[READ_DATA0][13] , \regfile_o[READ_DATA0][12] ,
         \regfile_o[READ_DATA0][11] , \regfile_o[READ_DATA0][10] ,
         \regfile_o[READ_DATA0][9] , \regfile_o[READ_DATA0][8] ,
         \regfile_o[READ_DATA0][7] , \regfile_o[READ_DATA0][6] ,
         \regfile_o[READ_DATA0][5] , \regfile_o[READ_DATA0][4] ,
         \regfile_o[READ_DATA0][3] , \regfile_o[READ_DATA0][2] ,
         \regfile_o[READ_DATA0][1] , \regfile_o[READ_DATA0][0] ,
         \regfile_o[READ_DATA1][31] , \regfile_o[READ_DATA1][30] ,
         \regfile_o[READ_DATA1][29] , \regfile_o[READ_DATA1][28] ,
         \regfile_o[READ_DATA1][27] , \regfile_o[READ_DATA1][26] ,
         \regfile_o[READ_DATA1][25] , \regfile_o[READ_DATA1][24] ,
         \regfile_o[READ_DATA1][23] , \regfile_o[READ_DATA1][22] ,
         \regfile_o[READ_DATA1][21] , \regfile_o[READ_DATA1][20] ,
         \regfile_o[READ_DATA1][19] , \regfile_o[READ_DATA1][18] ,
         \regfile_o[READ_DATA1][17] , \regfile_o[READ_DATA1][16] ,
         \regfile_o[READ_DATA1][15] , \regfile_o[READ_DATA1][14] ,
         \regfile_o[READ_DATA1][13] , \regfile_o[READ_DATA1][12] ,
         \regfile_o[READ_DATA1][11] , \regfile_o[READ_DATA1][10] ,
         \regfile_o[READ_DATA1][9] , \regfile_o[READ_DATA1][8] ,
         \regfile_o[READ_DATA1][7] , \regfile_o[READ_DATA1][6] ,
         \regfile_o[READ_DATA1][5] , \regfile_o[READ_DATA1][4] ,
         \regfile_o[READ_DATA1][3] , \regfile_o[READ_DATA1][2] ,
         \regfile_o[READ_DATA1][1] , \regfile_o[READ_DATA1][0] ;
  wire   \registers[31][31] , \registers[31][30] , \registers[31][29] ,
         \registers[31][28] , \registers[31][27] , \registers[31][26] ,
         \registers[31][25] , \registers[31][24] , \registers[31][23] ,
         \registers[31][22] , \registers[31][21] , \registers[31][20] ,
         \registers[31][19] , \registers[31][18] , \registers[31][17] ,
         \registers[31][16] , \registers[31][15] , \registers[31][14] ,
         \registers[31][13] , \registers[31][12] , \registers[31][11] ,
         \registers[31][10] , \registers[31][9] , \registers[31][8] ,
         \registers[31][7] , \registers[31][6] , \registers[31][5] ,
         \registers[31][4] , \registers[31][3] , \registers[31][2] ,
         \registers[31][1] , \registers[31][0] , \registers[30][31] ,
         \registers[30][30] , \registers[30][29] , \registers[30][28] ,
         \registers[30][27] , \registers[30][26] , \registers[30][25] ,
         \registers[30][24] , \registers[30][23] , \registers[30][22] ,
         \registers[30][21] , \registers[30][20] , \registers[30][19] ,
         \registers[30][18] , \registers[30][17] , \registers[30][16] ,
         \registers[30][15] , \registers[30][14] , \registers[30][13] ,
         \registers[30][12] , \registers[30][11] , \registers[30][10] ,
         \registers[30][9] , \registers[30][8] , \registers[30][7] ,
         \registers[30][6] , \registers[30][5] , \registers[30][4] ,
         \registers[30][3] , \registers[30][2] , \registers[30][1] ,
         \registers[30][0] , \registers[25][31] , \registers[25][30] ,
         \registers[25][29] , \registers[25][28] , \registers[25][27] ,
         \registers[25][26] , \registers[25][25] , \registers[25][24] ,
         \registers[25][23] , \registers[25][22] , \registers[25][21] ,
         \registers[25][20] , \registers[25][19] , \registers[25][18] ,
         \registers[25][17] , \registers[25][16] , \registers[25][15] ,
         \registers[25][14] , \registers[25][13] , \registers[25][12] ,
         \registers[25][11] , \registers[25][10] , \registers[25][9] ,
         \registers[25][8] , \registers[25][7] , \registers[25][6] ,
         \registers[25][5] , \registers[25][4] , \registers[25][3] ,
         \registers[25][2] , \registers[25][1] , \registers[25][0] ,
         \registers[24][31] , \registers[24][30] , \registers[24][29] ,
         \registers[24][28] , \registers[24][27] , \registers[24][26] ,
         \registers[24][25] , \registers[24][24] , \registers[24][23] ,
         \registers[24][22] , \registers[24][21] , \registers[24][20] ,
         \registers[24][19] , \registers[24][18] , \registers[24][17] ,
         \registers[24][16] , \registers[24][15] , \registers[24][14] ,
         \registers[24][13] , \registers[24][12] , \registers[24][11] ,
         \registers[24][10] , \registers[24][9] , \registers[24][8] ,
         \registers[24][7] , \registers[24][6] , \registers[24][5] ,
         \registers[24][4] , \registers[24][3] , \registers[24][2] ,
         \registers[24][1] , \registers[24][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[22][31] , \registers[22][30] ,
         \registers[22][29] , \registers[22][28] , \registers[22][27] ,
         \registers[22][26] , \registers[22][25] , \registers[22][24] ,
         \registers[22][23] , \registers[22][22] , \registers[22][21] ,
         \registers[22][20] , \registers[22][19] , \registers[22][18] ,
         \registers[22][17] , \registers[22][16] , \registers[22][15] ,
         \registers[22][14] , \registers[22][13] , \registers[22][12] ,
         \registers[22][11] , \registers[22][10] , \registers[22][9] ,
         \registers[22][8] , \registers[22][7] , \registers[22][6] ,
         \registers[22][5] , \registers[22][4] , \registers[22][3] ,
         \registers[22][2] , \registers[22][1] , \registers[22][0] ,
         \registers[21][31] , \registers[21][30] , \registers[21][29] ,
         \registers[21][28] , \registers[21][27] , \registers[21][26] ,
         \registers[21][25] , \registers[21][24] , \registers[21][23] ,
         \registers[21][22] , \registers[21][21] , \registers[21][20] ,
         \registers[21][19] , \registers[21][18] , \registers[21][17] ,
         \registers[21][16] , \registers[21][15] , \registers[21][14] ,
         \registers[21][13] , \registers[21][12] , \registers[21][11] ,
         \registers[21][10] , \registers[21][9] , \registers[21][8] ,
         \registers[21][7] , \registers[21][6] , \registers[21][5] ,
         \registers[21][4] , \registers[21][3] , \registers[21][2] ,
         \registers[21][1] , \registers[21][0] , \registers[20][31] ,
         \registers[20][30] , \registers[20][29] , \registers[20][28] ,
         \registers[20][27] , \registers[20][26] , \registers[20][25] ,
         \registers[20][24] , \registers[20][23] , \registers[20][22] ,
         \registers[20][21] , \registers[20][20] , \registers[20][19] ,
         \registers[20][18] , \registers[20][17] , \registers[20][16] ,
         \registers[20][15] , \registers[20][14] , \registers[20][13] ,
         \registers[20][12] , \registers[20][11] , \registers[20][10] ,
         \registers[20][9] , \registers[20][8] , \registers[20][7] ,
         \registers[20][6] , \registers[20][5] , \registers[20][4] ,
         \registers[20][3] , \registers[20][2] , \registers[20][1] ,
         \registers[20][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[18][31] , \registers[18][30] , \registers[18][29] ,
         \registers[18][28] , \registers[18][27] , \registers[18][26] ,
         \registers[18][25] , \registers[18][24] , \registers[18][23] ,
         \registers[18][22] , \registers[18][21] , \registers[18][20] ,
         \registers[18][19] , \registers[18][18] , \registers[18][17] ,
         \registers[18][16] , \registers[18][15] , \registers[18][14] ,
         \registers[18][13] , \registers[18][12] , \registers[18][11] ,
         \registers[18][10] , \registers[18][9] , \registers[18][8] ,
         \registers[18][7] , \registers[18][6] , \registers[18][5] ,
         \registers[18][4] , \registers[18][3] , \registers[18][2] ,
         \registers[18][1] , \registers[18][0] , \registers[17][31] ,
         \registers[17][30] , \registers[17][29] , \registers[17][28] ,
         \registers[17][27] , \registers[17][26] , \registers[17][25] ,
         \registers[17][24] , \registers[17][23] , \registers[17][22] ,
         \registers[17][21] , \registers[17][20] , \registers[17][19] ,
         \registers[17][18] , \registers[17][17] , \registers[17][16] ,
         \registers[17][15] , \registers[17][14] , \registers[17][13] ,
         \registers[17][12] , \registers[17][11] , \registers[17][10] ,
         \registers[17][9] , \registers[17][8] , \registers[17][7] ,
         \registers[17][6] , \registers[17][5] , \registers[17][4] ,
         \registers[17][3] , \registers[17][2] , \registers[17][1] ,
         \registers[17][0] , \registers[16][31] , \registers[16][30] ,
         \registers[16][29] , \registers[16][28] , \registers[16][27] ,
         \registers[16][26] , \registers[16][25] , \registers[16][24] ,
         \registers[16][23] , \registers[16][22] , \registers[16][21] ,
         \registers[16][20] , \registers[16][19] , \registers[16][18] ,
         \registers[16][17] , \registers[16][16] , \registers[16][15] ,
         \registers[16][14] , \registers[16][13] , \registers[16][12] ,
         \registers[16][11] , \registers[16][10] , \registers[16][9] ,
         \registers[16][8] , \registers[16][7] , \registers[16][6] ,
         \registers[16][5] , \registers[16][4] , \registers[16][3] ,
         \registers[16][2] , \registers[16][1] , \registers[16][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[12][31] ,
         \registers[12][30] , \registers[12][29] , \registers[12][28] ,
         \registers[12][27] , \registers[12][26] , \registers[12][25] ,
         \registers[12][24] , \registers[12][23] , \registers[12][22] ,
         \registers[12][21] , \registers[12][20] , \registers[12][19] ,
         \registers[12][18] , \registers[12][17] , \registers[12][16] ,
         \registers[12][15] , \registers[12][14] , \registers[12][13] ,
         \registers[12][12] , \registers[12][11] , \registers[12][10] ,
         \registers[12][9] , \registers[12][8] , \registers[12][7] ,
         \registers[12][6] , \registers[12][5] , \registers[12][4] ,
         \registers[12][3] , \registers[12][2] , \registers[12][1] ,
         \registers[12][0] , \registers[11][31] , \registers[11][30] ,
         \registers[11][29] , \registers[11][28] , \registers[11][27] ,
         \registers[11][26] , \registers[11][25] , \registers[11][24] ,
         \registers[11][23] , \registers[11][22] , \registers[11][21] ,
         \registers[11][20] , \registers[11][19] , \registers[11][18] ,
         \registers[11][17] , \registers[11][16] , \registers[11][15] ,
         \registers[11][14] , \registers[11][13] , \registers[11][12] ,
         \registers[11][11] , \registers[11][10] , \registers[11][9] ,
         \registers[11][8] , \registers[11][7] , \registers[11][6] ,
         \registers[11][5] , \registers[11][4] , \registers[11][3] ,
         \registers[11][2] , \registers[11][1] , \registers[11][0] ,
         \registers[10][31] , \registers[10][30] , \registers[10][29] ,
         \registers[10][28] , \registers[10][27] , \registers[10][26] ,
         \registers[10][25] , \registers[10][24] , \registers[10][23] ,
         \registers[10][22] , \registers[10][21] , \registers[10][20] ,
         \registers[10][19] , \registers[10][18] , \registers[10][17] ,
         \registers[10][16] , \registers[10][15] , \registers[10][14] ,
         \registers[10][13] , \registers[10][12] , \registers[10][11] ,
         \registers[10][10] , \registers[10][9] , \registers[10][8] ,
         \registers[10][7] , \registers[10][6] , \registers[10][5] ,
         \registers[10][4] , \registers[10][3] , \registers[10][2] ,
         \registers[10][1] , \registers[10][0] , \registers[7][31] ,
         \registers[7][30] , \registers[7][29] , \registers[7][28] ,
         \registers[7][27] , \registers[7][26] , \registers[7][25] ,
         \registers[7][24] , \registers[7][23] , \registers[7][22] ,
         \registers[7][21] , \registers[7][20] , \registers[7][19] ,
         \registers[7][18] , \registers[7][17] , \registers[7][16] ,
         \registers[7][15] , \registers[7][14] , \registers[7][13] ,
         \registers[7][12] , \registers[7][11] , \registers[7][10] ,
         \registers[7][9] , \registers[7][8] , \registers[7][7] ,
         \registers[7][6] , \registers[7][5] , \registers[7][4] ,
         \registers[7][3] , \registers[7][2] , \registers[7][1] ,
         \registers[7][0] , \registers[6][31] , \registers[6][30] ,
         \registers[6][29] , \registers[6][28] , \registers[6][27] ,
         \registers[6][26] , \registers[6][25] , \registers[6][24] ,
         \registers[6][23] , \registers[6][22] , \registers[6][21] ,
         \registers[6][20] , \registers[6][19] , \registers[6][18] ,
         \registers[6][17] , \registers[6][16] , \registers[6][15] ,
         \registers[6][14] , \registers[6][13] , \registers[6][12] ,
         \registers[6][11] , \registers[6][10] , \registers[6][9] ,
         \registers[6][8] , \registers[6][7] , \registers[6][6] ,
         \registers[6][5] , \registers[6][4] , \registers[6][3] ,
         \registers[6][2] , \registers[6][1] , \registers[6][0] ,
         \registers[5][31] , \registers[5][30] , \registers[5][29] ,
         \registers[5][28] , \registers[5][27] , \registers[5][26] ,
         \registers[5][25] , \registers[5][24] , \registers[5][23] ,
         \registers[5][22] , \registers[5][21] , \registers[5][20] ,
         \registers[5][19] , \registers[5][18] , \registers[5][17] ,
         \registers[5][16] , \registers[5][15] , \registers[5][14] ,
         \registers[5][13] , \registers[5][12] , \registers[5][11] ,
         \registers[5][10] , \registers[5][9] , \registers[5][8] ,
         \registers[5][7] , \registers[5][6] , \registers[5][5] ,
         \registers[5][4] , \registers[5][3] , \registers[5][2] ,
         \registers[5][1] , \registers[5][0] , \registers[4][31] ,
         \registers[4][30] , \registers[4][29] , \registers[4][28] ,
         \registers[4][27] , \registers[4][26] , \registers[4][25] ,
         \registers[4][24] , \registers[4][23] , \registers[4][22] ,
         \registers[4][21] , \registers[4][20] , \registers[4][19] ,
         \registers[4][18] , \registers[4][17] , \registers[4][16] ,
         \registers[4][15] , \registers[4][14] , \registers[4][13] ,
         \registers[4][12] , \registers[4][11] , \registers[4][10] ,
         \registers[4][9] , \registers[4][8] , \registers[4][7] ,
         \registers[4][6] , \registers[4][5] , \registers[4][4] ,
         \registers[4][3] , \registers[4][2] , \registers[4][1] ,
         \registers[4][0] , \registers[3][31] , \registers[3][30] ,
         \registers[3][29] , \registers[3][28] , \registers[3][27] ,
         \registers[3][26] , \registers[3][25] , \registers[3][24] ,
         \registers[3][23] , \registers[3][22] , \registers[3][21] ,
         \registers[3][20] , \registers[3][19] , \registers[3][18] ,
         \registers[3][17] , \registers[3][16] , \registers[3][15] ,
         \registers[3][14] , \registers[3][13] , \registers[3][12] ,
         \registers[3][11] , \registers[3][10] , \registers[3][9] ,
         \registers[3][8] , \registers[3][7] , \registers[3][6] ,
         \registers[3][5] , \registers[3][4] , \registers[3][3] ,
         \registers[3][2] , \registers[3][1] , \registers[3][0] ,
         \registers[2][31] , \registers[2][30] , \registers[2][29] ,
         \registers[2][28] , \registers[2][27] , \registers[2][26] ,
         \registers[2][25] , \registers[2][24] , \registers[2][23] ,
         \registers[2][22] , \registers[2][21] , \registers[2][20] ,
         \registers[2][19] , \registers[2][18] , \registers[2][17] ,
         \registers[2][16] , \registers[2][15] , \registers[2][14] ,
         \registers[2][13] , \registers[2][12] , \registers[2][11] ,
         \registers[2][10] , \registers[2][9] , \registers[2][8] ,
         \registers[2][7] , \registers[2][6] , \registers[2][5] ,
         \registers[2][4] , \registers[2][3] , \registers[2][2] ,
         \registers[2][1] , \registers[2][0] , \registers[1][31] ,
         \registers[1][30] , \registers[1][29] , \registers[1][28] ,
         \registers[1][27] , \registers[1][26] , \registers[1][25] ,
         \registers[1][24] , \registers[1][23] , \registers[1][22] ,
         \registers[1][21] , \registers[1][20] , \registers[1][19] ,
         \registers[1][18] , \registers[1][17] , \registers[1][16] ,
         \registers[1][15] , \registers[1][14] , \registers[1][13] ,
         \registers[1][12] , \registers[1][11] , \registers[1][10] ,
         \registers[1][9] , \registers[1][8] , \registers[1][7] ,
         \registers[1][6] , \registers[1][5] , \registers[1][4] ,
         \registers[1][3] , \registers[1][2] , \registers[1][1] ,
         \registers[1][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1393,
         n1394, n1396, n1398, n1400, n1402, n1404, n1406, n1407, n1408, n1409,
         n1414, n1415, n1416, n1417, n1425, n1426, n1428, n1429, n1430, n1431,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n352, n880, n1392, n1395, n1397, n1399, n1401,
         n1403, n1405, n1410, n1411, n1412, n1413, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1427, n1432, n1433, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099;

  HS65_LH_DFPRQX9 \registers_reg[31][31]  ( .D(n2425), .CP(clk), .RN(n2765), 
        .Q(\registers[31][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][30]  ( .D(n2424), .CP(clk), .RN(n2817), 
        .Q(\registers[31][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][29]  ( .D(n2423), .CP(clk), .RN(n2816), 
        .Q(\registers[31][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][28]  ( .D(n2422), .CP(clk), .RN(n2816), 
        .Q(\registers[31][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][27]  ( .D(n2421), .CP(clk), .RN(n2816), 
        .Q(\registers[31][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][26]  ( .D(n2420), .CP(clk), .RN(n2816), 
        .Q(\registers[31][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][25]  ( .D(n2419), .CP(clk), .RN(n2815), 
        .Q(\registers[31][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][24]  ( .D(n2418), .CP(clk), .RN(n2815), 
        .Q(\registers[31][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][23]  ( .D(n2417), .CP(clk), .RN(n2815), 
        .Q(\registers[31][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][22]  ( .D(n2416), .CP(clk), .RN(n2815), 
        .Q(\registers[31][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][21]  ( .D(n2415), .CP(clk), .RN(n2815), 
        .Q(\registers[31][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][20]  ( .D(n2414), .CP(clk), .RN(n2815), 
        .Q(\registers[31][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][19]  ( .D(n2413), .CP(clk), .RN(n2815), 
        .Q(\registers[31][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][18]  ( .D(n2412), .CP(clk), .RN(n2815), 
        .Q(\registers[31][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][17]  ( .D(n2411), .CP(clk), .RN(n2815), 
        .Q(\registers[31][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][16]  ( .D(n2410), .CP(clk), .RN(n2815), 
        .Q(\registers[31][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][15]  ( .D(n2409), .CP(clk), .RN(n2815), 
        .Q(\registers[31][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][14]  ( .D(n2408), .CP(clk), .RN(n2815), 
        .Q(\registers[31][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][13]  ( .D(n2407), .CP(clk), .RN(n2814), 
        .Q(\registers[31][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][12]  ( .D(n2406), .CP(clk), .RN(n2814), 
        .Q(\registers[31][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][11]  ( .D(n2405), .CP(clk), .RN(n2814), 
        .Q(\registers[31][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][10]  ( .D(n2404), .CP(clk), .RN(n2814), 
        .Q(\registers[31][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][9]  ( .D(n2403), .CP(clk), .RN(n2814), 
        .Q(\registers[31][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][8]  ( .D(n2402), .CP(clk), .RN(n2814), 
        .Q(\registers[31][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][7]  ( .D(n2401), .CP(clk), .RN(n2814), 
        .Q(\registers[31][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][6]  ( .D(n2400), .CP(clk), .RN(n2814), 
        .Q(\registers[31][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][5]  ( .D(n2399), .CP(clk), .RN(n2814), 
        .Q(\registers[31][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][4]  ( .D(n2398), .CP(clk), .RN(n2814), 
        .Q(\registers[31][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][3]  ( .D(n2397), .CP(clk), .RN(n2814), 
        .Q(\registers[31][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][2]  ( .D(n2396), .CP(clk), .RN(n2814), 
        .Q(\registers[31][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][1]  ( .D(n2395), .CP(clk), .RN(n2813), 
        .Q(\registers[31][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[31][0]  ( .D(n2394), .CP(clk), .RN(n2813), 
        .Q(\registers[31][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][31]  ( .D(n2393), .CP(clk), .RN(n2813), 
        .Q(\registers[30][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][30]  ( .D(n2392), .CP(clk), .RN(n2813), 
        .Q(\registers[30][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][29]  ( .D(n2391), .CP(clk), .RN(n2813), 
        .Q(\registers[30][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][28]  ( .D(n2390), .CP(clk), .RN(n2813), 
        .Q(\registers[30][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][27]  ( .D(n2389), .CP(clk), .RN(n2813), 
        .Q(\registers[30][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][26]  ( .D(n2388), .CP(clk), .RN(n2813), 
        .Q(\registers[30][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][25]  ( .D(n2387), .CP(clk), .RN(n2813), 
        .Q(\registers[30][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][24]  ( .D(n2386), .CP(clk), .RN(n2813), 
        .Q(\registers[30][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][23]  ( .D(n2385), .CP(clk), .RN(n2813), 
        .Q(\registers[30][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][22]  ( .D(n2384), .CP(clk), .RN(n2813), 
        .Q(\registers[30][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][21]  ( .D(n2383), .CP(clk), .RN(n2812), 
        .Q(\registers[30][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][20]  ( .D(n2382), .CP(clk), .RN(n2812), 
        .Q(\registers[30][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][19]  ( .D(n2381), .CP(clk), .RN(n2812), 
        .Q(\registers[30][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][18]  ( .D(n2380), .CP(clk), .RN(n2812), 
        .Q(\registers[30][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][17]  ( .D(n2379), .CP(clk), .RN(n2812), 
        .Q(\registers[30][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][16]  ( .D(n2378), .CP(clk), .RN(n2812), 
        .Q(\registers[30][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][15]  ( .D(n2377), .CP(clk), .RN(n2812), 
        .Q(\registers[30][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][14]  ( .D(n2376), .CP(clk), .RN(n2812), 
        .Q(\registers[30][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][13]  ( .D(n2375), .CP(clk), .RN(n2812), 
        .Q(\registers[30][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][12]  ( .D(n2374), .CP(clk), .RN(n2812), 
        .Q(\registers[30][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][11]  ( .D(n2373), .CP(clk), .RN(n2812), 
        .Q(\registers[30][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][10]  ( .D(n2372), .CP(clk), .RN(n2812), 
        .Q(\registers[30][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][9]  ( .D(n2371), .CP(clk), .RN(n2811), 
        .Q(\registers[30][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][8]  ( .D(n2370), .CP(clk), .RN(n2811), 
        .Q(\registers[30][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][7]  ( .D(n2369), .CP(clk), .RN(n2811), 
        .Q(\registers[30][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][6]  ( .D(n2368), .CP(clk), .RN(n2811), 
        .Q(\registers[30][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][5]  ( .D(n2367), .CP(clk), .RN(n2811), 
        .Q(\registers[30][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][4]  ( .D(n2366), .CP(clk), .RN(n2811), 
        .Q(\registers[30][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][3]  ( .D(n2365), .CP(clk), .RN(n2811), 
        .Q(\registers[30][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][2]  ( .D(n2364), .CP(clk), .RN(n2811), 
        .Q(\registers[30][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][1]  ( .D(n2363), .CP(clk), .RN(n2811), 
        .Q(\registers[30][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[30][0]  ( .D(n2362), .CP(clk), .RN(n2811), 
        .Q(\registers[30][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][31]  ( .D(n2233), .CP(clk), .RN(n2811), 
        .Q(\registers[25][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][30]  ( .D(n2232), .CP(clk), .RN(n2811), 
        .Q(\registers[25][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][29]  ( .D(n2231), .CP(clk), .RN(n2810), 
        .Q(\registers[25][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][28]  ( .D(n2230), .CP(clk), .RN(n2810), 
        .Q(\registers[25][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][27]  ( .D(n2229), .CP(clk), .RN(n2810), 
        .Q(\registers[25][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][26]  ( .D(n2228), .CP(clk), .RN(n2810), 
        .Q(\registers[25][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][25]  ( .D(n2227), .CP(clk), .RN(n2810), 
        .Q(\registers[25][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][24]  ( .D(n2226), .CP(clk), .RN(n2810), 
        .Q(\registers[25][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][23]  ( .D(n2225), .CP(clk), .RN(n2810), 
        .Q(\registers[25][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][22]  ( .D(n2224), .CP(clk), .RN(n2810), 
        .Q(\registers[25][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][21]  ( .D(n2223), .CP(clk), .RN(n2810), 
        .Q(\registers[25][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][20]  ( .D(n2222), .CP(clk), .RN(n2810), 
        .Q(\registers[25][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][19]  ( .D(n2221), .CP(clk), .RN(n2810), 
        .Q(\registers[25][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][18]  ( .D(n2220), .CP(clk), .RN(n2810), 
        .Q(\registers[25][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][17]  ( .D(n2219), .CP(clk), .RN(n2809), 
        .Q(\registers[25][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][16]  ( .D(n2218), .CP(clk), .RN(n2809), 
        .Q(\registers[25][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][15]  ( .D(n2217), .CP(clk), .RN(n2809), 
        .Q(\registers[25][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][14]  ( .D(n2216), .CP(clk), .RN(n2809), 
        .Q(\registers[25][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][13]  ( .D(n2215), .CP(clk), .RN(n2809), 
        .Q(\registers[25][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][12]  ( .D(n2214), .CP(clk), .RN(n2809), 
        .Q(\registers[25][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][11]  ( .D(n2213), .CP(clk), .RN(n2809), 
        .Q(\registers[25][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][10]  ( .D(n2212), .CP(clk), .RN(n2809), 
        .Q(\registers[25][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][9]  ( .D(n2211), .CP(clk), .RN(n2809), 
        .Q(\registers[25][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][8]  ( .D(n2210), .CP(clk), .RN(n2809), 
        .Q(\registers[25][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][7]  ( .D(n2209), .CP(clk), .RN(n2809), 
        .Q(\registers[25][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][6]  ( .D(n2208), .CP(clk), .RN(n2809), 
        .Q(\registers[25][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][5]  ( .D(n2207), .CP(clk), .RN(n2808), 
        .Q(\registers[25][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][4]  ( .D(n2206), .CP(clk), .RN(n2808), 
        .Q(\registers[25][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][3]  ( .D(n2205), .CP(clk), .RN(n2808), 
        .Q(\registers[25][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][2]  ( .D(n2204), .CP(clk), .RN(n2808), 
        .Q(\registers[25][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][1]  ( .D(n2203), .CP(clk), .RN(n2808), 
        .Q(\registers[25][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[25][0]  ( .D(n2202), .CP(clk), .RN(n2808), 
        .Q(\registers[25][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][31]  ( .D(n2201), .CP(clk), .RN(n2808), 
        .Q(\registers[24][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][30]  ( .D(n2200), .CP(clk), .RN(n2808), 
        .Q(\registers[24][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][29]  ( .D(n2199), .CP(clk), .RN(n2808), 
        .Q(\registers[24][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][28]  ( .D(n2198), .CP(clk), .RN(n2808), 
        .Q(\registers[24][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][27]  ( .D(n2197), .CP(clk), .RN(n2808), 
        .Q(\registers[24][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][26]  ( .D(n2196), .CP(clk), .RN(n2807), 
        .Q(\registers[24][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][25]  ( .D(n2195), .CP(clk), .RN(n2807), 
        .Q(\registers[24][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][24]  ( .D(n2194), .CP(clk), .RN(n2807), 
        .Q(\registers[24][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][23]  ( .D(n2193), .CP(clk), .RN(n2807), 
        .Q(\registers[24][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][22]  ( .D(n2192), .CP(clk), .RN(n2807), 
        .Q(\registers[24][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][21]  ( .D(n2191), .CP(clk), .RN(n2807), 
        .Q(\registers[24][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][20]  ( .D(n2190), .CP(clk), .RN(n2807), 
        .Q(\registers[24][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][19]  ( .D(n2189), .CP(clk), .RN(n2807), 
        .Q(\registers[24][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][18]  ( .D(n2188), .CP(clk), .RN(n2807), 
        .Q(\registers[24][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][17]  ( .D(n2187), .CP(clk), .RN(n2807), 
        .Q(\registers[24][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][16]  ( .D(n2186), .CP(clk), .RN(n2807), 
        .Q(\registers[24][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][15]  ( .D(n2185), .CP(clk), .RN(n2807), 
        .Q(\registers[24][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][14]  ( .D(n2184), .CP(clk), .RN(n2806), 
        .Q(\registers[24][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][13]  ( .D(n2183), .CP(clk), .RN(n2806), 
        .Q(\registers[24][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][12]  ( .D(n2182), .CP(clk), .RN(n2806), 
        .Q(\registers[24][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][11]  ( .D(n2181), .CP(clk), .RN(n2806), 
        .Q(\registers[24][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][10]  ( .D(n2180), .CP(clk), .RN(n2806), 
        .Q(\registers[24][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][9]  ( .D(n2179), .CP(clk), .RN(n2806), 
        .Q(\registers[24][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][8]  ( .D(n2178), .CP(clk), .RN(n2806), 
        .Q(\registers[24][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][7]  ( .D(n2177), .CP(clk), .RN(n2806), 
        .Q(\registers[24][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][6]  ( .D(n2176), .CP(clk), .RN(n2806), 
        .Q(\registers[24][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][5]  ( .D(n2175), .CP(clk), .RN(n2806), 
        .Q(\registers[24][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][4]  ( .D(n2174), .CP(clk), .RN(n2806), 
        .Q(\registers[24][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][3]  ( .D(n2173), .CP(clk), .RN(n2806), 
        .Q(\registers[24][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][2]  ( .D(n2172), .CP(clk), .RN(n2805), 
        .Q(\registers[24][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][1]  ( .D(n2171), .CP(clk), .RN(n2805), 
        .Q(\registers[24][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[24][0]  ( .D(n2170), .CP(clk), .RN(n2805), 
        .Q(\registers[24][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][31]  ( .D(n2169), .CP(clk), .RN(n2805), 
        .Q(\registers[23][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][30]  ( .D(n2168), .CP(clk), .RN(n2805), 
        .Q(\registers[23][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][29]  ( .D(n2167), .CP(clk), .RN(n2805), 
        .Q(\registers[23][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][28]  ( .D(n2166), .CP(clk), .RN(n2805), 
        .Q(\registers[23][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][27]  ( .D(n2165), .CP(clk), .RN(n2805), 
        .Q(\registers[23][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][26]  ( .D(n2164), .CP(clk), .RN(n2805), 
        .Q(\registers[23][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][25]  ( .D(n2163), .CP(clk), .RN(n2805), 
        .Q(\registers[23][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][24]  ( .D(n2162), .CP(clk), .RN(n2805), 
        .Q(\registers[23][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][23]  ( .D(n2161), .CP(clk), .RN(n2805), 
        .Q(\registers[23][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][22]  ( .D(n2160), .CP(clk), .RN(n2804), 
        .Q(\registers[23][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][21]  ( .D(n2159), .CP(clk), .RN(n2804), 
        .Q(\registers[23][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][20]  ( .D(n2158), .CP(clk), .RN(n2804), 
        .Q(\registers[23][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][19]  ( .D(n2157), .CP(clk), .RN(n2804), 
        .Q(\registers[23][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][18]  ( .D(n2156), .CP(clk), .RN(n2804), 
        .Q(\registers[23][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][17]  ( .D(n2155), .CP(clk), .RN(n2804), 
        .Q(\registers[23][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][16]  ( .D(n2154), .CP(clk), .RN(n2804), 
        .Q(\registers[23][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][15]  ( .D(n2153), .CP(clk), .RN(n2804), 
        .Q(\registers[23][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][14]  ( .D(n2152), .CP(clk), .RN(n2804), 
        .Q(\registers[23][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][13]  ( .D(n2151), .CP(clk), .RN(n2804), 
        .Q(\registers[23][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][12]  ( .D(n2150), .CP(clk), .RN(n2804), 
        .Q(\registers[23][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][11]  ( .D(n2149), .CP(clk), .RN(n2804), 
        .Q(\registers[23][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][10]  ( .D(n2148), .CP(clk), .RN(n2803), 
        .Q(\registers[23][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][9]  ( .D(n2147), .CP(clk), .RN(n2803), 
        .Q(\registers[23][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][8]  ( .D(n2146), .CP(clk), .RN(n2803), 
        .Q(\registers[23][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][7]  ( .D(n2145), .CP(clk), .RN(n2803), 
        .Q(\registers[23][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][6]  ( .D(n2144), .CP(clk), .RN(n2803), 
        .Q(\registers[23][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][5]  ( .D(n2143), .CP(clk), .RN(n2803), 
        .Q(\registers[23][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][4]  ( .D(n2142), .CP(clk), .RN(n2803), 
        .Q(\registers[23][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][3]  ( .D(n2141), .CP(clk), .RN(n2803), 
        .Q(\registers[23][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][2]  ( .D(n2140), .CP(clk), .RN(n2803), 
        .Q(\registers[23][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][1]  ( .D(n2139), .CP(clk), .RN(n2803), 
        .Q(\registers[23][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[23][0]  ( .D(n2138), .CP(clk), .RN(n2803), 
        .Q(\registers[23][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][31]  ( .D(n2137), .CP(clk), .RN(n2803), 
        .Q(\registers[22][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][30]  ( .D(n2136), .CP(clk), .RN(n2802), 
        .Q(\registers[22][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][29]  ( .D(n2135), .CP(clk), .RN(n2802), 
        .Q(\registers[22][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][28]  ( .D(n2134), .CP(clk), .RN(n2802), 
        .Q(\registers[22][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][27]  ( .D(n2133), .CP(clk), .RN(n2802), 
        .Q(\registers[22][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][26]  ( .D(n2132), .CP(clk), .RN(n2802), 
        .Q(\registers[22][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][25]  ( .D(n2131), .CP(clk), .RN(n2802), 
        .Q(\registers[22][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][24]  ( .D(n2130), .CP(clk), .RN(n2802), 
        .Q(\registers[22][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][23]  ( .D(n2129), .CP(clk), .RN(n2802), 
        .Q(\registers[22][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][22]  ( .D(n2128), .CP(clk), .RN(n2802), 
        .Q(\registers[22][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][21]  ( .D(n2127), .CP(clk), .RN(n2802), 
        .Q(\registers[22][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][20]  ( .D(n2126), .CP(clk), .RN(n2802), 
        .Q(\registers[22][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][19]  ( .D(n2125), .CP(clk), .RN(n2802), 
        .Q(\registers[22][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][18]  ( .D(n2124), .CP(clk), .RN(n2801), 
        .Q(\registers[22][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][17]  ( .D(n2123), .CP(clk), .RN(n2801), 
        .Q(\registers[22][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][16]  ( .D(n2122), .CP(clk), .RN(n2801), 
        .Q(\registers[22][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][15]  ( .D(n2121), .CP(clk), .RN(n2801), 
        .Q(\registers[22][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][14]  ( .D(n2120), .CP(clk), .RN(n2801), 
        .Q(\registers[22][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][13]  ( .D(n2119), .CP(clk), .RN(n2801), 
        .Q(\registers[22][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][12]  ( .D(n2118), .CP(clk), .RN(n2801), 
        .Q(\registers[22][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][11]  ( .D(n2117), .CP(clk), .RN(n2801), 
        .Q(\registers[22][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][10]  ( .D(n2116), .CP(clk), .RN(n2801), 
        .Q(\registers[22][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][9]  ( .D(n2115), .CP(clk), .RN(n2801), 
        .Q(\registers[22][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][8]  ( .D(n2114), .CP(clk), .RN(n2801), 
        .Q(\registers[22][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][7]  ( .D(n2113), .CP(clk), .RN(n2808), 
        .Q(\registers[22][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][6]  ( .D(n2112), .CP(clk), .RN(n2825), 
        .Q(\registers[22][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][5]  ( .D(n2111), .CP(clk), .RN(n2825), 
        .Q(\registers[22][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][4]  ( .D(n2110), .CP(clk), .RN(n2825), 
        .Q(\registers[22][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][3]  ( .D(n2109), .CP(clk), .RN(n2825), 
        .Q(\registers[22][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][2]  ( .D(n2108), .CP(clk), .RN(n2825), 
        .Q(\registers[22][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][1]  ( .D(n2107), .CP(clk), .RN(n2825), 
        .Q(\registers[22][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[22][0]  ( .D(n2106), .CP(clk), .RN(n2825), 
        .Q(\registers[22][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][31]  ( .D(n2105), .CP(clk), .RN(n2825), 
        .Q(\registers[21][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][30]  ( .D(n2104), .CP(clk), .RN(n2826), 
        .Q(\registers[21][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][29]  ( .D(n2103), .CP(clk), .RN(n2825), 
        .Q(\registers[21][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][28]  ( .D(n2102), .CP(clk), .RN(n2826), 
        .Q(\registers[21][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][27]  ( .D(n2101), .CP(clk), .RN(n2825), 
        .Q(\registers[21][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][26]  ( .D(n2100), .CP(clk), .RN(n2826), 
        .Q(\registers[21][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][25]  ( .D(n2099), .CP(clk), .RN(n2825), 
        .Q(\registers[21][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][24]  ( .D(n2098), .CP(clk), .RN(n2826), 
        .Q(\registers[21][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][23]  ( .D(n2097), .CP(clk), .RN(n2825), 
        .Q(\registers[21][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][22]  ( .D(n2096), .CP(clk), .RN(n2824), 
        .Q(\registers[21][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][21]  ( .D(n2095), .CP(clk), .RN(n2824), 
        .Q(\registers[21][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][20]  ( .D(n2094), .CP(clk), .RN(n2824), 
        .Q(\registers[21][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][19]  ( .D(n2093), .CP(clk), .RN(n2824), 
        .Q(\registers[21][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][18]  ( .D(n2092), .CP(clk), .RN(n2824), 
        .Q(\registers[21][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][17]  ( .D(n2091), .CP(clk), .RN(n2824), 
        .Q(\registers[21][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][16]  ( .D(n2090), .CP(clk), .RN(n2824), 
        .Q(\registers[21][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][15]  ( .D(n2089), .CP(clk), .RN(n2824), 
        .Q(\registers[21][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][14]  ( .D(n2088), .CP(clk), .RN(n2824), 
        .Q(\registers[21][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][13]  ( .D(n2087), .CP(clk), .RN(n2824), 
        .Q(\registers[21][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][12]  ( .D(n2086), .CP(clk), .RN(n2824), 
        .Q(\registers[21][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][11]  ( .D(n2085), .CP(clk), .RN(n2824), 
        .Q(\registers[21][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][10]  ( .D(n2084), .CP(clk), .RN(n2823), 
        .Q(\registers[21][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][9]  ( .D(n2083), .CP(clk), .RN(n2823), 
        .Q(\registers[21][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][8]  ( .D(n2082), .CP(clk), .RN(n2823), 
        .Q(\registers[21][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][7]  ( .D(n2081), .CP(clk), .RN(n2823), 
        .Q(\registers[21][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][6]  ( .D(n2080), .CP(clk), .RN(n2823), 
        .Q(\registers[21][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][5]  ( .D(n2079), .CP(clk), .RN(n2823), 
        .Q(\registers[21][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][4]  ( .D(n2078), .CP(clk), .RN(n2823), 
        .Q(\registers[21][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][3]  ( .D(n2077), .CP(clk), .RN(n2823), 
        .Q(\registers[21][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][2]  ( .D(n2076), .CP(clk), .RN(n2823), 
        .Q(\registers[21][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][1]  ( .D(n2075), .CP(clk), .RN(n2823), 
        .Q(\registers[21][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[21][0]  ( .D(n2074), .CP(clk), .RN(n2823), 
        .Q(\registers[21][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][31]  ( .D(n2073), .CP(clk), .RN(n2823), 
        .Q(\registers[20][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][30]  ( .D(n2072), .CP(clk), .RN(n2816), 
        .Q(\registers[20][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][29]  ( .D(n2071), .CP(clk), .RN(n2816), 
        .Q(\registers[20][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][28]  ( .D(n2070), .CP(clk), .RN(n2816), 
        .Q(\registers[20][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][27]  ( .D(n2069), .CP(clk), .RN(n2816), 
        .Q(\registers[20][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][26]  ( .D(n2068), .CP(clk), .RN(n2816), 
        .Q(\registers[20][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][25]  ( .D(n2067), .CP(clk), .RN(n2816), 
        .Q(\registers[20][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][24]  ( .D(n2066), .CP(clk), .RN(n2816), 
        .Q(\registers[20][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][23]  ( .D(n2065), .CP(clk), .RN(n2816), 
        .Q(\registers[20][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][22]  ( .D(n2064), .CP(clk), .RN(n2817), 
        .Q(\registers[20][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][21]  ( .D(n2063), .CP(clk), .RN(n2821), 
        .Q(\registers[20][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][20]  ( .D(n2062), .CP(clk), .RN(n2817), 
        .Q(\registers[20][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][19]  ( .D(n2061), .CP(clk), .RN(n2817), 
        .Q(\registers[20][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][18]  ( .D(n2060), .CP(clk), .RN(n2817), 
        .Q(\registers[20][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][17]  ( .D(n2059), .CP(clk), .RN(n2817), 
        .Q(\registers[20][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][16]  ( .D(n2058), .CP(clk), .RN(n2817), 
        .Q(\registers[20][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][15]  ( .D(n2057), .CP(clk), .RN(n2817), 
        .Q(\registers[20][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][14]  ( .D(n2056), .CP(clk), .RN(n2817), 
        .Q(\registers[20][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][13]  ( .D(n2055), .CP(clk), .RN(n2817), 
        .Q(\registers[20][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][12]  ( .D(n2054), .CP(clk), .RN(n2817), 
        .Q(\registers[20][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][11]  ( .D(n2053), .CP(clk), .RN(n2817), 
        .Q(\registers[20][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][10]  ( .D(n2052), .CP(clk), .RN(n2818), 
        .Q(\registers[20][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][9]  ( .D(n2051), .CP(clk), .RN(n2818), 
        .Q(\registers[20][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][8]  ( .D(n2050), .CP(clk), .RN(n2818), 
        .Q(\registers[20][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][7]  ( .D(n2049), .CP(clk), .RN(n2818), 
        .Q(\registers[20][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][6]  ( .D(n2048), .CP(clk), .RN(n2818), 
        .Q(\registers[20][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][5]  ( .D(n2047), .CP(clk), .RN(n2818), 
        .Q(\registers[20][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][4]  ( .D(n2046), .CP(clk), .RN(n2818), 
        .Q(\registers[20][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][3]  ( .D(n2045), .CP(clk), .RN(n2818), 
        .Q(\registers[20][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][2]  ( .D(n2044), .CP(clk), .RN(n2818), 
        .Q(\registers[20][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][1]  ( .D(n2043), .CP(clk), .RN(n2818), 
        .Q(\registers[20][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[20][0]  ( .D(n2042), .CP(clk), .RN(n2818), 
        .Q(\registers[20][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][31]  ( .D(n2041), .CP(clk), .RN(n2819), 
        .Q(\registers[19][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][30]  ( .D(n2040), .CP(clk), .RN(n2819), 
        .Q(\registers[19][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][29]  ( .D(n2039), .CP(clk), .RN(n2819), 
        .Q(\registers[19][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][28]  ( .D(n2038), .CP(clk), .RN(n2819), 
        .Q(\registers[19][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][27]  ( .D(n2037), .CP(clk), .RN(n2819), 
        .Q(\registers[19][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][26]  ( .D(n2036), .CP(clk), .RN(n2819), 
        .Q(\registers[19][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][25]  ( .D(n2035), .CP(clk), .RN(n2819), 
        .Q(\registers[19][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][24]  ( .D(n2034), .CP(clk), .RN(n2819), 
        .Q(\registers[19][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][23]  ( .D(n2033), .CP(clk), .RN(n2819), 
        .Q(\registers[19][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][22]  ( .D(n2032), .CP(clk), .RN(n2819), 
        .Q(\registers[19][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][21]  ( .D(n2031), .CP(clk), .RN(n2819), 
        .Q(\registers[19][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][20]  ( .D(n2030), .CP(clk), .RN(n2819), 
        .Q(\registers[19][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][19]  ( .D(n2029), .CP(clk), .RN(n2820), 
        .Q(\registers[19][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][18]  ( .D(n2028), .CP(clk), .RN(n2820), 
        .Q(\registers[19][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][17]  ( .D(n2027), .CP(clk), .RN(n2820), 
        .Q(\registers[19][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][16]  ( .D(n2026), .CP(clk), .RN(n2820), 
        .Q(\registers[19][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][15]  ( .D(n2025), .CP(clk), .RN(n2820), 
        .Q(\registers[19][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][14]  ( .D(n2024), .CP(clk), .RN(n2820), 
        .Q(\registers[19][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][13]  ( .D(n2023), .CP(clk), .RN(n2820), 
        .Q(\registers[19][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][12]  ( .D(n2022), .CP(clk), .RN(n2820), 
        .Q(\registers[19][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][11]  ( .D(n2021), .CP(clk), .RN(n2820), 
        .Q(\registers[19][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][10]  ( .D(n2020), .CP(clk), .RN(n2820), 
        .Q(\registers[19][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][9]  ( .D(n2019), .CP(clk), .RN(n2820), 
        .Q(\registers[19][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][8]  ( .D(n2018), .CP(clk), .RN(n2820), 
        .Q(\registers[19][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][7]  ( .D(n2017), .CP(clk), .RN(n2821), 
        .Q(\registers[19][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][6]  ( .D(n2016), .CP(clk), .RN(n2821), 
        .Q(\registers[19][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][5]  ( .D(n2015), .CP(clk), .RN(n2821), 
        .Q(\registers[19][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][4]  ( .D(n2014), .CP(clk), .RN(n2821), 
        .Q(\registers[19][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][3]  ( .D(n2013), .CP(clk), .RN(n2821), 
        .Q(\registers[19][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][2]  ( .D(n2012), .CP(clk), .RN(n2821), 
        .Q(\registers[19][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][1]  ( .D(n2011), .CP(clk), .RN(n2821), 
        .Q(\registers[19][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[19][0]  ( .D(n2010), .CP(clk), .RN(n2821), 
        .Q(\registers[19][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][31]  ( .D(n2009), .CP(clk), .RN(n2821), 
        .Q(\registers[18][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][30]  ( .D(n2008), .CP(clk), .RN(n2821), 
        .Q(\registers[18][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][29]  ( .D(n2007), .CP(clk), .RN(n2821), 
        .Q(\registers[18][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][28]  ( .D(n2006), .CP(clk), .RN(n2822), 
        .Q(\registers[18][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][27]  ( .D(n2005), .CP(clk), .RN(n2822), 
        .Q(\registers[18][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][26]  ( .D(n2004), .CP(clk), .RN(n2822), 
        .Q(\registers[18][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][25]  ( .D(n2003), .CP(clk), .RN(n2822), 
        .Q(\registers[18][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][24]  ( .D(n2002), .CP(clk), .RN(n2822), 
        .Q(\registers[18][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][23]  ( .D(n2001), .CP(clk), .RN(n2822), 
        .Q(\registers[18][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][22]  ( .D(n2000), .CP(clk), .RN(n2822), 
        .Q(\registers[18][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][21]  ( .D(n1999), .CP(clk), .RN(n2822), 
        .Q(\registers[18][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][20]  ( .D(n1998), .CP(clk), .RN(n2822), 
        .Q(\registers[18][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][19]  ( .D(n1997), .CP(clk), .RN(n2822), 
        .Q(\registers[18][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][18]  ( .D(n1996), .CP(clk), .RN(n2822), 
        .Q(\registers[18][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][17]  ( .D(n1995), .CP(clk), .RN(n2822), 
        .Q(\registers[18][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][16]  ( .D(n1994), .CP(clk), .RN(n2818), 
        .Q(\registers[18][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][15]  ( .D(n1993), .CP(clk), .RN(n2783), 
        .Q(\registers[18][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][14]  ( .D(n1992), .CP(clk), .RN(n2778), 
        .Q(\registers[18][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][13]  ( .D(n1991), .CP(clk), .RN(n2774), 
        .Q(\registers[18][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][12]  ( .D(n1990), .CP(clk), .RN(n2774), 
        .Q(\registers[18][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][11]  ( .D(n1989), .CP(clk), .RN(n2774), 
        .Q(\registers[18][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][10]  ( .D(n1988), .CP(clk), .RN(n2774), 
        .Q(\registers[18][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][9]  ( .D(n1987), .CP(clk), .RN(n2774), 
        .Q(\registers[18][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][8]  ( .D(n1986), .CP(clk), .RN(n2774), 
        .Q(\registers[18][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][7]  ( .D(n1985), .CP(clk), .RN(n2774), 
        .Q(\registers[18][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][6]  ( .D(n1984), .CP(clk), .RN(n2774), 
        .Q(\registers[18][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][5]  ( .D(n1983), .CP(clk), .RN(n2774), 
        .Q(\registers[18][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][4]  ( .D(n1982), .CP(clk), .RN(n2774), 
        .Q(\registers[18][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][3]  ( .D(n1981), .CP(clk), .RN(n2774), 
        .Q(\registers[18][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][2]  ( .D(n1980), .CP(clk), .RN(n2775), 
        .Q(\registers[18][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][1]  ( .D(n1979), .CP(clk), .RN(n2775), 
        .Q(\registers[18][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[18][0]  ( .D(n1978), .CP(clk), .RN(n2775), 
        .Q(\registers[18][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][31]  ( .D(n1977), .CP(clk), .RN(n2775), 
        .Q(\registers[17][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][30]  ( .D(n1976), .CP(clk), .RN(n2775), 
        .Q(\registers[17][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][29]  ( .D(n1975), .CP(clk), .RN(n2775), 
        .Q(\registers[17][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][28]  ( .D(n1974), .CP(clk), .RN(n2775), 
        .Q(\registers[17][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][27]  ( .D(n1973), .CP(clk), .RN(n2775), 
        .Q(\registers[17][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][26]  ( .D(n1972), .CP(clk), .RN(n2775), 
        .Q(\registers[17][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][25]  ( .D(n1971), .CP(clk), .RN(n2775), 
        .Q(\registers[17][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][24]  ( .D(n1970), .CP(clk), .RN(n2775), 
        .Q(\registers[17][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][23]  ( .D(n1969), .CP(clk), .RN(n2775), 
        .Q(\registers[17][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][22]  ( .D(n1968), .CP(clk), .RN(n2776), 
        .Q(\registers[17][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][21]  ( .D(n1967), .CP(clk), .RN(n2776), 
        .Q(\registers[17][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][20]  ( .D(n1966), .CP(clk), .RN(n2776), 
        .Q(\registers[17][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][19]  ( .D(n1965), .CP(clk), .RN(n2776), 
        .Q(\registers[17][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][18]  ( .D(n1964), .CP(clk), .RN(n2776), 
        .Q(\registers[17][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][17]  ( .D(n1963), .CP(clk), .RN(n2776), 
        .Q(\registers[17][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][16]  ( .D(n1962), .CP(clk), .RN(n2776), 
        .Q(\registers[17][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][15]  ( .D(n1961), .CP(clk), .RN(n2776), 
        .Q(\registers[17][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][14]  ( .D(n1960), .CP(clk), .RN(n2776), 
        .Q(\registers[17][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][13]  ( .D(n1959), .CP(clk), .RN(n2776), 
        .Q(\registers[17][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][12]  ( .D(n1958), .CP(clk), .RN(n2776), 
        .Q(\registers[17][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][11]  ( .D(n1957), .CP(clk), .RN(n2776), 
        .Q(\registers[17][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][10]  ( .D(n1956), .CP(clk), .RN(n2777), 
        .Q(\registers[17][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][9]  ( .D(n1955), .CP(clk), .RN(n2777), 
        .Q(\registers[17][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][8]  ( .D(n1954), .CP(clk), .RN(n2777), 
        .Q(\registers[17][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][7]  ( .D(n1953), .CP(clk), .RN(n2777), 
        .Q(\registers[17][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][6]  ( .D(n1952), .CP(clk), .RN(n2777), 
        .Q(\registers[17][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][5]  ( .D(n1951), .CP(clk), .RN(n2777), 
        .Q(\registers[17][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][4]  ( .D(n1950), .CP(clk), .RN(n2777), 
        .Q(\registers[17][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][3]  ( .D(n1949), .CP(clk), .RN(n2777), 
        .Q(\registers[17][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][2]  ( .D(n1948), .CP(clk), .RN(n2777), 
        .Q(\registers[17][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][1]  ( .D(n1947), .CP(clk), .RN(n2777), 
        .Q(\registers[17][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[17][0]  ( .D(n1946), .CP(clk), .RN(n2777), 
        .Q(\registers[17][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][31]  ( .D(n1945), .CP(clk), .RN(n2777), 
        .Q(\registers[16][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][30]  ( .D(n1944), .CP(clk), .RN(n2778), 
        .Q(\registers[16][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][29]  ( .D(n1943), .CP(clk), .RN(n2778), 
        .Q(\registers[16][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][28]  ( .D(n1942), .CP(clk), .RN(n2778), 
        .Q(\registers[16][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][27]  ( .D(n1941), .CP(clk), .RN(n2778), 
        .Q(\registers[16][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][26]  ( .D(n1940), .CP(clk), .RN(n2778), 
        .Q(\registers[16][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][25]  ( .D(n1939), .CP(clk), .RN(n2778), 
        .Q(\registers[16][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][24]  ( .D(n1938), .CP(clk), .RN(n2778), 
        .Q(\registers[16][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][23]  ( .D(n1937), .CP(clk), .RN(n2778), 
        .Q(\registers[16][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][22]  ( .D(n1936), .CP(clk), .RN(n2778), 
        .Q(\registers[16][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][21]  ( .D(n1935), .CP(clk), .RN(n2778), 
        .Q(\registers[16][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][20]  ( .D(n1934), .CP(clk), .RN(n2778), 
        .Q(\registers[16][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][19]  ( .D(n1933), .CP(clk), .RN(n2779), 
        .Q(\registers[16][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][18]  ( .D(n1932), .CP(clk), .RN(n2779), 
        .Q(\registers[16][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][17]  ( .D(n1931), .CP(clk), .RN(n2779), 
        .Q(\registers[16][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][16]  ( .D(n1930), .CP(clk), .RN(n2779), 
        .Q(\registers[16][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][15]  ( .D(n1929), .CP(clk), .RN(n2779), 
        .Q(\registers[16][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][14]  ( .D(n1928), .CP(clk), .RN(n2779), 
        .Q(\registers[16][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][13]  ( .D(n1927), .CP(clk), .RN(n2779), 
        .Q(\registers[16][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][12]  ( .D(n1926), .CP(clk), .RN(n2779), 
        .Q(\registers[16][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][11]  ( .D(n1925), .CP(clk), .RN(n2779), 
        .Q(\registers[16][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][10]  ( .D(n1924), .CP(clk), .RN(n2779), 
        .Q(\registers[16][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][9]  ( .D(n1923), .CP(clk), .RN(n2779), 
        .Q(\registers[16][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][8]  ( .D(n1922), .CP(clk), .RN(n2779), 
        .Q(\registers[16][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][7]  ( .D(n1921), .CP(clk), .RN(n2780), 
        .Q(\registers[16][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][6]  ( .D(n1920), .CP(clk), .RN(n2780), 
        .Q(\registers[16][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][5]  ( .D(n1919), .CP(clk), .RN(n2780), 
        .Q(\registers[16][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][4]  ( .D(n1918), .CP(clk), .RN(n2780), 
        .Q(\registers[16][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][3]  ( .D(n1917), .CP(clk), .RN(n2780), 
        .Q(\registers[16][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][2]  ( .D(n1916), .CP(clk), .RN(n2780), 
        .Q(\registers[16][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][1]  ( .D(n1915), .CP(clk), .RN(n2780), 
        .Q(\registers[16][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[16][0]  ( .D(n1914), .CP(clk), .RN(n2780), 
        .Q(\registers[16][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][31]  ( .D(n1849), .CP(clk), .RN(n2780), 
        .Q(\registers[13][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][30]  ( .D(n1848), .CP(clk), .RN(n2780), 
        .Q(\registers[13][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][29]  ( .D(n1847), .CP(clk), .RN(n2780), 
        .Q(\registers[13][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][28]  ( .D(n1846), .CP(clk), .RN(n2780), 
        .Q(\registers[13][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][27]  ( .D(n1845), .CP(clk), .RN(n2781), 
        .Q(\registers[13][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][26]  ( .D(n1844), .CP(clk), .RN(n2781), 
        .Q(\registers[13][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][25]  ( .D(n1843), .CP(clk), .RN(n2781), 
        .Q(\registers[13][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][24]  ( .D(n1842), .CP(clk), .RN(n2781), 
        .Q(\registers[13][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][23]  ( .D(n1841), .CP(clk), .RN(n2781), 
        .Q(\registers[13][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][22]  ( .D(n1840), .CP(clk), .RN(n2781), 
        .Q(\registers[13][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][21]  ( .D(n1839), .CP(clk), .RN(n2781), 
        .Q(\registers[13][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][20]  ( .D(n1838), .CP(clk), .RN(n2781), 
        .Q(\registers[13][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][19]  ( .D(n1837), .CP(clk), .RN(n2781), 
        .Q(\registers[13][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][18]  ( .D(n1836), .CP(clk), .RN(n2781), 
        .Q(\registers[13][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][17]  ( .D(n1835), .CP(clk), .RN(n2781), 
        .Q(\registers[13][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][16]  ( .D(n1834), .CP(clk), .RN(n2781), 
        .Q(\registers[13][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][15]  ( .D(n1833), .CP(clk), .RN(n2782), 
        .Q(\registers[13][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][14]  ( .D(n1832), .CP(clk), .RN(n2782), 
        .Q(\registers[13][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][13]  ( .D(n1831), .CP(clk), .RN(n2782), 
        .Q(\registers[13][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][12]  ( .D(n1830), .CP(clk), .RN(n2782), 
        .Q(\registers[13][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][11]  ( .D(n1829), .CP(clk), .RN(n2782), 
        .Q(\registers[13][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][10]  ( .D(n1828), .CP(clk), .RN(n2782), 
        .Q(\registers[13][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][9]  ( .D(n1827), .CP(clk), .RN(n2782), 
        .Q(\registers[13][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][8]  ( .D(n1826), .CP(clk), .RN(n2782), 
        .Q(\registers[13][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][7]  ( .D(n1825), .CP(clk), .RN(n2782), 
        .Q(\registers[13][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][6]  ( .D(n1824), .CP(clk), .RN(n2782), 
        .Q(\registers[13][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][5]  ( .D(n1823), .CP(clk), .RN(n2782), 
        .Q(\registers[13][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][4]  ( .D(n1822), .CP(clk), .RN(n2782), 
        .Q(\registers[13][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][3]  ( .D(n1821), .CP(clk), .RN(n2769), 
        .Q(\registers[13][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][2]  ( .D(n1820), .CP(clk), .RN(n2765), 
        .Q(\registers[13][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][1]  ( .D(n1819), .CP(clk), .RN(n2765), 
        .Q(\registers[13][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[13][0]  ( .D(n1818), .CP(clk), .RN(n2765), 
        .Q(\registers[13][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][31]  ( .D(n1817), .CP(clk), .RN(n2765), 
        .Q(\registers[12][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][30]  ( .D(n1816), .CP(clk), .RN(n2765), 
        .Q(\registers[12][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][29]  ( .D(n1815), .CP(clk), .RN(n2765), 
        .Q(\registers[12][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][28]  ( .D(n1814), .CP(clk), .RN(n2765), 
        .Q(\registers[12][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][27]  ( .D(n1813), .CP(clk), .RN(n2765), 
        .Q(\registers[12][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][26]  ( .D(n1812), .CP(clk), .RN(n2765), 
        .Q(\registers[12][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][25]  ( .D(n1811), .CP(clk), .RN(n2765), 
        .Q(\registers[12][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][24]  ( .D(n1810), .CP(clk), .RN(n2765), 
        .Q(\registers[12][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][23]  ( .D(n1809), .CP(clk), .RN(n2766), 
        .Q(\registers[12][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][22]  ( .D(n1808), .CP(clk), .RN(n2766), 
        .Q(\registers[12][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][21]  ( .D(n1807), .CP(clk), .RN(n2766), 
        .Q(\registers[12][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][20]  ( .D(n1806), .CP(clk), .RN(n2766), 
        .Q(\registers[12][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][19]  ( .D(n1805), .CP(clk), .RN(n2766), 
        .Q(\registers[12][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][18]  ( .D(n1804), .CP(clk), .RN(n2766), 
        .Q(\registers[12][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][17]  ( .D(n1803), .CP(clk), .RN(n2766), 
        .Q(\registers[12][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][16]  ( .D(n1802), .CP(clk), .RN(n2766), 
        .Q(\registers[12][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][15]  ( .D(n1801), .CP(clk), .RN(n2766), 
        .Q(\registers[12][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][14]  ( .D(n1800), .CP(clk), .RN(n2766), 
        .Q(\registers[12][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][13]  ( .D(n1799), .CP(clk), .RN(n2766), 
        .Q(\registers[12][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][12]  ( .D(n1798), .CP(clk), .RN(n2766), 
        .Q(\registers[12][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][11]  ( .D(n1797), .CP(clk), .RN(n2767), 
        .Q(\registers[12][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][10]  ( .D(n1796), .CP(clk), .RN(n2767), 
        .Q(\registers[12][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][9]  ( .D(n1795), .CP(clk), .RN(n2767), 
        .Q(\registers[12][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][8]  ( .D(n1794), .CP(clk), .RN(n2767), 
        .Q(\registers[12][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][7]  ( .D(n1793), .CP(clk), .RN(n2767), 
        .Q(\registers[12][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][6]  ( .D(n1792), .CP(clk), .RN(n2767), 
        .Q(\registers[12][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][5]  ( .D(n1791), .CP(clk), .RN(n2767), 
        .Q(\registers[12][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][4]  ( .D(n1790), .CP(clk), .RN(n2767), 
        .Q(\registers[12][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][3]  ( .D(n1789), .CP(clk), .RN(n2767), 
        .Q(\registers[12][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][2]  ( .D(n1788), .CP(clk), .RN(n2767), 
        .Q(\registers[12][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][1]  ( .D(n1787), .CP(clk), .RN(n2767), 
        .Q(\registers[12][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[12][0]  ( .D(n1786), .CP(clk), .RN(n2767), 
        .Q(\registers[12][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][31]  ( .D(n1785), .CP(clk), .RN(n2768), 
        .Q(\registers[11][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][30]  ( .D(n1784), .CP(clk), .RN(n2768), 
        .Q(\registers[11][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][29]  ( .D(n1783), .CP(clk), .RN(n2768), 
        .Q(\registers[11][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][28]  ( .D(n1782), .CP(clk), .RN(n2768), 
        .Q(\registers[11][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][27]  ( .D(n1781), .CP(clk), .RN(n2768), 
        .Q(\registers[11][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][26]  ( .D(n1780), .CP(clk), .RN(n2768), 
        .Q(\registers[11][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][25]  ( .D(n1779), .CP(clk), .RN(n2768), 
        .Q(\registers[11][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][24]  ( .D(n1778), .CP(clk), .RN(n2768), 
        .Q(\registers[11][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][23]  ( .D(n1777), .CP(clk), .RN(n2768), 
        .Q(\registers[11][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][22]  ( .D(n1776), .CP(clk), .RN(n2768), 
        .Q(\registers[11][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][21]  ( .D(n1775), .CP(clk), .RN(n2768), 
        .Q(\registers[11][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][20]  ( .D(n1774), .CP(clk), .RN(n2768), 
        .Q(\registers[11][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][19]  ( .D(n1773), .CP(clk), .RN(n2769), 
        .Q(\registers[11][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][18]  ( .D(n1772), .CP(clk), .RN(n2769), 
        .Q(\registers[11][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][17]  ( .D(n1771), .CP(clk), .RN(n2769), 
        .Q(\registers[11][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][16]  ( .D(n1770), .CP(clk), .RN(n2769), 
        .Q(\registers[11][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][15]  ( .D(n1769), .CP(clk), .RN(n2769), 
        .Q(\registers[11][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][14]  ( .D(n1768), .CP(clk), .RN(n2769), 
        .Q(\registers[11][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][13]  ( .D(n1767), .CP(clk), .RN(n2769), 
        .Q(\registers[11][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][12]  ( .D(n1766), .CP(clk), .RN(n2769), 
        .Q(\registers[11][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][11]  ( .D(n1765), .CP(clk), .RN(n2769), 
        .Q(\registers[11][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][10]  ( .D(n1764), .CP(clk), .RN(n2769), 
        .Q(\registers[11][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][9]  ( .D(n1763), .CP(clk), .RN(n2769), 
        .Q(\registers[11][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][8]  ( .D(n1762), .CP(clk), .RN(n2770), 
        .Q(\registers[11][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][7]  ( .D(n1761), .CP(clk), .RN(n2770), 
        .Q(\registers[11][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][6]  ( .D(n1760), .CP(clk), .RN(n2770), 
        .Q(\registers[11][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][5]  ( .D(n1759), .CP(clk), .RN(n2770), 
        .Q(\registers[11][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][4]  ( .D(n1758), .CP(clk), .RN(n2770), 
        .Q(\registers[11][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][3]  ( .D(n1757), .CP(clk), .RN(n2770), 
        .Q(\registers[11][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][2]  ( .D(n1756), .CP(clk), .RN(n2770), 
        .Q(\registers[11][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][1]  ( .D(n1755), .CP(clk), .RN(n2770), 
        .Q(\registers[11][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[11][0]  ( .D(n1754), .CP(clk), .RN(n2770), 
        .Q(\registers[11][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][31]  ( .D(n1753), .CP(clk), .RN(n2770), 
        .Q(\registers[10][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][30]  ( .D(n1752), .CP(clk), .RN(n2770), 
        .Q(\registers[10][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][29]  ( .D(n1751), .CP(clk), .RN(n2770), 
        .Q(\registers[10][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][28]  ( .D(n1750), .CP(clk), .RN(n2771), 
        .Q(\registers[10][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][27]  ( .D(n1749), .CP(clk), .RN(n2771), 
        .Q(\registers[10][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][26]  ( .D(n1748), .CP(clk), .RN(n2771), 
        .Q(\registers[10][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][25]  ( .D(n1747), .CP(clk), .RN(n2771), 
        .Q(\registers[10][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][24]  ( .D(n1746), .CP(clk), .RN(n2771), 
        .Q(\registers[10][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][23]  ( .D(n1745), .CP(clk), .RN(n2771), 
        .Q(\registers[10][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][22]  ( .D(n1744), .CP(clk), .RN(n2771), 
        .Q(\registers[10][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][21]  ( .D(n1743), .CP(clk), .RN(n2771), 
        .Q(\registers[10][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][20]  ( .D(n1742), .CP(clk), .RN(n2771), 
        .Q(\registers[10][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][19]  ( .D(n1741), .CP(clk), .RN(n2771), 
        .Q(\registers[10][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][18]  ( .D(n1740), .CP(clk), .RN(n2771), 
        .Q(\registers[10][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][17]  ( .D(n1739), .CP(clk), .RN(n2771), 
        .Q(\registers[10][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][16]  ( .D(n1738), .CP(clk), .RN(n2772), 
        .Q(\registers[10][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][15]  ( .D(n1737), .CP(clk), .RN(n2772), 
        .Q(\registers[10][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][14]  ( .D(n1736), .CP(clk), .RN(n2772), 
        .Q(\registers[10][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][13]  ( .D(n1735), .CP(clk), .RN(n2772), 
        .Q(\registers[10][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][12]  ( .D(n1734), .CP(clk), .RN(n2772), 
        .Q(\registers[10][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][11]  ( .D(n1733), .CP(clk), .RN(n2772), 
        .Q(\registers[10][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][10]  ( .D(n1732), .CP(clk), .RN(n2772), 
        .Q(\registers[10][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][9]  ( .D(n1731), .CP(clk), .RN(n2772), 
        .Q(\registers[10][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][8]  ( .D(n1730), .CP(clk), .RN(n2772), 
        .Q(\registers[10][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][7]  ( .D(n1729), .CP(clk), .RN(n2772), 
        .Q(\registers[10][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][6]  ( .D(n1728), .CP(clk), .RN(n2772), 
        .Q(\registers[10][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][5]  ( .D(n1727), .CP(clk), .RN(n2772), 
        .Q(\registers[10][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][4]  ( .D(n1726), .CP(clk), .RN(n2773), 
        .Q(\registers[10][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][3]  ( .D(n1725), .CP(clk), .RN(n2773), 
        .Q(\registers[10][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][2]  ( .D(n1724), .CP(clk), .RN(n2773), 
        .Q(\registers[10][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][1]  ( .D(n1723), .CP(clk), .RN(n2773), 
        .Q(\registers[10][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[10][0]  ( .D(n1722), .CP(clk), .RN(n2773), 
        .Q(\registers[10][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][31]  ( .D(n1657), .CP(clk), .RN(n2773), 
        .Q(\registers[7][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][30]  ( .D(n1656), .CP(clk), .RN(n2773), 
        .Q(\registers[7][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][29]  ( .D(n1655), .CP(clk), .RN(n2773), 
        .Q(\registers[7][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][28]  ( .D(n1654), .CP(clk), .RN(n2773), 
        .Q(\registers[7][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][27]  ( .D(n1653), .CP(clk), .RN(n2773), 
        .Q(\registers[7][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][26]  ( .D(n1652), .CP(clk), .RN(n2773), 
        .Q(\registers[7][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][25]  ( .D(n1651), .CP(clk), .RN(n2773), 
        .Q(\registers[7][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][24]  ( .D(n1650), .CP(clk), .RN(n2774), 
        .Q(\registers[7][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][23]  ( .D(n1649), .CP(clk), .RN(n2796), 
        .Q(\registers[7][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][22]  ( .D(n1648), .CP(clk), .RN(n2792), 
        .Q(\registers[7][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][21]  ( .D(n1647), .CP(clk), .RN(n2792), 
        .Q(\registers[7][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][20]  ( .D(n1646), .CP(clk), .RN(n2792), 
        .Q(\registers[7][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][19]  ( .D(n1645), .CP(clk), .RN(n2792), 
        .Q(\registers[7][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][18]  ( .D(n1644), .CP(clk), .RN(n2792), 
        .Q(\registers[7][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][17]  ( .D(n1643), .CP(clk), .RN(n2792), 
        .Q(\registers[7][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][16]  ( .D(n1642), .CP(clk), .RN(n2792), 
        .Q(\registers[7][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][15]  ( .D(n1641), .CP(clk), .RN(n2792), 
        .Q(\registers[7][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][14]  ( .D(n1640), .CP(clk), .RN(n2792), 
        .Q(\registers[7][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][13]  ( .D(n1639), .CP(clk), .RN(n2792), 
        .Q(\registers[7][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][12]  ( .D(n1638), .CP(clk), .RN(n2792), 
        .Q(\registers[7][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][11]  ( .D(n1637), .CP(clk), .RN(n2793), 
        .Q(\registers[7][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][10]  ( .D(n1636), .CP(clk), .RN(n2793), 
        .Q(\registers[7][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][9]  ( .D(n1635), .CP(clk), .RN(n2793), .Q(
        \registers[7][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][8]  ( .D(n1634), .CP(clk), .RN(n2793), .Q(
        \registers[7][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][7]  ( .D(n1633), .CP(clk), .RN(n2793), .Q(
        \registers[7][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][6]  ( .D(n1632), .CP(clk), .RN(n2793), .Q(
        \registers[7][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][5]  ( .D(n1631), .CP(clk), .RN(n2793), .Q(
        \registers[7][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][4]  ( .D(n1630), .CP(clk), .RN(n2793), .Q(
        \registers[7][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][3]  ( .D(n1629), .CP(clk), .RN(n2793), .Q(
        \registers[7][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][2]  ( .D(n1628), .CP(clk), .RN(n2793), .Q(
        \registers[7][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][1]  ( .D(n1627), .CP(clk), .RN(n2793), .Q(
        \registers[7][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[7][0]  ( .D(n1626), .CP(clk), .RN(n2793), .Q(
        \registers[7][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][31]  ( .D(n1625), .CP(clk), .RN(n2794), 
        .Q(\registers[6][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][30]  ( .D(n1624), .CP(clk), .RN(n2794), 
        .Q(\registers[6][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][29]  ( .D(n1623), .CP(clk), .RN(n2794), 
        .Q(\registers[6][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][28]  ( .D(n1622), .CP(clk), .RN(n2794), 
        .Q(\registers[6][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][27]  ( .D(n1621), .CP(clk), .RN(n2794), 
        .Q(\registers[6][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][26]  ( .D(n1620), .CP(clk), .RN(n2794), 
        .Q(\registers[6][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][25]  ( .D(n1619), .CP(clk), .RN(n2794), 
        .Q(\registers[6][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][24]  ( .D(n1618), .CP(clk), .RN(n2794), 
        .Q(\registers[6][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][23]  ( .D(n1617), .CP(clk), .RN(n2794), 
        .Q(\registers[6][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][22]  ( .D(n1616), .CP(clk), .RN(n2794), 
        .Q(\registers[6][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][21]  ( .D(n1615), .CP(clk), .RN(n2794), 
        .Q(\registers[6][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][20]  ( .D(n1614), .CP(clk), .RN(n2794), 
        .Q(\registers[6][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][19]  ( .D(n1613), .CP(clk), .RN(n2795), 
        .Q(\registers[6][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][18]  ( .D(n1612), .CP(clk), .RN(n2795), 
        .Q(\registers[6][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][17]  ( .D(n1611), .CP(clk), .RN(n2795), 
        .Q(\registers[6][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][16]  ( .D(n1610), .CP(clk), .RN(n2795), 
        .Q(\registers[6][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][15]  ( .D(n1609), .CP(clk), .RN(n2795), 
        .Q(\registers[6][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][14]  ( .D(n1608), .CP(clk), .RN(n2795), 
        .Q(\registers[6][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][13]  ( .D(n1607), .CP(clk), .RN(n2795), 
        .Q(\registers[6][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][12]  ( .D(n1606), .CP(clk), .RN(n2795), 
        .Q(\registers[6][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][11]  ( .D(n1605), .CP(clk), .RN(n2795), 
        .Q(\registers[6][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][10]  ( .D(n1604), .CP(clk), .RN(n2795), 
        .Q(\registers[6][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][9]  ( .D(n1603), .CP(clk), .RN(n2795), .Q(
        \registers[6][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][8]  ( .D(n1602), .CP(clk), .RN(n2795), .Q(
        \registers[6][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][7]  ( .D(n1601), .CP(clk), .RN(n2796), .Q(
        \registers[6][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][6]  ( .D(n1600), .CP(clk), .RN(n2796), .Q(
        \registers[6][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][5]  ( .D(n1599), .CP(clk), .RN(n2796), .Q(
        \registers[6][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][4]  ( .D(n1598), .CP(clk), .RN(n2796), .Q(
        \registers[6][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][3]  ( .D(n1597), .CP(clk), .RN(n2796), .Q(
        \registers[6][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][2]  ( .D(n1596), .CP(clk), .RN(n2796), .Q(
        \registers[6][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][1]  ( .D(n1595), .CP(clk), .RN(n2796), .Q(
        \registers[6][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[6][0]  ( .D(n1594), .CP(clk), .RN(n2796), .Q(
        \registers[6][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][31]  ( .D(n1593), .CP(clk), .RN(n2796), 
        .Q(\registers[5][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][30]  ( .D(n1592), .CP(clk), .RN(n2796), 
        .Q(\registers[5][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][29]  ( .D(n1591), .CP(clk), .RN(n2796), 
        .Q(\registers[5][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][28]  ( .D(n1590), .CP(clk), .RN(n2797), 
        .Q(\registers[5][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][27]  ( .D(n1589), .CP(clk), .RN(n2797), 
        .Q(\registers[5][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][26]  ( .D(n1588), .CP(clk), .RN(n2797), 
        .Q(\registers[5][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][25]  ( .D(n1587), .CP(clk), .RN(n2797), 
        .Q(\registers[5][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][24]  ( .D(n1586), .CP(clk), .RN(n2797), 
        .Q(\registers[5][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][23]  ( .D(n1585), .CP(clk), .RN(n2797), 
        .Q(\registers[5][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][22]  ( .D(n1584), .CP(clk), .RN(n2797), 
        .Q(\registers[5][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][21]  ( .D(n1583), .CP(clk), .RN(n2797), 
        .Q(\registers[5][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][20]  ( .D(n1582), .CP(clk), .RN(n2797), 
        .Q(\registers[5][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][19]  ( .D(n1581), .CP(clk), .RN(n2797), 
        .Q(\registers[5][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][18]  ( .D(n1580), .CP(clk), .RN(n2797), 
        .Q(\registers[5][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][17]  ( .D(n1579), .CP(clk), .RN(n2797), 
        .Q(\registers[5][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][16]  ( .D(n1578), .CP(clk), .RN(n2798), 
        .Q(\registers[5][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][15]  ( .D(n1577), .CP(clk), .RN(n2798), 
        .Q(\registers[5][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][14]  ( .D(n1576), .CP(clk), .RN(n2798), 
        .Q(\registers[5][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][13]  ( .D(n1575), .CP(clk), .RN(n2798), 
        .Q(\registers[5][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][12]  ( .D(n1574), .CP(clk), .RN(n2798), 
        .Q(\registers[5][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][11]  ( .D(n1573), .CP(clk), .RN(n2798), 
        .Q(\registers[5][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][10]  ( .D(n1572), .CP(clk), .RN(n2798), 
        .Q(\registers[5][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][9]  ( .D(n1571), .CP(clk), .RN(n2798), .Q(
        \registers[5][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][8]  ( .D(n1570), .CP(clk), .RN(n2798), .Q(
        \registers[5][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][7]  ( .D(n1569), .CP(clk), .RN(n2798), .Q(
        \registers[5][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][6]  ( .D(n1568), .CP(clk), .RN(n2798), .Q(
        \registers[5][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][5]  ( .D(n1567), .CP(clk), .RN(n2798), .Q(
        \registers[5][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][4]  ( .D(n1566), .CP(clk), .RN(n2799), .Q(
        \registers[5][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][3]  ( .D(n1565), .CP(clk), .RN(n2799), .Q(
        \registers[5][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][2]  ( .D(n1564), .CP(clk), .RN(n2799), .Q(
        \registers[5][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][1]  ( .D(n1563), .CP(clk), .RN(n2799), .Q(
        \registers[5][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[5][0]  ( .D(n1562), .CP(clk), .RN(n2799), .Q(
        \registers[5][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][31]  ( .D(n1561), .CP(clk), .RN(n2799), 
        .Q(\registers[4][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][30]  ( .D(n1560), .CP(clk), .RN(n2799), 
        .Q(\registers[4][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][29]  ( .D(n1559), .CP(clk), .RN(n2799), 
        .Q(\registers[4][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][28]  ( .D(n1558), .CP(clk), .RN(n2801), 
        .Q(\registers[4][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][27]  ( .D(n1557), .CP(clk), .RN(n2799), 
        .Q(\registers[4][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][26]  ( .D(n1556), .CP(clk), .RN(n2799), 
        .Q(\registers[4][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][25]  ( .D(n1555), .CP(clk), .RN(n2799), 
        .Q(\registers[4][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][24]  ( .D(n1554), .CP(clk), .RN(n2800), 
        .Q(\registers[4][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][23]  ( .D(n1553), .CP(clk), .RN(n2800), 
        .Q(\registers[4][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][22]  ( .D(n1552), .CP(clk), .RN(n2800), 
        .Q(\registers[4][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][21]  ( .D(n1551), .CP(clk), .RN(n2800), 
        .Q(\registers[4][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][20]  ( .D(n1550), .CP(clk), .RN(n2800), 
        .Q(\registers[4][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][19]  ( .D(n1549), .CP(clk), .RN(n2800), 
        .Q(\registers[4][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][18]  ( .D(n1548), .CP(clk), .RN(n2800), 
        .Q(\registers[4][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][17]  ( .D(n1547), .CP(clk), .RN(n2800), 
        .Q(\registers[4][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][16]  ( .D(n1546), .CP(clk), .RN(n2800), 
        .Q(\registers[4][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][15]  ( .D(n1545), .CP(clk), .RN(n2800), 
        .Q(\registers[4][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][14]  ( .D(n1544), .CP(clk), .RN(n2800), 
        .Q(\registers[4][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][13]  ( .D(n1543), .CP(clk), .RN(n2800), 
        .Q(\registers[4][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][12]  ( .D(n1542), .CP(clk), .RN(n2787), 
        .Q(\registers[4][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][11]  ( .D(n1541), .CP(clk), .RN(n2783), 
        .Q(\registers[4][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][10]  ( .D(n1540), .CP(clk), .RN(n2783), 
        .Q(\registers[4][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][9]  ( .D(n1539), .CP(clk), .RN(n2783), .Q(
        \registers[4][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][8]  ( .D(n1538), .CP(clk), .RN(n2783), .Q(
        \registers[4][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][7]  ( .D(n1537), .CP(clk), .RN(n2783), .Q(
        \registers[4][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][6]  ( .D(n1536), .CP(clk), .RN(n2783), .Q(
        \registers[4][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][5]  ( .D(n1535), .CP(clk), .RN(n2783), .Q(
        \registers[4][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][4]  ( .D(n1534), .CP(clk), .RN(n2783), .Q(
        \registers[4][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][3]  ( .D(n1533), .CP(clk), .RN(n2783), .Q(
        \registers[4][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][2]  ( .D(n1532), .CP(clk), .RN(n2783), .Q(
        \registers[4][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][1]  ( .D(n1531), .CP(clk), .RN(n2783), .Q(
        \registers[4][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[4][0]  ( .D(n1530), .CP(clk), .RN(n2784), .Q(
        \registers[4][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][31]  ( .D(n1529), .CP(clk), .RN(n2784), 
        .Q(\registers[3][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][30]  ( .D(n1528), .CP(clk), .RN(n2784), 
        .Q(\registers[3][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][29]  ( .D(n1527), .CP(clk), .RN(n2784), 
        .Q(\registers[3][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][28]  ( .D(n1526), .CP(clk), .RN(n2784), 
        .Q(\registers[3][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][27]  ( .D(n1525), .CP(clk), .RN(n2784), 
        .Q(\registers[3][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][26]  ( .D(n1524), .CP(clk), .RN(n2784), 
        .Q(\registers[3][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][25]  ( .D(n1523), .CP(clk), .RN(n2784), 
        .Q(\registers[3][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][24]  ( .D(n1522), .CP(clk), .RN(n2784), 
        .Q(\registers[3][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][23]  ( .D(n1521), .CP(clk), .RN(n2784), 
        .Q(\registers[3][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][22]  ( .D(n1520), .CP(clk), .RN(n2784), 
        .Q(\registers[3][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][21]  ( .D(n1519), .CP(clk), .RN(n2784), 
        .Q(\registers[3][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][20]  ( .D(n1518), .CP(clk), .RN(n2785), 
        .Q(\registers[3][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][19]  ( .D(n1517), .CP(clk), .RN(n2785), 
        .Q(\registers[3][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][18]  ( .D(n1516), .CP(clk), .RN(n2785), 
        .Q(\registers[3][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][17]  ( .D(n1515), .CP(clk), .RN(n2785), 
        .Q(\registers[3][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][16]  ( .D(n1514), .CP(clk), .RN(n2785), 
        .Q(\registers[3][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][15]  ( .D(n1513), .CP(clk), .RN(n2785), 
        .Q(\registers[3][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][14]  ( .D(n1512), .CP(clk), .RN(n2785), 
        .Q(\registers[3][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][13]  ( .D(n1511), .CP(clk), .RN(n2785), 
        .Q(\registers[3][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][12]  ( .D(n1510), .CP(clk), .RN(n2785), 
        .Q(\registers[3][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][11]  ( .D(n1509), .CP(clk), .RN(n2785), 
        .Q(\registers[3][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][10]  ( .D(n1508), .CP(clk), .RN(n2785), 
        .Q(\registers[3][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][9]  ( .D(n1507), .CP(clk), .RN(n2785), .Q(
        \registers[3][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][8]  ( .D(n1506), .CP(clk), .RN(n2786), .Q(
        \registers[3][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][7]  ( .D(n1505), .CP(clk), .RN(n2786), .Q(
        \registers[3][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][6]  ( .D(n1504), .CP(clk), .RN(n2786), .Q(
        \registers[3][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][5]  ( .D(n1503), .CP(clk), .RN(n2786), .Q(
        \registers[3][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][4]  ( .D(n1502), .CP(clk), .RN(n2786), .Q(
        \registers[3][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][3]  ( .D(n1501), .CP(clk), .RN(n2786), .Q(
        \registers[3][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][2]  ( .D(n1500), .CP(clk), .RN(n2786), .Q(
        \registers[3][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][1]  ( .D(n1499), .CP(clk), .RN(n2786), .Q(
        \registers[3][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[3][0]  ( .D(n1498), .CP(clk), .RN(n2786), .Q(
        \registers[3][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][31]  ( .D(n1497), .CP(clk), .RN(n2786), 
        .Q(\registers[2][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][30]  ( .D(n1496), .CP(clk), .RN(n2786), 
        .Q(\registers[2][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][29]  ( .D(n1495), .CP(clk), .RN(n2786), 
        .Q(\registers[2][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][28]  ( .D(n1494), .CP(clk), .RN(n2787), 
        .Q(\registers[2][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][27]  ( .D(n1493), .CP(clk), .RN(n2787), 
        .Q(\registers[2][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][26]  ( .D(n1492), .CP(clk), .RN(n2787), 
        .Q(\registers[2][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][25]  ( .D(n1491), .CP(clk), .RN(n2787), 
        .Q(\registers[2][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][24]  ( .D(n1490), .CP(clk), .RN(n2787), 
        .Q(\registers[2][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][23]  ( .D(n1489), .CP(clk), .RN(n2787), 
        .Q(\registers[2][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][22]  ( .D(n1488), .CP(clk), .RN(n2787), 
        .Q(\registers[2][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][21]  ( .D(n1487), .CP(clk), .RN(n2787), 
        .Q(\registers[2][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][20]  ( .D(n1486), .CP(clk), .RN(n2787), 
        .Q(\registers[2][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][19]  ( .D(n1485), .CP(clk), .RN(n2787), 
        .Q(\registers[2][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][18]  ( .D(n1484), .CP(clk), .RN(n2787), 
        .Q(\registers[2][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][17]  ( .D(n1483), .CP(clk), .RN(n2788), 
        .Q(\registers[2][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][16]  ( .D(n1482), .CP(clk), .RN(n2788), 
        .Q(\registers[2][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][15]  ( .D(n1481), .CP(clk), .RN(n2788), 
        .Q(\registers[2][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][14]  ( .D(n1480), .CP(clk), .RN(n2788), 
        .Q(\registers[2][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][13]  ( .D(n1479), .CP(clk), .RN(n2788), 
        .Q(\registers[2][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][12]  ( .D(n1478), .CP(clk), .RN(n2788), 
        .Q(\registers[2][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][11]  ( .D(n1477), .CP(clk), .RN(n2788), 
        .Q(\registers[2][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][10]  ( .D(n1476), .CP(clk), .RN(n2788), 
        .Q(\registers[2][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][9]  ( .D(n1475), .CP(clk), .RN(n2788), .Q(
        \registers[2][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][8]  ( .D(n1474), .CP(clk), .RN(n2788), .Q(
        \registers[2][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][7]  ( .D(n1473), .CP(clk), .RN(n2788), .Q(
        \registers[2][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][6]  ( .D(n1472), .CP(clk), .RN(n2788), .Q(
        \registers[2][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][5]  ( .D(n1471), .CP(clk), .RN(n2789), .Q(
        \registers[2][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][4]  ( .D(n1470), .CP(clk), .RN(n2789), .Q(
        \registers[2][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][3]  ( .D(n1469), .CP(clk), .RN(n2789), .Q(
        \registers[2][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][2]  ( .D(n1468), .CP(clk), .RN(n2789), .Q(
        \registers[2][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][1]  ( .D(n1467), .CP(clk), .RN(n2789), .Q(
        \registers[2][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[2][0]  ( .D(n1466), .CP(clk), .RN(n2789), .Q(
        \registers[2][0] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][31]  ( .D(n1465), .CP(clk), .RN(n2789), 
        .Q(\registers[1][31] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][30]  ( .D(n1464), .CP(clk), .RN(n2789), 
        .Q(\registers[1][30] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][29]  ( .D(n1463), .CP(clk), .RN(n2789), 
        .Q(\registers[1][29] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][28]  ( .D(n1462), .CP(clk), .RN(n2789), 
        .Q(\registers[1][28] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][27]  ( .D(n1461), .CP(clk), .RN(n2789), 
        .Q(\registers[1][27] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][26]  ( .D(n1460), .CP(clk), .RN(n2789), 
        .Q(\registers[1][26] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][25]  ( .D(n1459), .CP(clk), .RN(n2790), 
        .Q(\registers[1][25] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][24]  ( .D(n1458), .CP(clk), .RN(n2790), 
        .Q(\registers[1][24] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][23]  ( .D(n1457), .CP(clk), .RN(n2790), 
        .Q(\registers[1][23] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][22]  ( .D(n1456), .CP(clk), .RN(n2790), 
        .Q(\registers[1][22] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][21]  ( .D(n1455), .CP(clk), .RN(n2790), 
        .Q(\registers[1][21] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][20]  ( .D(n1454), .CP(clk), .RN(n2790), 
        .Q(\registers[1][20] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][19]  ( .D(n1453), .CP(clk), .RN(n2790), 
        .Q(\registers[1][19] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][18]  ( .D(n1452), .CP(clk), .RN(n2790), 
        .Q(\registers[1][18] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][17]  ( .D(n1451), .CP(clk), .RN(n2790), 
        .Q(\registers[1][17] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][16]  ( .D(n1450), .CP(clk), .RN(n2790), 
        .Q(\registers[1][16] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][15]  ( .D(n1449), .CP(clk), .RN(n2790), 
        .Q(\registers[1][15] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][14]  ( .D(n1448), .CP(clk), .RN(n2790), 
        .Q(\registers[1][14] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][13]  ( .D(n1447), .CP(clk), .RN(n2791), 
        .Q(\registers[1][13] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][12]  ( .D(n1446), .CP(clk), .RN(n2791), 
        .Q(\registers[1][12] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][11]  ( .D(n1445), .CP(clk), .RN(n2791), 
        .Q(\registers[1][11] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][10]  ( .D(n1444), .CP(clk), .RN(n2791), 
        .Q(\registers[1][10] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][9]  ( .D(n1443), .CP(clk), .RN(n2791), .Q(
        \registers[1][9] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][8]  ( .D(n1442), .CP(clk), .RN(n2791), .Q(
        \registers[1][8] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][7]  ( .D(n1441), .CP(clk), .RN(n2791), .Q(
        \registers[1][7] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][6]  ( .D(n1440), .CP(clk), .RN(n2791), .Q(
        \registers[1][6] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][5]  ( .D(n1439), .CP(clk), .RN(n2791), .Q(
        \registers[1][5] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][4]  ( .D(n1438), .CP(clk), .RN(n2791), .Q(
        \registers[1][4] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][3]  ( .D(n1437), .CP(clk), .RN(n2791), .Q(
        \registers[1][3] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][2]  ( .D(n1436), .CP(clk), .RN(n2791), .Q(
        \registers[1][2] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][1]  ( .D(n1435), .CP(clk), .RN(n2792), .Q(
        \registers[1][1] ) );
  HS65_LH_DFPRQX9 \registers_reg[1][0]  ( .D(n1434), .CP(clk), .RN(n2799), .Q(
        \registers[1][0] ) );
  HS65_LH_DFPRQNX9 \registers_reg[29][31]  ( .D(n2361), .CP(clk), .RN(n2833), 
        .QN(n1) );
  HS65_LH_DFPRQNX9 \registers_reg[29][30]  ( .D(n2360), .CP(clk), .RN(n2833), 
        .QN(n2) );
  HS65_LH_DFPRQNX9 \registers_reg[29][29]  ( .D(n2359), .CP(clk), .RN(n2833), 
        .QN(n3) );
  HS65_LH_DFPRQNX9 \registers_reg[29][28]  ( .D(n2358), .CP(clk), .RN(n2832), 
        .QN(n4) );
  HS65_LH_DFPRQNX9 \registers_reg[29][27]  ( .D(n2357), .CP(clk), .RN(n2832), 
        .QN(n5) );
  HS65_LH_DFPRQNX9 \registers_reg[29][26]  ( .D(n2356), .CP(clk), .RN(n2832), 
        .QN(n6) );
  HS65_LH_DFPRQNX9 \registers_reg[29][25]  ( .D(n2355), .CP(clk), .RN(n2832), 
        .QN(n7) );
  HS65_LH_DFPRQNX9 \registers_reg[29][24]  ( .D(n2354), .CP(clk), .RN(n2832), 
        .QN(n8) );
  HS65_LH_DFPRQNX9 \registers_reg[29][23]  ( .D(n2353), .CP(clk), .RN(n2832), 
        .QN(n9) );
  HS65_LH_DFPRQNX9 \registers_reg[29][22]  ( .D(n2352), .CP(clk), .RN(n2832), 
        .QN(n10) );
  HS65_LH_DFPRQNX9 \registers_reg[29][21]  ( .D(n2351), .CP(clk), .RN(n2832), 
        .QN(n11) );
  HS65_LH_DFPRQNX9 \registers_reg[29][20]  ( .D(n2350), .CP(clk), .RN(n2832), 
        .QN(n12) );
  HS65_LH_DFPRQNX9 \registers_reg[29][19]  ( .D(n2349), .CP(clk), .RN(n2832), 
        .QN(n13) );
  HS65_LH_DFPRQNX9 \registers_reg[29][18]  ( .D(n2348), .CP(clk), .RN(n2832), 
        .QN(n14) );
  HS65_LH_DFPRQNX9 \registers_reg[29][17]  ( .D(n2347), .CP(clk), .RN(n2832), 
        .QN(n15) );
  HS65_LH_DFPRQNX9 \registers_reg[29][16]  ( .D(n2346), .CP(clk), .RN(n2832), 
        .QN(n16) );
  HS65_LH_DFPRQNX9 \registers_reg[29][15]  ( .D(n2345), .CP(clk), .RN(n2832), 
        .QN(n17) );
  HS65_LH_DFPRQNX9 \registers_reg[29][14]  ( .D(n2344), .CP(clk), .RN(n2831), 
        .QN(n18) );
  HS65_LH_DFPRQNX9 \registers_reg[29][13]  ( .D(n2343), .CP(clk), .RN(n2831), 
        .QN(n19) );
  HS65_LH_DFPRQNX9 \registers_reg[29][12]  ( .D(n2342), .CP(clk), .RN(n2831), 
        .QN(n20) );
  HS65_LH_DFPRQNX9 \registers_reg[29][11]  ( .D(n2341), .CP(clk), .RN(n2831), 
        .QN(n21) );
  HS65_LH_DFPRQNX9 \registers_reg[29][10]  ( .D(n2340), .CP(clk), .RN(n2831), 
        .QN(n22) );
  HS65_LH_DFPRQNX9 \registers_reg[29][9]  ( .D(n2339), .CP(clk), .RN(n2831), 
        .QN(n23) );
  HS65_LH_DFPRQNX9 \registers_reg[29][8]  ( .D(n2338), .CP(clk), .RN(n2831), 
        .QN(n24) );
  HS65_LH_DFPRQNX9 \registers_reg[29][7]  ( .D(n2337), .CP(clk), .RN(n2831), 
        .QN(n25) );
  HS65_LH_DFPRQNX9 \registers_reg[29][6]  ( .D(n2336), .CP(clk), .RN(n2831), 
        .QN(n26) );
  HS65_LH_DFPRQNX9 \registers_reg[29][5]  ( .D(n2335), .CP(clk), .RN(n2831), 
        .QN(n27) );
  HS65_LH_DFPRQNX9 \registers_reg[29][4]  ( .D(n2334), .CP(clk), .RN(n2831), 
        .QN(n28) );
  HS65_LH_DFPRQNX9 \registers_reg[29][3]  ( .D(n2333), .CP(clk), .RN(n2831), 
        .QN(n29) );
  HS65_LH_DFPRQNX9 \registers_reg[29][2]  ( .D(n2332), .CP(clk), .RN(n2831), 
        .QN(n30) );
  HS65_LH_DFPRQNX9 \registers_reg[29][1]  ( .D(n2331), .CP(clk), .RN(n2831), 
        .QN(n31) );
  HS65_LH_DFPRQNX9 \registers_reg[29][0]  ( .D(n2330), .CP(clk), .RN(n2830), 
        .QN(n32) );
  HS65_LH_DFPRQNX9 \registers_reg[27][31]  ( .D(n2297), .CP(clk), .RN(n2826), 
        .QN(n65) );
  HS65_LH_DFPRQNX9 \registers_reg[27][30]  ( .D(n2296), .CP(clk), .RN(n2826), 
        .QN(n66) );
  HS65_LH_DFPRQNX9 \registers_reg[27][29]  ( .D(n2295), .CP(clk), .RN(n2827), 
        .QN(n67) );
  HS65_LH_DFPRQNX9 \registers_reg[27][28]  ( .D(n2294), .CP(clk), .RN(n2827), 
        .QN(n68) );
  HS65_LH_DFPRQNX9 \registers_reg[27][27]  ( .D(n2293), .CP(clk), .RN(n2827), 
        .QN(n69) );
  HS65_LH_DFPRQNX9 \registers_reg[27][26]  ( .D(n2292), .CP(clk), .RN(n2827), 
        .QN(n70) );
  HS65_LH_DFPRQNX9 \registers_reg[27][25]  ( .D(n2291), .CP(clk), .RN(n2827), 
        .QN(n71) );
  HS65_LH_DFPRQNX9 \registers_reg[27][24]  ( .D(n2290), .CP(clk), .RN(n2827), 
        .QN(n72) );
  HS65_LH_DFPRQNX9 \registers_reg[27][23]  ( .D(n2289), .CP(clk), .RN(n2827), 
        .QN(n73) );
  HS65_LH_DFPRQNX9 \registers_reg[27][22]  ( .D(n2288), .CP(clk), .RN(n2827), 
        .QN(n74) );
  HS65_LH_DFPRQNX9 \registers_reg[27][21]  ( .D(n2287), .CP(clk), .RN(n2827), 
        .QN(n75) );
  HS65_LH_DFPRQNX9 \registers_reg[27][20]  ( .D(n2286), .CP(clk), .RN(n2827), 
        .QN(n76) );
  HS65_LH_DFPRQNX9 \registers_reg[27][19]  ( .D(n2285), .CP(clk), .RN(n2827), 
        .QN(n77) );
  HS65_LH_DFPRQNX9 \registers_reg[27][18]  ( .D(n2284), .CP(clk), .RN(n2827), 
        .QN(n78) );
  HS65_LH_DFPRQNX9 \registers_reg[27][17]  ( .D(n2283), .CP(clk), .RN(n2827), 
        .QN(n79) );
  HS65_LH_DFPRQNX9 \registers_reg[27][16]  ( .D(n2282), .CP(clk), .RN(n2828), 
        .QN(n80) );
  HS65_LH_DFPRQNX9 \registers_reg[27][15]  ( .D(n2281), .CP(clk), .RN(n2828), 
        .QN(n81) );
  HS65_LH_DFPRQNX9 \registers_reg[27][14]  ( .D(n2280), .CP(clk), .RN(n2828), 
        .QN(n82) );
  HS65_LH_DFPRQNX9 \registers_reg[27][13]  ( .D(n2279), .CP(clk), .RN(n2828), 
        .QN(n83) );
  HS65_LH_DFPRQNX9 \registers_reg[27][12]  ( .D(n2278), .CP(clk), .RN(n2828), 
        .QN(n84) );
  HS65_LH_DFPRQNX9 \registers_reg[27][11]  ( .D(n2277), .CP(clk), .RN(n2828), 
        .QN(n85) );
  HS65_LH_DFPRQNX9 \registers_reg[27][10]  ( .D(n2276), .CP(clk), .RN(n2828), 
        .QN(n86) );
  HS65_LH_DFPRQNX9 \registers_reg[27][9]  ( .D(n2275), .CP(clk), .RN(n2828), 
        .QN(n87) );
  HS65_LH_DFPRQNX9 \registers_reg[27][8]  ( .D(n2274), .CP(clk), .RN(n2828), 
        .QN(n88) );
  HS65_LH_DFPRQNX9 \registers_reg[27][7]  ( .D(n2273), .CP(clk), .RN(n2828), 
        .QN(n89) );
  HS65_LH_DFPRQNX9 \registers_reg[27][6]  ( .D(n2272), .CP(clk), .RN(n2828), 
        .QN(n90) );
  HS65_LH_DFPRQNX9 \registers_reg[27][5]  ( .D(n2271), .CP(clk), .RN(n2828), 
        .QN(n91) );
  HS65_LH_DFPRQNX9 \registers_reg[27][4]  ( .D(n2270), .CP(clk), .RN(n2828), 
        .QN(n92) );
  HS65_LH_DFPRQNX9 \registers_reg[27][3]  ( .D(n2269), .CP(clk), .RN(n2828), 
        .QN(n93) );
  HS65_LH_DFPRQNX9 \registers_reg[27][2]  ( .D(n2268), .CP(clk), .RN(n2829), 
        .QN(n94) );
  HS65_LH_DFPRQNX9 \registers_reg[27][1]  ( .D(n2267), .CP(clk), .RN(n2829), 
        .QN(n95) );
  HS65_LH_DFPRQNX9 \registers_reg[27][0]  ( .D(n2266), .CP(clk), .RN(n2829), 
        .QN(n96) );
  HS65_LH_DFPRQNX9 \registers_reg[15][31]  ( .D(n1913), .CP(clk), .RN(n2842), 
        .QN(n129) );
  HS65_LH_DFPRQNX9 \registers_reg[15][30]  ( .D(n1912), .CP(clk), .RN(n2842), 
        .QN(n130) );
  HS65_LH_DFPRQNX9 \registers_reg[15][29]  ( .D(n1911), .CP(clk), .RN(n2842), 
        .QN(n131) );
  HS65_LH_DFPRQNX9 \registers_reg[15][28]  ( .D(n1910), .CP(clk), .RN(n2842), 
        .QN(n132) );
  HS65_LH_DFPRQNX9 \registers_reg[15][27]  ( .D(n1909), .CP(clk), .RN(n2841), 
        .QN(n133) );
  HS65_LH_DFPRQNX9 \registers_reg[15][26]  ( .D(n1908), .CP(clk), .RN(n2841), 
        .QN(n134) );
  HS65_LH_DFPRQNX9 \registers_reg[15][25]  ( .D(n1907), .CP(clk), .RN(n2841), 
        .QN(n135) );
  HS65_LH_DFPRQNX9 \registers_reg[15][24]  ( .D(n1906), .CP(clk), .RN(n2841), 
        .QN(n136) );
  HS65_LH_DFPRQNX9 \registers_reg[15][23]  ( .D(n1905), .CP(clk), .RN(n2841), 
        .QN(n137) );
  HS65_LH_DFPRQNX9 \registers_reg[15][22]  ( .D(n1904), .CP(clk), .RN(n2841), 
        .QN(n138) );
  HS65_LH_DFPRQNX9 \registers_reg[15][21]  ( .D(n1903), .CP(clk), .RN(n2841), 
        .QN(n139) );
  HS65_LH_DFPRQNX9 \registers_reg[15][20]  ( .D(n1902), .CP(clk), .RN(n2841), 
        .QN(n140) );
  HS65_LH_DFPRQNX9 \registers_reg[15][19]  ( .D(n1901), .CP(clk), .RN(n2841), 
        .QN(n141) );
  HS65_LH_DFPRQNX9 \registers_reg[15][18]  ( .D(n1900), .CP(clk), .RN(n2841), 
        .QN(n142) );
  HS65_LH_DFPRQNX9 \registers_reg[15][17]  ( .D(n1899), .CP(clk), .RN(n2841), 
        .QN(n143) );
  HS65_LH_DFPRQNX9 \registers_reg[15][16]  ( .D(n1898), .CP(clk), .RN(n2841), 
        .QN(n144) );
  HS65_LH_DFPRQNX9 \registers_reg[15][15]  ( .D(n1897), .CP(clk), .RN(n2841), 
        .QN(n145) );
  HS65_LH_DFPRQNX9 \registers_reg[15][14]  ( .D(n1896), .CP(clk), .RN(n2836), 
        .QN(n146) );
  HS65_LH_DFPRQNX9 \registers_reg[15][13]  ( .D(n1895), .CP(clk), .RN(n2836), 
        .QN(n147) );
  HS65_LH_DFPRQNX9 \registers_reg[15][12]  ( .D(n1894), .CP(clk), .RN(n2836), 
        .QN(n148) );
  HS65_LH_DFPRQNX9 \registers_reg[15][11]  ( .D(n1893), .CP(clk), .RN(n2836), 
        .QN(n149) );
  HS65_LH_DFPRQNX9 \registers_reg[15][10]  ( .D(n1892), .CP(clk), .RN(n2836), 
        .QN(n150) );
  HS65_LH_DFPRQNX9 \registers_reg[15][9]  ( .D(n1891), .CP(clk), .RN(n2836), 
        .QN(n151) );
  HS65_LH_DFPRQNX9 \registers_reg[15][8]  ( .D(n1890), .CP(clk), .RN(n2836), 
        .QN(n152) );
  HS65_LH_DFPRQNX9 \registers_reg[15][7]  ( .D(n1889), .CP(clk), .RN(n2835), 
        .QN(n153) );
  HS65_LH_DFPRQNX9 \registers_reg[15][6]  ( .D(n1888), .CP(clk), .RN(n2835), 
        .QN(n154) );
  HS65_LH_DFPRQNX9 \registers_reg[15][5]  ( .D(n1887), .CP(clk), .RN(n2835), 
        .QN(n155) );
  HS65_LH_DFPRQNX9 \registers_reg[15][4]  ( .D(n1886), .CP(clk), .RN(n2835), 
        .QN(n156) );
  HS65_LH_DFPRQNX9 \registers_reg[15][3]  ( .D(n1885), .CP(clk), .RN(n2835), 
        .QN(n157) );
  HS65_LH_DFPRQNX9 \registers_reg[15][2]  ( .D(n1884), .CP(clk), .RN(n2835), 
        .QN(n158) );
  HS65_LH_DFPRQNX9 \registers_reg[15][1]  ( .D(n1883), .CP(clk), .RN(n2835), 
        .QN(n159) );
  HS65_LH_DFPRQNX9 \registers_reg[15][0]  ( .D(n1882), .CP(clk), .RN(n2835), 
        .QN(n160) );
  HS65_LH_DFPRQNX9 \registers_reg[9][31]  ( .D(n1721), .CP(clk), .RN(n2836), 
        .QN(n193) );
  HS65_LH_DFPRQNX9 \registers_reg[9][30]  ( .D(n1720), .CP(clk), .RN(n2836), 
        .QN(n194) );
  HS65_LH_DFPRQNX9 \registers_reg[9][29]  ( .D(n1719), .CP(clk), .RN(n2836), 
        .QN(n195) );
  HS65_LH_DFPRQNX9 \registers_reg[9][28]  ( .D(n1718), .CP(clk), .RN(n2836), 
        .QN(n196) );
  HS65_LH_DFPRQNX9 \registers_reg[9][27]  ( .D(n1717), .CP(clk), .RN(n2836), 
        .QN(n197) );
  HS65_LH_DFPRQNX9 \registers_reg[9][26]  ( .D(n1716), .CP(clk), .RN(n2836), 
        .QN(n198) );
  HS65_LH_DFPRQNX9 \registers_reg[9][25]  ( .D(n1715), .CP(clk), .RN(n2833), 
        .QN(n199) );
  HS65_LH_DFPRQNX9 \registers_reg[9][24]  ( .D(n1714), .CP(clk), .RN(n2836), 
        .QN(n200) );
  HS65_LH_DFPRQNX9 \registers_reg[9][23]  ( .D(n1713), .CP(clk), .RN(n2837), 
        .QN(n201) );
  HS65_LH_DFPRQNX9 \registers_reg[9][22]  ( .D(n1712), .CP(clk), .RN(n2837), 
        .QN(n202) );
  HS65_LH_DFPRQNX9 \registers_reg[9][21]  ( .D(n1711), .CP(clk), .RN(n2837), 
        .QN(n203) );
  HS65_LH_DFPRQNX9 \registers_reg[9][20]  ( .D(n1710), .CP(clk), .RN(n2837), 
        .QN(n204) );
  HS65_LH_DFPRQNX9 \registers_reg[9][19]  ( .D(n1709), .CP(clk), .RN(n2837), 
        .QN(n205) );
  HS65_LH_DFPRQNX9 \registers_reg[9][18]  ( .D(n1708), .CP(clk), .RN(n2837), 
        .QN(n206) );
  HS65_LH_DFPRQNX9 \registers_reg[9][17]  ( .D(n1707), .CP(clk), .RN(n2837), 
        .QN(n207) );
  HS65_LH_DFPRQNX9 \registers_reg[9][16]  ( .D(n1706), .CP(clk), .RN(n2837), 
        .QN(n208) );
  HS65_LH_DFPRQNX9 \registers_reg[9][15]  ( .D(n1705), .CP(clk), .RN(n2837), 
        .QN(n209) );
  HS65_LH_DFPRQNX9 \registers_reg[9][14]  ( .D(n1704), .CP(clk), .RN(n2837), 
        .QN(n210) );
  HS65_LH_DFPRQNX9 \registers_reg[9][13]  ( .D(n1703), .CP(clk), .RN(n2837), 
        .QN(n211) );
  HS65_LH_DFPRQNX9 \registers_reg[9][12]  ( .D(n1702), .CP(clk), .RN(n2837), 
        .QN(n212) );
  HS65_LH_DFPRQNX9 \registers_reg[9][11]  ( .D(n1701), .CP(clk), .RN(n2837), 
        .QN(n213) );
  HS65_LH_DFPRQNX9 \registers_reg[9][10]  ( .D(n1700), .CP(clk), .RN(n2837), 
        .QN(n214) );
  HS65_LH_DFPRQNX9 \registers_reg[9][9]  ( .D(n1699), .CP(clk), .RN(n2838), 
        .QN(n215) );
  HS65_LH_DFPRQNX9 \registers_reg[9][8]  ( .D(n1698), .CP(clk), .RN(n2838), 
        .QN(n216) );
  HS65_LH_DFPRQNX9 \registers_reg[9][7]  ( .D(n1697), .CP(clk), .RN(n2838), 
        .QN(n217) );
  HS65_LH_DFPRQNX9 \registers_reg[9][6]  ( .D(n1696), .CP(clk), .RN(n2838), 
        .QN(n218) );
  HS65_LH_DFPRQNX9 \registers_reg[9][5]  ( .D(n1695), .CP(clk), .RN(n2838), 
        .QN(n219) );
  HS65_LH_DFPRQNX9 \registers_reg[9][4]  ( .D(n1694), .CP(clk), .RN(n2838), 
        .QN(n220) );
  HS65_LH_DFPRQNX9 \registers_reg[9][3]  ( .D(n1693), .CP(clk), .RN(n2838), 
        .QN(n221) );
  HS65_LH_DFPRQNX9 \registers_reg[9][2]  ( .D(n1692), .CP(clk), .RN(n2838), 
        .QN(n222) );
  HS65_LH_DFPRQNX9 \registers_reg[9][1]  ( .D(n1691), .CP(clk), .RN(n2838), 
        .QN(n223) );
  HS65_LH_DFPRQNX9 \registers_reg[9][0]  ( .D(n1690), .CP(clk), .RN(n2838), 
        .QN(n224) );
  HS65_LH_DFPRQNX9 \registers_reg[28][31]  ( .D(n2329), .CP(clk), .RN(n2830), 
        .QN(n33) );
  HS65_LH_DFPRQNX9 \registers_reg[28][30]  ( .D(n2328), .CP(clk), .RN(n2830), 
        .QN(n34) );
  HS65_LH_DFPRQNX9 \registers_reg[28][29]  ( .D(n2327), .CP(clk), .RN(n2830), 
        .QN(n35) );
  HS65_LH_DFPRQNX9 \registers_reg[28][28]  ( .D(n2326), .CP(clk), .RN(n2830), 
        .QN(n36) );
  HS65_LH_DFPRQNX9 \registers_reg[28][27]  ( .D(n2325), .CP(clk), .RN(n2830), 
        .QN(n37) );
  HS65_LH_DFPRQNX9 \registers_reg[28][26]  ( .D(n2324), .CP(clk), .RN(n2830), 
        .QN(n38) );
  HS65_LH_DFPRQNX9 \registers_reg[28][25]  ( .D(n2323), .CP(clk), .RN(n2830), 
        .QN(n39) );
  HS65_LH_DFPRQNX9 \registers_reg[28][24]  ( .D(n2322), .CP(clk), .RN(n2830), 
        .QN(n40) );
  HS65_LH_DFPRQNX9 \registers_reg[28][23]  ( .D(n2321), .CP(clk), .RN(n2830), 
        .QN(n41) );
  HS65_LH_DFPRQNX9 \registers_reg[28][22]  ( .D(n2320), .CP(clk), .RN(n2830), 
        .QN(n42) );
  HS65_LH_DFPRQNX9 \registers_reg[28][21]  ( .D(n2319), .CP(clk), .RN(n2830), 
        .QN(n43) );
  HS65_LH_DFPRQNX9 \registers_reg[28][20]  ( .D(n2318), .CP(clk), .RN(n2830), 
        .QN(n44) );
  HS65_LH_DFPRQNX9 \registers_reg[28][19]  ( .D(n2317), .CP(clk), .RN(n2830), 
        .QN(n45) );
  HS65_LH_DFPRQNX9 \registers_reg[28][18]  ( .D(n2316), .CP(clk), .RN(n2829), 
        .QN(n46) );
  HS65_LH_DFPRQNX9 \registers_reg[28][17]  ( .D(n2315), .CP(clk), .RN(n2829), 
        .QN(n47) );
  HS65_LH_DFPRQNX9 \registers_reg[28][16]  ( .D(n2314), .CP(clk), .RN(n2829), 
        .QN(n48) );
  HS65_LH_DFPRQNX9 \registers_reg[28][15]  ( .D(n2313), .CP(clk), .RN(n2829), 
        .QN(n49) );
  HS65_LH_DFPRQNX9 \registers_reg[28][14]  ( .D(n2312), .CP(clk), .RN(n2829), 
        .QN(n50) );
  HS65_LH_DFPRQNX9 \registers_reg[28][13]  ( .D(n2311), .CP(clk), .RN(n2829), 
        .QN(n51) );
  HS65_LH_DFPRQNX9 \registers_reg[28][12]  ( .D(n2310), .CP(clk), .RN(n2829), 
        .QN(n52) );
  HS65_LH_DFPRQNX9 \registers_reg[28][11]  ( .D(n2309), .CP(clk), .RN(n2829), 
        .QN(n53) );
  HS65_LH_DFPRQNX9 \registers_reg[28][10]  ( .D(n2308), .CP(clk), .RN(n2829), 
        .QN(n54) );
  HS65_LH_DFPRQNX9 \registers_reg[28][9]  ( .D(n2307), .CP(clk), .RN(n2829), 
        .QN(n55) );
  HS65_LH_DFPRQNX9 \registers_reg[28][8]  ( .D(n2306), .CP(clk), .RN(n2829), 
        .QN(n56) );
  HS65_LH_DFPRQNX9 \registers_reg[28][7]  ( .D(n2305), .CP(clk), .RN(n2827), 
        .QN(n57) );
  HS65_LH_DFPRQNX9 \registers_reg[28][6]  ( .D(n2304), .CP(clk), .RN(n2826), 
        .QN(n58) );
  HS65_LH_DFPRQNX9 \registers_reg[28][5]  ( .D(n2303), .CP(clk), .RN(n2826), 
        .QN(n59) );
  HS65_LH_DFPRQNX9 \registers_reg[28][4]  ( .D(n2302), .CP(clk), .RN(n2826), 
        .QN(n60) );
  HS65_LH_DFPRQNX9 \registers_reg[28][3]  ( .D(n2301), .CP(clk), .RN(n2826), 
        .QN(n61) );
  HS65_LH_DFPRQNX9 \registers_reg[28][2]  ( .D(n2300), .CP(clk), .RN(n2826), 
        .QN(n62) );
  HS65_LH_DFPRQNX9 \registers_reg[28][1]  ( .D(n2299), .CP(clk), .RN(n2826), 
        .QN(n63) );
  HS65_LH_DFPRQNX9 \registers_reg[28][0]  ( .D(n2298), .CP(clk), .RN(n2826), 
        .QN(n64) );
  HS65_LH_DFPRQNX9 \registers_reg[26][31]  ( .D(n2265), .CP(clk), .RN(n2844), 
        .QN(n97) );
  HS65_LH_DFPRQNX9 \registers_reg[26][30]  ( .D(n2264), .CP(clk), .RN(n2844), 
        .QN(n98) );
  HS65_LH_DFPRQNX9 \registers_reg[26][29]  ( .D(n2263), .CP(clk), .RN(n2844), 
        .QN(n99) );
  HS65_LH_DFPRQNX9 \registers_reg[26][28]  ( .D(n2262), .CP(clk), .RN(n2844), 
        .QN(n100) );
  HS65_LH_DFPRQNX9 \registers_reg[26][27]  ( .D(n2261), .CP(clk), .RN(n2844), 
        .QN(n101) );
  HS65_LH_DFPRQNX9 \registers_reg[26][26]  ( .D(n2260), .CP(clk), .RN(n2844), 
        .QN(n102) );
  HS65_LH_DFPRQNX9 \registers_reg[26][25]  ( .D(n2259), .CP(clk), .RN(n2844), 
        .QN(n103) );
  HS65_LH_DFPRQNX9 \registers_reg[26][24]  ( .D(n2258), .CP(clk), .RN(n2844), 
        .QN(n104) );
  HS65_LH_DFPRQNX9 \registers_reg[26][23]  ( .D(n2257), .CP(clk), .RN(n2843), 
        .QN(n105) );
  HS65_LH_DFPRQNX9 \registers_reg[26][22]  ( .D(n2256), .CP(clk), .RN(n2843), 
        .QN(n106) );
  HS65_LH_DFPRQNX9 \registers_reg[26][21]  ( .D(n2255), .CP(clk), .RN(n2843), 
        .QN(n107) );
  HS65_LH_DFPRQNX9 \registers_reg[26][20]  ( .D(n2254), .CP(clk), .RN(n2843), 
        .QN(n108) );
  HS65_LH_DFPRQNX9 \registers_reg[26][19]  ( .D(n2253), .CP(clk), .RN(n2843), 
        .QN(n109) );
  HS65_LH_DFPRQNX9 \registers_reg[26][18]  ( .D(n2252), .CP(clk), .RN(n2843), 
        .QN(n110) );
  HS65_LH_DFPRQNX9 \registers_reg[26][17]  ( .D(n2251), .CP(clk), .RN(n2843), 
        .QN(n111) );
  HS65_LH_DFPRQNX9 \registers_reg[26][16]  ( .D(n2250), .CP(clk), .RN(n2843), 
        .QN(n112) );
  HS65_LH_DFPRQNX9 \registers_reg[26][15]  ( .D(n2249), .CP(clk), .RN(n2843), 
        .QN(n113) );
  HS65_LH_DFPRQNX9 \registers_reg[26][14]  ( .D(n2248), .CP(clk), .RN(n2843), 
        .QN(n114) );
  HS65_LH_DFPRQNX9 \registers_reg[26][13]  ( .D(n2247), .CP(clk), .RN(n2843), 
        .QN(n115) );
  HS65_LH_DFPRQNX9 \registers_reg[26][12]  ( .D(n2246), .CP(clk), .RN(n2843), 
        .QN(n116) );
  HS65_LH_DFPRQNX9 \registers_reg[26][11]  ( .D(n2245), .CP(clk), .RN(n2843), 
        .QN(n117) );
  HS65_LH_DFPRQNX9 \registers_reg[26][10]  ( .D(n2244), .CP(clk), .RN(n2843), 
        .QN(n118) );
  HS65_LH_DFPRQNX9 \registers_reg[26][9]  ( .D(n2243), .CP(clk), .RN(n2842), 
        .QN(n119) );
  HS65_LH_DFPRQNX9 \registers_reg[26][8]  ( .D(n2242), .CP(clk), .RN(n2842), 
        .QN(n120) );
  HS65_LH_DFPRQNX9 \registers_reg[26][7]  ( .D(n2241), .CP(clk), .RN(n2842), 
        .QN(n121) );
  HS65_LH_DFPRQNX9 \registers_reg[26][6]  ( .D(n2240), .CP(clk), .RN(n2842), 
        .QN(n122) );
  HS65_LH_DFPRQNX9 \registers_reg[26][5]  ( .D(n2239), .CP(clk), .RN(n2842), 
        .QN(n123) );
  HS65_LH_DFPRQNX9 \registers_reg[26][4]  ( .D(n2238), .CP(clk), .RN(n2842), 
        .QN(n124) );
  HS65_LH_DFPRQNX9 \registers_reg[26][3]  ( .D(n2237), .CP(clk), .RN(n2842), 
        .QN(n125) );
  HS65_LH_DFPRQNX9 \registers_reg[26][2]  ( .D(n2236), .CP(clk), .RN(n2842), 
        .QN(n126) );
  HS65_LH_DFPRQNX9 \registers_reg[26][1]  ( .D(n2235), .CP(clk), .RN(n2842), 
        .QN(n127) );
  HS65_LH_DFPRQNX9 \registers_reg[26][0]  ( .D(n2234), .CP(clk), .RN(n2842), 
        .QN(n128) );
  HS65_LH_DFPRQNX9 \registers_reg[14][31]  ( .D(n1881), .CP(clk), .RN(n2835), 
        .QN(n161) );
  HS65_LH_DFPRQNX9 \registers_reg[14][30]  ( .D(n1880), .CP(clk), .RN(n2835), 
        .QN(n162) );
  HS65_LH_DFPRQNX9 \registers_reg[14][29]  ( .D(n1879), .CP(clk), .RN(n2835), 
        .QN(n163) );
  HS65_LH_DFPRQNX9 \registers_reg[14][28]  ( .D(n1878), .CP(clk), .RN(n2835), 
        .QN(n164) );
  HS65_LH_DFPRQNX9 \registers_reg[14][27]  ( .D(n1877), .CP(clk), .RN(n2835), 
        .QN(n165) );
  HS65_LH_DFPRQNX9 \registers_reg[14][26]  ( .D(n1876), .CP(clk), .RN(n2835), 
        .QN(n166) );
  HS65_LH_DFPRQNX9 \registers_reg[14][25]  ( .D(n1875), .CP(clk), .RN(n2834), 
        .QN(n167) );
  HS65_LH_DFPRQNX9 \registers_reg[14][24]  ( .D(n1874), .CP(clk), .RN(n2834), 
        .QN(n168) );
  HS65_LH_DFPRQNX9 \registers_reg[14][23]  ( .D(n1873), .CP(clk), .RN(n2834), 
        .QN(n169) );
  HS65_LH_DFPRQNX9 \registers_reg[14][22]  ( .D(n1872), .CP(clk), .RN(n2834), 
        .QN(n170) );
  HS65_LH_DFPRQNX9 \registers_reg[14][21]  ( .D(n1871), .CP(clk), .RN(n2834), 
        .QN(n171) );
  HS65_LH_DFPRQNX9 \registers_reg[14][20]  ( .D(n1870), .CP(clk), .RN(n2834), 
        .QN(n172) );
  HS65_LH_DFPRQNX9 \registers_reg[14][19]  ( .D(n1869), .CP(clk), .RN(n2834), 
        .QN(n173) );
  HS65_LH_DFPRQNX9 \registers_reg[14][18]  ( .D(n1868), .CP(clk), .RN(n2834), 
        .QN(n174) );
  HS65_LH_DFPRQNX9 \registers_reg[14][17]  ( .D(n1867), .CP(clk), .RN(n2834), 
        .QN(n175) );
  HS65_LH_DFPRQNX9 \registers_reg[14][16]  ( .D(n1866), .CP(clk), .RN(n2834), 
        .QN(n176) );
  HS65_LH_DFPRQNX9 \registers_reg[14][15]  ( .D(n1865), .CP(clk), .RN(n2834), 
        .QN(n177) );
  HS65_LH_DFPRQNX9 \registers_reg[14][14]  ( .D(n1864), .CP(clk), .RN(n2834), 
        .QN(n178) );
  HS65_LH_DFPRQNX9 \registers_reg[14][13]  ( .D(n1863), .CP(clk), .RN(n2834), 
        .QN(n179) );
  HS65_LH_DFPRQNX9 \registers_reg[14][12]  ( .D(n1862), .CP(clk), .RN(n2834), 
        .QN(n180) );
  HS65_LH_DFPRQNX9 \registers_reg[14][11]  ( .D(n1861), .CP(clk), .RN(n2833), 
        .QN(n181) );
  HS65_LH_DFPRQNX9 \registers_reg[14][10]  ( .D(n1860), .CP(clk), .RN(n2833), 
        .QN(n182) );
  HS65_LH_DFPRQNX9 \registers_reg[14][9]  ( .D(n1859), .CP(clk), .RN(n2833), 
        .QN(n183) );
  HS65_LH_DFPRQNX9 \registers_reg[14][8]  ( .D(n1858), .CP(clk), .RN(n2833), 
        .QN(n184) );
  HS65_LH_DFPRQNX9 \registers_reg[14][7]  ( .D(n1857), .CP(clk), .RN(n2833), 
        .QN(n185) );
  HS65_LH_DFPRQNX9 \registers_reg[14][6]  ( .D(n1856), .CP(clk), .RN(n2833), 
        .QN(n186) );
  HS65_LH_DFPRQNX9 \registers_reg[14][5]  ( .D(n1855), .CP(clk), .RN(n2833), 
        .QN(n187) );
  HS65_LH_DFPRQNX9 \registers_reg[14][4]  ( .D(n1854), .CP(clk), .RN(n2833), 
        .QN(n188) );
  HS65_LH_DFPRQNX9 \registers_reg[14][3]  ( .D(n1853), .CP(clk), .RN(n2833), 
        .QN(n189) );
  HS65_LH_DFPRQNX9 \registers_reg[14][2]  ( .D(n1852), .CP(clk), .RN(n2833), 
        .QN(n190) );
  HS65_LH_DFPRQNX9 \registers_reg[14][1]  ( .D(n1851), .CP(clk), .RN(n2838), 
        .QN(n191) );
  HS65_LH_DFPRQNX9 \registers_reg[14][0]  ( .D(n1850), .CP(clk), .RN(n2826), 
        .QN(n192) );
  HS65_LH_DFPRQNX9 \registers_reg[8][31]  ( .D(n1689), .CP(clk), .RN(n2838), 
        .QN(n225) );
  HS65_LH_DFPRQNX9 \registers_reg[8][30]  ( .D(n1688), .CP(clk), .RN(n2838), 
        .QN(n226) );
  HS65_LH_DFPRQNX9 \registers_reg[8][29]  ( .D(n1687), .CP(clk), .RN(n2838), 
        .QN(n227) );
  HS65_LH_DFPRQNX9 \registers_reg[8][28]  ( .D(n1686), .CP(clk), .RN(n2839), 
        .QN(n228) );
  HS65_LH_DFPRQNX9 \registers_reg[8][27]  ( .D(n1685), .CP(clk), .RN(n2839), 
        .QN(n229) );
  HS65_LH_DFPRQNX9 \registers_reg[8][26]  ( .D(n1684), .CP(clk), .RN(n2839), 
        .QN(n230) );
  HS65_LH_DFPRQNX9 \registers_reg[8][25]  ( .D(n1683), .CP(clk), .RN(n2839), 
        .QN(n231) );
  HS65_LH_DFPRQNX9 \registers_reg[8][24]  ( .D(n1682), .CP(clk), .RN(n2839), 
        .QN(n232) );
  HS65_LH_DFPRQNX9 \registers_reg[8][23]  ( .D(n1681), .CP(clk), .RN(n2839), 
        .QN(n233) );
  HS65_LH_DFPRQNX9 \registers_reg[8][22]  ( .D(n1680), .CP(clk), .RN(n2839), 
        .QN(n234) );
  HS65_LH_DFPRQNX9 \registers_reg[8][21]  ( .D(n1679), .CP(clk), .RN(n2839), 
        .QN(n235) );
  HS65_LH_DFPRQNX9 \registers_reg[8][20]  ( .D(n1678), .CP(clk), .RN(n2839), 
        .QN(n236) );
  HS65_LH_DFPRQNX9 \registers_reg[8][19]  ( .D(n1677), .CP(clk), .RN(n2839), 
        .QN(n237) );
  HS65_LH_DFPRQNX9 \registers_reg[8][18]  ( .D(n1676), .CP(clk), .RN(n2839), 
        .QN(n238) );
  HS65_LH_DFPRQNX9 \registers_reg[8][17]  ( .D(n1675), .CP(clk), .RN(n2839), 
        .QN(n239) );
  HS65_LH_DFPRQNX9 \registers_reg[8][16]  ( .D(n1674), .CP(clk), .RN(n2839), 
        .QN(n240) );
  HS65_LH_DFPRQNX9 \registers_reg[8][15]  ( .D(n1673), .CP(clk), .RN(n2839), 
        .QN(n241) );
  HS65_LH_DFPRQNX9 \registers_reg[8][14]  ( .D(n1672), .CP(clk), .RN(n2840), 
        .QN(n242) );
  HS65_LH_DFPRQNX9 \registers_reg[8][13]  ( .D(n1671), .CP(clk), .RN(n2840), 
        .QN(n243) );
  HS65_LH_DFPRQNX9 \registers_reg[8][12]  ( .D(n1670), .CP(clk), .RN(n2840), 
        .QN(n244) );
  HS65_LH_DFPRQNX9 \registers_reg[8][11]  ( .D(n1669), .CP(clk), .RN(n2840), 
        .QN(n245) );
  HS65_LH_DFPRQNX9 \registers_reg[8][10]  ( .D(n1668), .CP(clk), .RN(n2840), 
        .QN(n246) );
  HS65_LH_DFPRQNX9 \registers_reg[8][9]  ( .D(n1667), .CP(clk), .RN(n2840), 
        .QN(n247) );
  HS65_LH_DFPRQNX9 \registers_reg[8][8]  ( .D(n1666), .CP(clk), .RN(n2840), 
        .QN(n248) );
  HS65_LH_DFPRQNX9 \registers_reg[8][7]  ( .D(n1665), .CP(clk), .RN(n2840), 
        .QN(n249) );
  HS65_LH_DFPRQNX9 \registers_reg[8][6]  ( .D(n1664), .CP(clk), .RN(n2840), 
        .QN(n250) );
  HS65_LH_DFPRQNX9 \registers_reg[8][5]  ( .D(n1663), .CP(clk), .RN(n2840), 
        .QN(n251) );
  HS65_LH_DFPRQNX9 \registers_reg[8][4]  ( .D(n1662), .CP(clk), .RN(n2840), 
        .QN(n252) );
  HS65_LH_DFPRQNX9 \registers_reg[8][3]  ( .D(n1661), .CP(clk), .RN(n2840), 
        .QN(n253) );
  HS65_LH_DFPRQNX9 \registers_reg[8][2]  ( .D(n1660), .CP(clk), .RN(n2840), 
        .QN(n254) );
  HS65_LH_DFPRQNX9 \registers_reg[8][1]  ( .D(n1659), .CP(clk), .RN(n2840), 
        .QN(n255) );
  HS65_LH_DFPRQNX9 \registers_reg[8][0]  ( .D(n1658), .CP(clk), .RN(n2841), 
        .QN(n256) );
  HS65_LH_AND2X4 U3 ( .A(n1393), .B(n1394), .Z(n257) );
  HS65_LH_AND2X4 U4 ( .A(n1396), .B(n1394), .Z(n258) );
  HS65_LH_AND2X4 U5 ( .A(n1398), .B(n1394), .Z(n259) );
  HS65_LH_AND2X4 U6 ( .A(n1406), .B(n1394), .Z(n260) );
  HS65_LH_AND2X4 U7 ( .A(n1402), .B(n1394), .Z(n261) );
  HS65_LH_AND2X4 U8 ( .A(n1404), .B(n1394), .Z(n262) );
  HS65_LH_AND2X4 U9 ( .A(n1400), .B(n1394), .Z(n263) );
  HS65_LH_AND2X4 U10 ( .A(n1408), .B(n1398), .Z(n264) );
  HS65_LH_AND2X4 U11 ( .A(n1408), .B(n1402), .Z(n265) );
  HS65_LH_AND2X4 U12 ( .A(n1408), .B(n1396), .Z(n266) );
  HS65_LH_AND2X4 U13 ( .A(n1408), .B(n1400), .Z(n267) );
  HS65_LH_AND2X4 U14 ( .A(n1417), .B(n1402), .Z(n268) );
  HS65_LH_AND2X4 U15 ( .A(n1417), .B(n1400), .Z(n269) );
  HS65_LH_AND2X4 U16 ( .A(n1426), .B(n1404), .Z(n270) );
  HS65_LH_AND2X4 U17 ( .A(n1417), .B(n1404), .Z(n271) );
  HS65_LH_AND2X4 U18 ( .A(n1426), .B(n1406), .Z(n272) );
  HS65_LH_AND2X4 U19 ( .A(n1417), .B(n1406), .Z(n273) );
  HS65_LH_AND2X4 U20 ( .A(n1426), .B(n1393), .Z(n274) );
  HS65_LH_AND2X4 U21 ( .A(n1417), .B(n1398), .Z(n275) );
  HS65_LH_AND2X4 U22 ( .A(n1417), .B(n1393), .Z(n276) );
  HS65_LH_AND2X4 U23 ( .A(n1417), .B(n1396), .Z(n277) );
  HS65_LH_AND2X4 U24 ( .A(n861), .B(n841), .Z(n380) );
  HS65_LH_AND2X4 U25 ( .A(n849), .B(n841), .Z(n358) );
  HS65_LH_AND2X4 U26 ( .A(n1389), .B(n1369), .Z(n908) );
  HS65_LH_AND2X4 U27 ( .A(n1377), .B(n1369), .Z(n886) );
  HS65_LH_AND2X4 U28 ( .A(n857), .B(n841), .Z(n365) );
  HS65_LH_AND2X4 U29 ( .A(n1385), .B(n1369), .Z(n893) );
  HS65_LH_AND2X4 U30 ( .A(n861), .B(n843), .Z(n378) );
  HS65_LH_AND2X4 U31 ( .A(n860), .B(n843), .Z(n379) );
  HS65_LH_AND2X4 U32 ( .A(n861), .B(n846), .Z(n376) );
  HS65_LH_AND2X4 U33 ( .A(n860), .B(n846), .Z(n377) );
  HS65_LH_AND2X4 U34 ( .A(n849), .B(n843), .Z(n356) );
  HS65_LH_AND2X4 U35 ( .A(n848), .B(n843), .Z(n357) );
  HS65_LH_AND2X4 U36 ( .A(n1389), .B(n1371), .Z(n906) );
  HS65_LH_AND2X4 U37 ( .A(n1388), .B(n1371), .Z(n907) );
  HS65_LH_AND2X4 U38 ( .A(n1389), .B(n1374), .Z(n904) );
  HS65_LH_AND2X4 U39 ( .A(n1388), .B(n1374), .Z(n905) );
  HS65_LH_AND2X4 U40 ( .A(n1377), .B(n1371), .Z(n884) );
  HS65_LH_AND2X4 U41 ( .A(n1376), .B(n1371), .Z(n885) );
  HS65_LH_AND2X4 U42 ( .A(n1368), .B(n1374), .Z(n875) );
  HS65_LH_AND2X4 U43 ( .A(n860), .B(n841), .Z(n381) );
  HS65_LH_AND2X4 U44 ( .A(n1388), .B(n1369), .Z(n909) );
  HS65_LH_AND2X4 U45 ( .A(n1376), .B(n1369), .Z(n887) );
  HS65_LH_AND2X4 U46 ( .A(n861), .B(n845), .Z(n374) );
  HS65_LH_AND2X4 U47 ( .A(n860), .B(n845), .Z(n375) );
  HS65_LH_AND2X4 U48 ( .A(n1389), .B(n1373), .Z(n902) );
  HS65_LH_AND2X4 U49 ( .A(n1388), .B(n1373), .Z(n903) );
  HS65_LH_AND2X4 U50 ( .A(n1373), .B(n1384), .Z(n897) );
  HS65_LH_IVX9 U51 ( .A(\regfile_i[WRITE_DATA][6] ), .Z(n2710) );
  HS65_LH_IVX9 U52 ( .A(\regfile_i[WRITE_DATA][7] ), .Z(n2712) );
  HS65_LH_IVX9 U53 ( .A(\regfile_i[WRITE_DATA][8] ), .Z(n2714) );
  HS65_LH_IVX9 U54 ( .A(\regfile_i[WRITE_DATA][10] ), .Z(n2718) );
  HS65_LH_IVX9 U55 ( .A(\regfile_i[WRITE_DATA][11] ), .Z(n2720) );
  HS65_LH_IVX9 U56 ( .A(\regfile_i[WRITE_DATA][12] ), .Z(n2722) );
  HS65_LH_IVX9 U57 ( .A(\regfile_i[WRITE_DATA][13] ), .Z(n2724) );
  HS65_LH_IVX9 U58 ( .A(\regfile_i[WRITE_DATA][14] ), .Z(n2726) );
  HS65_LH_IVX9 U59 ( .A(\regfile_i[WRITE_DATA][15] ), .Z(n2728) );
  HS65_LH_IVX9 U60 ( .A(\regfile_i[WRITE_DATA][16] ), .Z(n2730) );
  HS65_LH_IVX9 U61 ( .A(\regfile_i[WRITE_DATA][17] ), .Z(n2732) );
  HS65_LH_IVX9 U62 ( .A(\regfile_i[WRITE_DATA][18] ), .Z(n2734) );
  HS65_LH_IVX9 U63 ( .A(\regfile_i[WRITE_DATA][19] ), .Z(n2736) );
  HS65_LH_IVX9 U64 ( .A(\regfile_i[WRITE_DATA][20] ), .Z(n2738) );
  HS65_LH_IVX9 U65 ( .A(\regfile_i[WRITE_DATA][21] ), .Z(n2740) );
  HS65_LH_IVX9 U66 ( .A(\regfile_i[WRITE_DATA][22] ), .Z(n2742) );
  HS65_LH_IVX9 U67 ( .A(\regfile_i[WRITE_DATA][23] ), .Z(n2744) );
  HS65_LH_IVX9 U68 ( .A(\regfile_i[WRITE_DATA][24] ), .Z(n2746) );
  HS65_LH_IVX9 U69 ( .A(\regfile_i[WRITE_DATA][25] ), .Z(n2748) );
  HS65_LH_IVX9 U70 ( .A(\regfile_i[WRITE_DATA][26] ), .Z(n2750) );
  HS65_LH_IVX9 U71 ( .A(\regfile_i[WRITE_DATA][27] ), .Z(n2752) );
  HS65_LH_IVX9 U72 ( .A(\regfile_i[WRITE_DATA][28] ), .Z(n2754) );
  HS65_LH_IVX9 U73 ( .A(\regfile_i[WRITE_DATA][29] ), .Z(n2756) );
  HS65_LH_IVX9 U74 ( .A(\regfile_i[WRITE_DATA][30] ), .Z(n2758) );
  HS65_LH_IVX9 U75 ( .A(\regfile_i[WRITE_DATA][31] ), .Z(n2760) );
  HS65_LH_AND2X4 U76 ( .A(n849), .B(n846), .Z(n354) );
  HS65_LH_AND2X4 U77 ( .A(n848), .B(n846), .Z(n355) );
  HS65_LH_AND2X4 U78 ( .A(n1377), .B(n1374), .Z(n882) );
  HS65_LH_AND2X4 U79 ( .A(n1376), .B(n1374), .Z(n883) );
  HS65_LH_AND2X4 U80 ( .A(n840), .B(n846), .Z(n347) );
  HS65_LH_AND2X4 U81 ( .A(n842), .B(n846), .Z(n348) );
  HS65_LH_AND2X4 U82 ( .A(n840), .B(n843), .Z(n342) );
  HS65_LH_AND2X4 U83 ( .A(n842), .B(n843), .Z(n343) );
  HS65_LH_AND2X4 U84 ( .A(n1370), .B(n1374), .Z(n876) );
  HS65_LH_AND2X4 U85 ( .A(n1368), .B(n1371), .Z(n870) );
  HS65_LH_AND2X4 U86 ( .A(n1370), .B(n1371), .Z(n871) );
  HS65_LH_AND2X4 U87 ( .A(n848), .B(n841), .Z(n359) );
  HS65_LH_AND2X4 U88 ( .A(n848), .B(n845), .Z(n353) );
  HS65_LH_AND2X4 U89 ( .A(n1376), .B(n1373), .Z(n881) );
  HS65_LH_AND2X4 U90 ( .A(n841), .B(n856), .Z(n364) );
  HS65_LH_AND2X4 U91 ( .A(n1369), .B(n1384), .Z(n892) );
  HS65_LH_AND2X4 U92 ( .A(n845), .B(n856), .Z(n369) );
  HS65_LH_AND2X4 U93 ( .A(n845), .B(n857), .Z(n370) );
  HS65_LH_AND2X4 U94 ( .A(n1373), .B(n1385), .Z(n898) );
  HS65_LH_IVX9 U95 ( .A(\regfile_i[WRITE_DATA][1] ), .Z(n2700) );
  HS65_LH_IVX9 U96 ( .A(\regfile_i[WRITE_DATA][2] ), .Z(n2702) );
  HS65_LH_IVX9 U97 ( .A(\regfile_i[WRITE_DATA][3] ), .Z(n2704) );
  HS65_LH_IVX9 U98 ( .A(\regfile_i[WRITE_DATA][4] ), .Z(n2706) );
  HS65_LH_IVX9 U99 ( .A(\regfile_i[WRITE_DATA][5] ), .Z(n2708) );
  HS65_LH_IVX9 U100 ( .A(\regfile_i[WRITE_DATA][9] ), .Z(n2716) );
  HS65_LH_IVX9 U101 ( .A(\regfile_i[WRITE_DATA][0] ), .Z(n2698) );
  HS65_LH_IVX9 U102 ( .A(\regfile_i[FORWARD_A] ), .Z(n2893) );
  HS65_LH_NOR3AX2 U103 ( .A(\regfile_i[ADRWRITE][2] ), .B(
        \regfile_i[ADRWRITE][0] ), .C(\regfile_i[ADRWRITE][1] ), .Z(n1400) );
  HS65_LH_NOR3AX2 U104 ( .A(\regfile_i[ADRWRITE][2] ), .B(n2897), .C(
        \regfile_i[ADRWRITE][1] ), .Z(n1402) );
  HS65_LH_NOR3AX2 U105 ( .A(\regfile_i[ADRWRITE][2] ), .B(n2896), .C(
        \regfile_i[ADRWRITE][0] ), .Z(n1404) );
  HS65_LH_NOR3AX2 U106 ( .A(\regfile_i[WR_EN] ), .B(\regfile_i[ADRWRITE][4] ), 
        .C(n2895), .Z(n1408) );
  HS65_LH_NOR3AX2 U107 ( .A(\regfile_i[ADRWRITE][2] ), .B(n2896), .C(n2897), 
        .Z(n1406) );
  HS65_LH_NOR3AX2 U108 ( .A(\regfile_i[WR_EN] ), .B(\regfile_i[ADRWRITE][3] ), 
        .C(\regfile_i[ADRWRITE][4] ), .Z(n1394) );
  HS65_LH_BFX9 U109 ( .A(n2854), .Z(n2826) );
  HS65_LH_BFX9 U110 ( .A(n2847), .Z(n2840) );
  HS65_LH_BFX9 U111 ( .A(n2847), .Z(n2839) );
  HS65_LH_BFX9 U112 ( .A(n2848), .Z(n2837) );
  HS65_LH_BFX9 U113 ( .A(n2848), .Z(n2838) );
  HS65_LH_BFX9 U114 ( .A(n2850), .Z(n2834) );
  HS65_LH_BFX9 U115 ( .A(n2849), .Z(n2835) );
  HS65_LH_BFX9 U116 ( .A(n2849), .Z(n2836) );
  HS65_LH_BFX9 U117 ( .A(n2846), .Z(n2841) );
  HS65_LH_BFX9 U118 ( .A(n2846), .Z(n2842) );
  HS65_LH_BFX9 U119 ( .A(n2845), .Z(n2843) );
  HS65_LH_BFX9 U120 ( .A(n2853), .Z(n2828) );
  HS65_LH_BFX9 U121 ( .A(n2853), .Z(n2827) );
  HS65_LH_BFX9 U122 ( .A(n2852), .Z(n2829) );
  HS65_LH_BFX9 U123 ( .A(n2852), .Z(n2830) );
  HS65_LH_BFX9 U124 ( .A(n2851), .Z(n2831) );
  HS65_LH_BFX9 U125 ( .A(n2851), .Z(n2832) );
  HS65_LH_BFX9 U126 ( .A(n2850), .Z(n2833) );
  HS65_LH_BFX9 U127 ( .A(n2871), .Z(n2791) );
  HS65_LH_BFX9 U128 ( .A(n2872), .Z(n2790) );
  HS65_LH_BFX9 U129 ( .A(n2872), .Z(n2789) );
  HS65_LH_BFX9 U130 ( .A(n2873), .Z(n2788) );
  HS65_LH_BFX9 U131 ( .A(n2874), .Z(n2786) );
  HS65_LH_BFX9 U132 ( .A(n2874), .Z(n2785) );
  HS65_LH_BFX9 U133 ( .A(n2875), .Z(n2784) );
  HS65_LH_BFX9 U134 ( .A(n2873), .Z(n2787) );
  HS65_LH_BFX9 U135 ( .A(n2867), .Z(n2800) );
  HS65_LH_BFX9 U136 ( .A(n2867), .Z(n2799) );
  HS65_LH_BFX9 U137 ( .A(n2868), .Z(n2798) );
  HS65_LH_BFX9 U138 ( .A(n2868), .Z(n2797) );
  HS65_LH_BFX9 U139 ( .A(n2869), .Z(n2795) );
  HS65_LH_BFX9 U140 ( .A(n2870), .Z(n2794) );
  HS65_LH_BFX9 U141 ( .A(n2870), .Z(n2793) );
  HS65_LH_BFX9 U142 ( .A(n2871), .Z(n2792) );
  HS65_LH_BFX9 U143 ( .A(n2869), .Z(n2796) );
  HS65_LH_BFX9 U144 ( .A(n2880), .Z(n2773) );
  HS65_LH_BFX9 U145 ( .A(n2881), .Z(n2772) );
  HS65_LH_BFX9 U146 ( .A(n2881), .Z(n2771) );
  HS65_LH_BFX9 U147 ( .A(n2882), .Z(n2770) );
  HS65_LH_BFX9 U148 ( .A(n2883), .Z(n2768) );
  HS65_LH_BFX9 U149 ( .A(n2883), .Z(n2767) );
  HS65_LH_BFX9 U150 ( .A(n2884), .Z(n2766) );
  HS65_LH_BFX9 U151 ( .A(n2882), .Z(n2769) );
  HS65_LH_BFX9 U152 ( .A(n2876), .Z(n2782) );
  HS65_LH_BFX9 U153 ( .A(n2876), .Z(n2781) );
  HS65_LH_BFX9 U154 ( .A(n2877), .Z(n2780) );
  HS65_LH_BFX9 U155 ( .A(n2877), .Z(n2779) );
  HS65_LH_BFX9 U156 ( .A(n2878), .Z(n2777) );
  HS65_LH_BFX9 U157 ( .A(n2879), .Z(n2776) );
  HS65_LH_BFX9 U158 ( .A(n2879), .Z(n2775) );
  HS65_LH_BFX9 U159 ( .A(n2880), .Z(n2774) );
  HS65_LH_BFX9 U160 ( .A(n2878), .Z(n2778) );
  HS65_LH_BFX9 U161 ( .A(n2875), .Z(n2783) );
  HS65_LH_BFX9 U162 ( .A(n2856), .Z(n2822) );
  HS65_LH_BFX9 U163 ( .A(n2857), .Z(n2820) );
  HS65_LH_BFX9 U164 ( .A(n2857), .Z(n2819) );
  HS65_LH_BFX9 U165 ( .A(n2858), .Z(n2818) );
  HS65_LH_BFX9 U166 ( .A(n2856), .Z(n2821) );
  HS65_LH_BFX9 U167 ( .A(n2855), .Z(n2823) );
  HS65_LH_BFX9 U168 ( .A(n2855), .Z(n2824) );
  HS65_LH_BFX9 U169 ( .A(n2854), .Z(n2825) );
  HS65_LH_BFX9 U170 ( .A(n2866), .Z(n2801) );
  HS65_LH_BFX9 U171 ( .A(n2866), .Z(n2802) );
  HS65_LH_BFX9 U172 ( .A(n2865), .Z(n2803) );
  HS65_LH_BFX9 U173 ( .A(n2865), .Z(n2804) );
  HS65_LH_BFX9 U174 ( .A(n2864), .Z(n2805) );
  HS65_LH_BFX9 U175 ( .A(n2864), .Z(n2806) );
  HS65_LH_BFX9 U176 ( .A(n2863), .Z(n2807) );
  HS65_LH_BFX9 U177 ( .A(n2863), .Z(n2808) );
  HS65_LH_BFX9 U178 ( .A(n2862), .Z(n2809) );
  HS65_LH_BFX9 U179 ( .A(n2862), .Z(n2810) );
  HS65_LH_BFX9 U180 ( .A(n2861), .Z(n2811) );
  HS65_LH_BFX9 U181 ( .A(n2861), .Z(n2812) );
  HS65_LH_BFX9 U182 ( .A(n2860), .Z(n2813) );
  HS65_LH_BFX9 U183 ( .A(n2860), .Z(n2814) );
  HS65_LH_BFX9 U184 ( .A(n2859), .Z(n2815) );
  HS65_LH_BFX9 U185 ( .A(n2859), .Z(n2816) );
  HS65_LH_BFX9 U186 ( .A(n2858), .Z(n2817) );
  HS65_LH_BFX9 U187 ( .A(n2884), .Z(n2765) );
  HS65_LH_BFX9 U188 ( .A(n2845), .Z(n2844) );
  HS65_LH_BFX9 U189 ( .A(n2887), .Z(n2872) );
  HS65_LH_BFX9 U190 ( .A(n2887), .Z(n2874) );
  HS65_LH_BFX9 U191 ( .A(n2887), .Z(n2873) );
  HS65_LH_BFX9 U192 ( .A(n2888), .Z(n2867) );
  HS65_LH_BFX9 U193 ( .A(n2888), .Z(n2868) );
  HS65_LH_BFX9 U194 ( .A(n2887), .Z(n2870) );
  HS65_LH_BFX9 U195 ( .A(n2887), .Z(n2871) );
  HS65_LH_BFX9 U196 ( .A(n2888), .Z(n2869) );
  HS65_LH_BFX9 U197 ( .A(n2885), .Z(n2881) );
  HS65_LH_BFX9 U198 ( .A(n2885), .Z(n2883) );
  HS65_LH_BFX9 U199 ( .A(n2885), .Z(n2882) );
  HS65_LH_BFX9 U200 ( .A(n2886), .Z(n2876) );
  HS65_LH_BFX9 U201 ( .A(n2886), .Z(n2877) );
  HS65_LH_BFX9 U202 ( .A(n2886), .Z(n2879) );
  HS65_LH_BFX9 U203 ( .A(n2885), .Z(n2880) );
  HS65_LH_BFX9 U204 ( .A(n2886), .Z(n2878) );
  HS65_LH_BFX9 U205 ( .A(n2886), .Z(n2875) );
  HS65_LH_BFX9 U206 ( .A(n2890), .Z(n2857) );
  HS65_LH_BFX9 U207 ( .A(n2890), .Z(n2856) );
  HS65_LH_BFX9 U208 ( .A(n2890), .Z(n2855) );
  HS65_LH_BFX9 U209 ( .A(n2888), .Z(n2866) );
  HS65_LH_BFX9 U210 ( .A(n2888), .Z(n2865) );
  HS65_LH_BFX9 U211 ( .A(n2889), .Z(n2864) );
  HS65_LH_BFX9 U212 ( .A(n2889), .Z(n2863) );
  HS65_LH_BFX9 U213 ( .A(n2889), .Z(n2862) );
  HS65_LH_BFX9 U214 ( .A(n2889), .Z(n2861) );
  HS65_LH_BFX9 U215 ( .A(n2889), .Z(n2860) );
  HS65_LH_BFX9 U216 ( .A(n2890), .Z(n2859) );
  HS65_LH_BFX9 U217 ( .A(n2890), .Z(n2858) );
  HS65_LH_BFX9 U218 ( .A(n2885), .Z(n2884) );
  HS65_LH_BFX9 U219 ( .A(n2892), .Z(n2847) );
  HS65_LH_BFX9 U220 ( .A(n2892), .Z(n2848) );
  HS65_LH_BFX9 U221 ( .A(n2892), .Z(n2849) );
  HS65_LH_BFX9 U222 ( .A(n2892), .Z(n2846) );
  HS65_LH_BFX9 U223 ( .A(n2892), .Z(n2845) );
  HS65_LH_BFX9 U224 ( .A(n2891), .Z(n2854) );
  HS65_LH_BFX9 U225 ( .A(n2891), .Z(n2853) );
  HS65_LH_BFX9 U226 ( .A(n2891), .Z(n2852) );
  HS65_LH_BFX9 U227 ( .A(n2891), .Z(n2851) );
  HS65_LH_BFX9 U228 ( .A(n2891), .Z(n2850) );
  HS65_LH_BFX9 U229 ( .A(n2761), .Z(n2887) );
  HS65_LH_BFX9 U230 ( .A(n2761), .Z(n2886) );
  HS65_LH_BFX9 U231 ( .A(n2762), .Z(n2888) );
  HS65_LH_BFX9 U232 ( .A(n2762), .Z(n2889) );
  HS65_LH_BFX9 U233 ( .A(n2762), .Z(n2890) );
  HS65_LH_BFX9 U234 ( .A(n2761), .Z(n2885) );
  HS65_LH_BFX9 U235 ( .A(n2763), .Z(n2892) );
  HS65_LH_BFX9 U236 ( .A(n2763), .Z(n2891) );
  HS65_LH_BFX9 U237 ( .A(n908), .Z(n2514) );
  HS65_LH_BFX9 U238 ( .A(n886), .Z(n2562) );
  HS65_LH_BFX9 U239 ( .A(n908), .Z(n2515) );
  HS65_LH_BFX9 U240 ( .A(n886), .Z(n2563) );
  HS65_LH_BFX9 U241 ( .A(n380), .Z(n2607) );
  HS65_LH_BFX9 U242 ( .A(n358), .Z(n2655) );
  HS65_LH_BFX9 U243 ( .A(n380), .Z(n2608) );
  HS65_LH_BFX9 U244 ( .A(n358), .Z(n2656) );
  HS65_LH_BFX9 U245 ( .A(n380), .Z(n2609) );
  HS65_LH_BFX9 U246 ( .A(n358), .Z(n2657) );
  HS65_LH_BFX9 U247 ( .A(n908), .Z(n2516) );
  HS65_LH_BFX9 U248 ( .A(n886), .Z(n2564) );
  HS65_LH_BFX9 U249 ( .A(n893), .Z(n2553) );
  HS65_LH_BFX9 U250 ( .A(n893), .Z(n2554) );
  HS65_LH_BFX9 U251 ( .A(n345), .Z(n2688) );
  HS65_LH_BFX9 U252 ( .A(n345), .Z(n2689) );
  HS65_LH_BFX9 U253 ( .A(n365), .Z(n2646) );
  HS65_LH_BFX9 U254 ( .A(n365), .Z(n2647) );
  HS65_LH_BFX9 U255 ( .A(n873), .Z(n2595) );
  HS65_LH_BFX9 U256 ( .A(n873), .Z(n2596) );
  HS65_LH_BFX9 U257 ( .A(n345), .Z(n2690) );
  HS65_LH_BFX9 U258 ( .A(n873), .Z(n2597) );
  HS65_LH_BFX9 U259 ( .A(n893), .Z(n2555) );
  HS65_LH_BFX9 U260 ( .A(n365), .Z(n2648) );
  HS65_LH_IVX9 U261 ( .A(n2473), .Z(n2472) );
  HS65_LH_IVX9 U262 ( .A(n2473), .Z(n2471) );
  HS65_LH_IVX9 U263 ( .A(n2468), .Z(n2467) );
  HS65_LH_IVX9 U264 ( .A(n2468), .Z(n2466) );
  HS65_LH_IVX9 U265 ( .A(n2443), .Z(n2442) );
  HS65_LH_IVX9 U266 ( .A(n2443), .Z(n2441) );
  HS65_LH_IVX9 U267 ( .A(n2438), .Z(n2437) );
  HS65_LH_IVX9 U268 ( .A(n2438), .Z(n2436) );
  HS65_LH_IVX9 U269 ( .A(n300), .Z(n299) );
  HS65_LH_IVX9 U270 ( .A(n300), .Z(n298) );
  HS65_LH_BFX9 U271 ( .A(n259), .Z(n2499) );
  HS65_LH_BFX9 U272 ( .A(n263), .Z(n2494) );
  HS65_LH_BFX9 U273 ( .A(n261), .Z(n2489) );
  HS65_LH_BFX9 U274 ( .A(n262), .Z(n2484) );
  HS65_LH_BFX9 U275 ( .A(n260), .Z(n2479) );
  HS65_LH_BFX9 U276 ( .A(n266), .Z(n2464) );
  HS65_LH_BFX9 U277 ( .A(n264), .Z(n2459) );
  HS65_LH_BFX9 U278 ( .A(n267), .Z(n2454) );
  HS65_LH_BFX9 U279 ( .A(n265), .Z(n2449) );
  HS65_LH_BFX9 U280 ( .A(n269), .Z(n1412) );
  HS65_LH_BFX9 U281 ( .A(n268), .Z(n1401) );
  HS65_LH_BFX9 U282 ( .A(n271), .Z(n880) );
  HS65_LH_BFX9 U283 ( .A(n270), .Z(n296) );
  HS65_LH_IVX9 U284 ( .A(n2463), .Z(n2462) );
  HS65_LH_IVX9 U285 ( .A(n2463), .Z(n2461) );
  HS65_LH_IVX9 U286 ( .A(n2458), .Z(n2457) );
  HS65_LH_IVX9 U287 ( .A(n2458), .Z(n2456) );
  HS65_LH_IVX9 U288 ( .A(n2453), .Z(n2452) );
  HS65_LH_IVX9 U289 ( .A(n2453), .Z(n2451) );
  HS65_LH_IVX9 U290 ( .A(n2448), .Z(n2447) );
  HS65_LH_IVX9 U291 ( .A(n2448), .Z(n2446) );
  HS65_LH_IVX9 U292 ( .A(n2508), .Z(n2507) );
  HS65_LH_IVX9 U293 ( .A(n2508), .Z(n2506) );
  HS65_LH_IVX9 U294 ( .A(n2503), .Z(n2502) );
  HS65_LH_IVX9 U295 ( .A(n2503), .Z(n2501) );
  HS65_LH_IVX9 U296 ( .A(n2498), .Z(n2497) );
  HS65_LH_IVX9 U297 ( .A(n2498), .Z(n2496) );
  HS65_LH_IVX9 U298 ( .A(n2493), .Z(n2492) );
  HS65_LH_IVX9 U299 ( .A(n2493), .Z(n2491) );
  HS65_LH_IVX9 U300 ( .A(n2488), .Z(n2487) );
  HS65_LH_IVX9 U301 ( .A(n2488), .Z(n2486) );
  HS65_LH_IVX9 U302 ( .A(n2483), .Z(n2482) );
  HS65_LH_IVX9 U303 ( .A(n2483), .Z(n2481) );
  HS65_LH_IVX9 U304 ( .A(n2478), .Z(n2477) );
  HS65_LH_IVX9 U305 ( .A(n2478), .Z(n2476) );
  HS65_LH_IVX9 U306 ( .A(n2428), .Z(n2427) );
  HS65_LH_IVX9 U307 ( .A(n2428), .Z(n2426) );
  HS65_LH_IVX9 U308 ( .A(n1427), .Z(n1424) );
  HS65_LH_IVX9 U309 ( .A(n1427), .Z(n1423) );
  HS65_LH_IVX9 U310 ( .A(n1420), .Z(n1419) );
  HS65_LH_IVX9 U311 ( .A(n1420), .Z(n1418) );
  HS65_LH_IVX9 U312 ( .A(n1411), .Z(n1410) );
  HS65_LH_IVX9 U313 ( .A(n1411), .Z(n1405) );
  HS65_LH_IVX9 U314 ( .A(n1399), .Z(n1397) );
  HS65_LH_IVX9 U315 ( .A(n1399), .Z(n1395) );
  HS65_LH_IVX9 U316 ( .A(n352), .Z(n334) );
  HS65_LH_IVX9 U317 ( .A(n352), .Z(n333) );
  HS65_LH_IVX9 U318 ( .A(n320), .Z(n319) );
  HS65_LH_IVX9 U319 ( .A(n320), .Z(n318) );
  HS65_LH_IVX9 U320 ( .A(n295), .Z(n294) );
  HS65_LH_IVX9 U321 ( .A(n295), .Z(n293) );
  HS65_LH_IVX9 U322 ( .A(n330), .Z(n329) );
  HS65_LH_IVX9 U323 ( .A(n330), .Z(n328) );
  HS65_LH_IVX9 U324 ( .A(n290), .Z(n289) );
  HS65_LH_IVX9 U325 ( .A(n290), .Z(n288) );
  HS65_LH_BFX9 U326 ( .A(n259), .Z(n2500) );
  HS65_LH_BFX9 U327 ( .A(n263), .Z(n2495) );
  HS65_LH_BFX9 U328 ( .A(n261), .Z(n2490) );
  HS65_LH_BFX9 U329 ( .A(n262), .Z(n2485) );
  HS65_LH_BFX9 U330 ( .A(n266), .Z(n2465) );
  HS65_LH_BFX9 U331 ( .A(n264), .Z(n2460) );
  HS65_LH_BFX9 U332 ( .A(n267), .Z(n2455) );
  HS65_LH_BFX9 U333 ( .A(n265), .Z(n2450) );
  HS65_LH_IVX9 U334 ( .A(n305), .Z(n304) );
  HS65_LH_IVX9 U335 ( .A(n305), .Z(n303) );
  HS65_LH_IVX9 U336 ( .A(n315), .Z(n314) );
  HS65_LH_IVX9 U337 ( .A(n315), .Z(n313) );
  HS65_LH_IVX9 U338 ( .A(n310), .Z(n309) );
  HS65_LH_IVX9 U339 ( .A(n310), .Z(n308) );
  HS65_LH_BFX9 U340 ( .A(n257), .Z(n2509) );
  HS65_LH_BFX9 U341 ( .A(n258), .Z(n2504) );
  HS65_LH_BFX9 U342 ( .A(n276), .Z(n2429) );
  HS65_LH_BFX9 U343 ( .A(n277), .Z(n1432) );
  HS65_LH_BFX9 U344 ( .A(n275), .Z(n1421) );
  HS65_LH_BFX9 U345 ( .A(n274), .Z(n321) );
  HS65_LH_BFX9 U346 ( .A(n273), .Z(n331) );
  HS65_LH_BFX9 U347 ( .A(n272), .Z(n291) );
  HS65_LH_BFX9 U348 ( .A(n2435), .Z(n2433) );
  HS65_LH_BFX9 U349 ( .A(n327), .Z(n325) );
  HS65_LH_IVX9 U350 ( .A(n2432), .Z(n2431) );
  HS65_LH_IVX9 U351 ( .A(n324), .Z(n323) );
  HS65_LH_BFX9 U352 ( .A(n257), .Z(n2510) );
  HS65_LH_BFX9 U353 ( .A(n258), .Z(n2505) );
  HS65_LH_BFX9 U354 ( .A(n260), .Z(n2480) );
  HS65_LH_BFX9 U355 ( .A(n269), .Z(n1413) );
  HS65_LH_BFX9 U356 ( .A(n268), .Z(n1403) );
  HS65_LH_BFX9 U357 ( .A(n271), .Z(n1392) );
  HS65_LH_BFX9 U358 ( .A(n270), .Z(n297) );
  HS65_LH_BFX9 U359 ( .A(n2428), .Z(n2430) );
  HS65_LH_BFX9 U360 ( .A(n1427), .Z(n1433) );
  HS65_LH_BFX9 U361 ( .A(n1420), .Z(n1422) );
  HS65_LH_BFX9 U362 ( .A(n320), .Z(n322) );
  HS65_LH_BFX9 U363 ( .A(n273), .Z(n332) );
  HS65_LH_BFX9 U364 ( .A(n272), .Z(n292) );
  HS65_LH_BFX9 U365 ( .A(n2432), .Z(n2434) );
  HS65_LH_BFX9 U366 ( .A(n324), .Z(n326) );
  HS65_LH_BFX9 U367 ( .A(n2764), .Z(n2762) );
  HS65_LH_BFX9 U368 ( .A(n2764), .Z(n2761) );
  HS65_LH_BFX9 U369 ( .A(n2764), .Z(n2763) );
  HS65_LH_BFX9 U370 ( .A(n897), .Z(n2544) );
  HS65_LH_BFX9 U371 ( .A(n892), .Z(n2556) );
  HS65_LH_BFX9 U372 ( .A(n897), .Z(n2545) );
  HS65_LH_BFX9 U373 ( .A(n892), .Z(n2557) );
  HS65_LH_BFX9 U374 ( .A(n875), .Z(n2589) );
  HS65_LH_BFX9 U375 ( .A(n870), .Z(n2601) );
  HS65_LH_BFX9 U376 ( .A(n875), .Z(n2590) );
  HS65_LH_BFX9 U377 ( .A(n870), .Z(n2602) );
  HS65_LH_BFX9 U378 ( .A(n369), .Z(n2637) );
  HS65_LH_BFX9 U379 ( .A(n369), .Z(n2638) );
  HS65_LH_BFX9 U380 ( .A(n347), .Z(n2682) );
  HS65_LH_BFX9 U381 ( .A(n347), .Z(n2683) );
  HS65_LH_BFX9 U382 ( .A(n372), .Z(n2631) );
  HS65_LH_BFX9 U383 ( .A(n372), .Z(n2632) );
  HS65_LH_BFX9 U384 ( .A(n904), .Z(n2526) );
  HS65_LH_BFX9 U385 ( .A(n904), .Z(n2527) );
  HS65_LH_BFX9 U386 ( .A(n906), .Z(n2520) );
  HS65_LH_BFX9 U387 ( .A(n902), .Z(n2532) );
  HS65_LH_BFX9 U388 ( .A(n884), .Z(n2568) );
  HS65_LH_BFX9 U389 ( .A(n906), .Z(n2521) );
  HS65_LH_BFX9 U390 ( .A(n902), .Z(n2533) );
  HS65_LH_BFX9 U391 ( .A(n884), .Z(n2569) );
  HS65_LH_BFX9 U392 ( .A(n907), .Z(n2517) );
  HS65_LH_BFX9 U393 ( .A(n903), .Z(n2529) );
  HS65_LH_BFX9 U394 ( .A(n885), .Z(n2565) );
  HS65_LH_BFX9 U395 ( .A(n907), .Z(n2518) );
  HS65_LH_BFX9 U396 ( .A(n903), .Z(n2530) );
  HS65_LH_BFX9 U397 ( .A(n885), .Z(n2566) );
  HS65_LH_BFX9 U398 ( .A(n909), .Z(n2511) );
  HS65_LH_BFX9 U399 ( .A(n905), .Z(n2523) );
  HS65_LH_BFX9 U400 ( .A(n887), .Z(n2559) );
  HS65_LH_BFX9 U401 ( .A(n909), .Z(n2512) );
  HS65_LH_BFX9 U402 ( .A(n905), .Z(n2524) );
  HS65_LH_BFX9 U403 ( .A(n887), .Z(n2560) );
  HS65_LH_BFX9 U404 ( .A(n381), .Z(n2604) );
  HS65_LH_BFX9 U405 ( .A(n377), .Z(n2616) );
  HS65_LH_BFX9 U406 ( .A(n359), .Z(n2652) );
  HS65_LH_BFX9 U407 ( .A(n381), .Z(n2605) );
  HS65_LH_BFX9 U408 ( .A(n377), .Z(n2617) );
  HS65_LH_BFX9 U409 ( .A(n359), .Z(n2653) );
  HS65_LH_BFX9 U410 ( .A(n379), .Z(n2610) );
  HS65_LH_BFX9 U411 ( .A(n375), .Z(n2622) );
  HS65_LH_BFX9 U412 ( .A(n357), .Z(n2658) );
  HS65_LH_BFX9 U413 ( .A(n379), .Z(n2611) );
  HS65_LH_BFX9 U414 ( .A(n375), .Z(n2623) );
  HS65_LH_BFX9 U415 ( .A(n357), .Z(n2659) );
  HS65_LH_BFX9 U416 ( .A(n378), .Z(n2613) );
  HS65_LH_BFX9 U417 ( .A(n374), .Z(n2625) );
  HS65_LH_BFX9 U418 ( .A(n356), .Z(n2661) );
  HS65_LH_BFX9 U419 ( .A(n378), .Z(n2614) );
  HS65_LH_BFX9 U420 ( .A(n374), .Z(n2626) );
  HS65_LH_BFX9 U421 ( .A(n356), .Z(n2662) );
  HS65_LH_BFX9 U422 ( .A(n376), .Z(n2619) );
  HS65_LH_BFX9 U423 ( .A(n376), .Z(n2620) );
  HS65_LH_BFX9 U424 ( .A(n897), .Z(n2546) );
  HS65_LH_BFX9 U425 ( .A(n875), .Z(n2591) );
  HS65_LH_BFX9 U426 ( .A(n907), .Z(n2519) );
  HS65_LH_BFX9 U427 ( .A(n903), .Z(n2531) );
  HS65_LH_BFX9 U428 ( .A(n885), .Z(n2567) );
  HS65_LH_BFX9 U429 ( .A(n909), .Z(n2513) );
  HS65_LH_BFX9 U430 ( .A(n905), .Z(n2525) );
  HS65_LH_BFX9 U431 ( .A(n887), .Z(n2561) );
  HS65_LH_BFX9 U432 ( .A(n381), .Z(n2606) );
  HS65_LH_BFX9 U433 ( .A(n377), .Z(n2618) );
  HS65_LH_BFX9 U434 ( .A(n359), .Z(n2654) );
  HS65_LH_BFX9 U435 ( .A(n379), .Z(n2612) );
  HS65_LH_BFX9 U436 ( .A(n375), .Z(n2624) );
  HS65_LH_BFX9 U437 ( .A(n357), .Z(n2660) );
  HS65_LH_BFX9 U438 ( .A(n378), .Z(n2615) );
  HS65_LH_BFX9 U439 ( .A(n374), .Z(n2627) );
  HS65_LH_BFX9 U440 ( .A(n356), .Z(n2663) );
  HS65_LH_BFX9 U441 ( .A(n376), .Z(n2621) );
  HS65_LH_BFX9 U442 ( .A(n904), .Z(n2528) );
  HS65_LH_BFX9 U443 ( .A(n906), .Z(n2522) );
  HS65_LH_BFX9 U444 ( .A(n902), .Z(n2534) );
  HS65_LH_BFX9 U445 ( .A(n884), .Z(n2570) );
  HS65_LH_NAND2X7 U446 ( .A(n842), .B(n841), .Z(n345) );
  HS65_LH_NAND2X7 U447 ( .A(n1370), .B(n1369), .Z(n873) );
  HS65_LH_BFX9 U448 ( .A(n882), .Z(n2574) );
  HS65_LH_BFX9 U449 ( .A(n883), .Z(n2571) );
  HS65_LH_BFX9 U450 ( .A(n881), .Z(n2577) );
  HS65_LH_BFX9 U451 ( .A(n882), .Z(n2575) );
  HS65_LH_BFX9 U452 ( .A(n883), .Z(n2572) );
  HS65_LH_BFX9 U453 ( .A(n881), .Z(n2578) );
  HS65_LH_BFX9 U454 ( .A(n373), .Z(n2628) );
  HS65_LH_BFX9 U455 ( .A(n368), .Z(n2640) );
  HS65_LH_BFX9 U456 ( .A(n373), .Z(n2629) );
  HS65_LH_BFX9 U457 ( .A(n368), .Z(n2641) );
  HS65_LH_BFX9 U458 ( .A(n346), .Z(n2685) );
  HS65_LH_BFX9 U459 ( .A(n346), .Z(n2686) );
  HS65_LH_BFX9 U460 ( .A(n354), .Z(n2667) );
  HS65_LH_BFX9 U461 ( .A(n355), .Z(n2664) );
  HS65_LH_BFX9 U462 ( .A(n353), .Z(n2670) );
  HS65_LH_BFX9 U463 ( .A(n354), .Z(n2668) );
  HS65_LH_BFX9 U464 ( .A(n355), .Z(n2665) );
  HS65_LH_BFX9 U465 ( .A(n353), .Z(n2671) );
  HS65_LH_BFX9 U466 ( .A(n351), .Z(n2673) );
  HS65_LH_BFX9 U467 ( .A(n351), .Z(n2674) );
  HS65_LH_BFX9 U468 ( .A(n898), .Z(n2541) );
  HS65_LH_BFX9 U469 ( .A(n898), .Z(n2542) );
  HS65_LH_BFX9 U470 ( .A(n876), .Z(n2586) );
  HS65_LH_BFX9 U471 ( .A(n871), .Z(n2598) );
  HS65_LH_BFX9 U472 ( .A(n876), .Z(n2587) );
  HS65_LH_BFX9 U473 ( .A(n871), .Z(n2599) );
  HS65_LH_BFX9 U474 ( .A(n364), .Z(n2649) );
  HS65_LH_BFX9 U475 ( .A(n364), .Z(n2650) );
  HS65_LH_BFX9 U476 ( .A(n342), .Z(n2694) );
  HS65_LH_BFX9 U477 ( .A(n342), .Z(n2695) );
  HS65_LH_BFX9 U478 ( .A(n901), .Z(n2535) );
  HS65_LH_BFX9 U479 ( .A(n896), .Z(n2547) );
  HS65_LH_BFX9 U480 ( .A(n901), .Z(n2536) );
  HS65_LH_BFX9 U481 ( .A(n896), .Z(n2548) );
  HS65_LH_BFX9 U482 ( .A(n367), .Z(n2643) );
  HS65_LH_BFX9 U483 ( .A(n367), .Z(n2644) );
  HS65_LH_BFX9 U484 ( .A(n874), .Z(n2592) );
  HS65_LH_BFX9 U485 ( .A(n874), .Z(n2593) );
  HS65_LH_BFX9 U486 ( .A(n370), .Z(n2634) );
  HS65_LH_BFX9 U487 ( .A(n370), .Z(n2635) );
  HS65_LH_BFX9 U488 ( .A(n348), .Z(n2679) );
  HS65_LH_BFX9 U489 ( .A(n343), .Z(n2691) );
  HS65_LH_BFX9 U490 ( .A(n348), .Z(n2680) );
  HS65_LH_BFX9 U491 ( .A(n343), .Z(n2692) );
  HS65_LH_BFX9 U492 ( .A(n879), .Z(n2580) );
  HS65_LH_BFX9 U493 ( .A(n879), .Z(n2581) );
  HS65_LH_BFX9 U494 ( .A(n350), .Z(n2676) );
  HS65_LH_BFX9 U495 ( .A(n350), .Z(n2677) );
  HS65_LH_BFX9 U496 ( .A(n900), .Z(n2538) );
  HS65_LH_BFX9 U497 ( .A(n895), .Z(n2550) );
  HS65_LH_BFX9 U498 ( .A(n900), .Z(n2539) );
  HS65_LH_BFX9 U499 ( .A(n895), .Z(n2551) );
  HS65_LH_BFX9 U500 ( .A(n878), .Z(n2583) );
  HS65_LH_BFX9 U501 ( .A(n878), .Z(n2584) );
  HS65_LH_BFX9 U502 ( .A(n354), .Z(n2669) );
  HS65_LH_BFX9 U503 ( .A(n355), .Z(n2666) );
  HS65_LH_BFX9 U504 ( .A(n353), .Z(n2672) );
  HS65_LH_BFX9 U505 ( .A(n369), .Z(n2639) );
  HS65_LH_BFX9 U506 ( .A(n364), .Z(n2651) );
  HS65_LH_BFX9 U507 ( .A(n347), .Z(n2684) );
  HS65_LH_BFX9 U508 ( .A(n342), .Z(n2696) );
  HS65_LH_BFX9 U509 ( .A(n372), .Z(n2633) );
  HS65_LH_BFX9 U510 ( .A(n367), .Z(n2645) );
  HS65_LH_BFX9 U511 ( .A(n350), .Z(n2678) );
  HS65_LH_BFX9 U512 ( .A(n878), .Z(n2585) );
  HS65_LH_IVX9 U513 ( .A(n2710), .Z(n2709) );
  HS65_LH_IVX9 U514 ( .A(n2712), .Z(n2711) );
  HS65_LH_IVX9 U515 ( .A(n2714), .Z(n2713) );
  HS65_LH_IVX9 U516 ( .A(n2716), .Z(n2715) );
  HS65_LH_IVX9 U517 ( .A(n2718), .Z(n2717) );
  HS65_LH_IVX9 U518 ( .A(n2720), .Z(n2719) );
  HS65_LH_IVX9 U519 ( .A(n2722), .Z(n2721) );
  HS65_LH_IVX9 U520 ( .A(n2724), .Z(n2723) );
  HS65_LH_IVX9 U521 ( .A(n2726), .Z(n2725) );
  HS65_LH_IVX9 U522 ( .A(n2728), .Z(n2727) );
  HS65_LH_IVX9 U523 ( .A(n2730), .Z(n2729) );
  HS65_LH_IVX9 U524 ( .A(n2732), .Z(n2731) );
  HS65_LH_IVX9 U525 ( .A(n2734), .Z(n2733) );
  HS65_LH_IVX9 U526 ( .A(n2736), .Z(n2735) );
  HS65_LH_IVX9 U527 ( .A(n2738), .Z(n2737) );
  HS65_LH_IVX9 U528 ( .A(n2740), .Z(n2739) );
  HS65_LH_IVX9 U529 ( .A(n2742), .Z(n2741) );
  HS65_LH_IVX9 U530 ( .A(n2744), .Z(n2743) );
  HS65_LH_IVX9 U531 ( .A(n2746), .Z(n2745) );
  HS65_LH_IVX9 U532 ( .A(n2748), .Z(n2747) );
  HS65_LH_IVX9 U533 ( .A(n2750), .Z(n2749) );
  HS65_LH_IVX9 U534 ( .A(n2752), .Z(n2751) );
  HS65_LH_IVX9 U535 ( .A(n2754), .Z(n2753) );
  HS65_LH_IVX9 U536 ( .A(n2756), .Z(n2755) );
  HS65_LH_IVX9 U537 ( .A(n2758), .Z(n2757) );
  HS65_LH_IVX9 U538 ( .A(n2760), .Z(n2759) );
  HS65_LH_BFX9 U539 ( .A(n900), .Z(n2540) );
  HS65_LH_BFX9 U540 ( .A(n895), .Z(n2552) );
  HS65_LH_BFX9 U541 ( .A(n882), .Z(n2576) );
  HS65_LH_BFX9 U542 ( .A(n883), .Z(n2573) );
  HS65_LH_BFX9 U543 ( .A(n881), .Z(n2579) );
  HS65_LH_IVX9 U544 ( .A(n2698), .Z(n2697) );
  HS65_LH_IVX9 U545 ( .A(n2700), .Z(n2699) );
  HS65_LH_IVX9 U546 ( .A(n2702), .Z(n2701) );
  HS65_LH_IVX9 U547 ( .A(n2704), .Z(n2703) );
  HS65_LH_IVX9 U548 ( .A(n2706), .Z(n2705) );
  HS65_LH_IVX9 U549 ( .A(n2708), .Z(n2707) );
  HS65_LH_BFX9 U550 ( .A(n892), .Z(n2558) );
  HS65_LH_BFX9 U551 ( .A(n870), .Z(n2603) );
  HS65_LH_BFX9 U552 ( .A(n346), .Z(n2687) );
  HS65_LH_BFX9 U553 ( .A(n351), .Z(n2675) );
  HS65_LH_BFX9 U554 ( .A(n373), .Z(n2630) );
  HS65_LH_BFX9 U555 ( .A(n368), .Z(n2642) );
  HS65_LH_BFX9 U556 ( .A(n874), .Z(n2594) );
  HS65_LH_BFX9 U557 ( .A(n879), .Z(n2582) );
  HS65_LH_BFX9 U558 ( .A(n901), .Z(n2537) );
  HS65_LH_BFX9 U559 ( .A(n896), .Z(n2549) );
  HS65_LH_BFX9 U560 ( .A(n898), .Z(n2543) );
  HS65_LH_BFX9 U561 ( .A(n876), .Z(n2588) );
  HS65_LH_BFX9 U562 ( .A(n871), .Z(n2600) );
  HS65_LH_BFX9 U563 ( .A(n370), .Z(n2636) );
  HS65_LH_BFX9 U564 ( .A(n348), .Z(n2681) );
  HS65_LH_BFX9 U565 ( .A(n343), .Z(n2693) );
  HS65_LH_BFX9 U566 ( .A(n257), .Z(n2508) );
  HS65_LH_BFX9 U567 ( .A(n258), .Z(n2503) );
  HS65_LH_BFX9 U568 ( .A(n261), .Z(n2488) );
  HS65_LH_BFX9 U569 ( .A(n262), .Z(n2483) );
  HS65_LH_BFX9 U570 ( .A(n1407), .Z(n2473) );
  HS65_LH_BFX9 U571 ( .A(n1409), .Z(n2468) );
  HS65_LH_BFX9 U572 ( .A(n1414), .Z(n2443) );
  HS65_LH_BFX9 U573 ( .A(n1415), .Z(n2438) );
  HS65_LH_BFX9 U574 ( .A(n1431), .Z(n300) );
  HS65_LH_BFX9 U575 ( .A(n259), .Z(n2498) );
  HS65_LH_BFX9 U576 ( .A(n263), .Z(n2493) );
  HS65_LH_BFX9 U577 ( .A(n260), .Z(n2478) );
  HS65_LH_BFX9 U578 ( .A(n266), .Z(n2463) );
  HS65_LH_BFX9 U579 ( .A(n264), .Z(n2458) );
  HS65_LH_BFX9 U580 ( .A(n267), .Z(n2453) );
  HS65_LH_BFX9 U581 ( .A(n265), .Z(n2448) );
  HS65_LH_BFX9 U582 ( .A(n269), .Z(n1411) );
  HS65_LH_BFX9 U583 ( .A(n268), .Z(n1399) );
  HS65_LH_BFX9 U584 ( .A(n271), .Z(n352) );
  HS65_LH_BFX9 U585 ( .A(n270), .Z(n295) );
  HS65_LH_BFX9 U586 ( .A(n276), .Z(n2428) );
  HS65_LH_BFX9 U587 ( .A(n277), .Z(n1427) );
  HS65_LH_BFX9 U588 ( .A(n275), .Z(n1420) );
  HS65_LH_BFX9 U589 ( .A(n274), .Z(n320) );
  HS65_LH_BFX9 U590 ( .A(n273), .Z(n330) );
  HS65_LH_BFX9 U591 ( .A(n272), .Z(n290) );
  HS65_LH_BFX9 U592 ( .A(n1428), .Z(n315) );
  HS65_LH_BFX9 U593 ( .A(n1429), .Z(n310) );
  HS65_LH_BFX9 U594 ( .A(n1430), .Z(n305) );
  HS65_LH_BFX9 U595 ( .A(n1407), .Z(n2474) );
  HS65_LH_BFX9 U596 ( .A(n1409), .Z(n2469) );
  HS65_LH_BFX9 U597 ( .A(n1414), .Z(n2444) );
  HS65_LH_BFX9 U598 ( .A(n1415), .Z(n2439) );
  HS65_LH_BFX9 U599 ( .A(n1428), .Z(n316) );
  HS65_LH_BFX9 U600 ( .A(n1429), .Z(n311) );
  HS65_LH_BFX9 U601 ( .A(n1430), .Z(n306) );
  HS65_LH_BFX9 U602 ( .A(n1431), .Z(n301) );
  HS65_LH_BFX9 U603 ( .A(n2435), .Z(n2432) );
  HS65_LH_IVX9 U604 ( .A(n1416), .Z(n2435) );
  HS65_LH_BFX9 U605 ( .A(n327), .Z(n324) );
  HS65_LH_IVX9 U606 ( .A(n1425), .Z(n327) );
  HS65_LH_BFX9 U607 ( .A(n1407), .Z(n2475) );
  HS65_LH_BFX9 U608 ( .A(n1409), .Z(n2470) );
  HS65_LH_BFX9 U609 ( .A(n1414), .Z(n2445) );
  HS65_LH_BFX9 U610 ( .A(n1415), .Z(n2440) );
  HS65_LH_BFX9 U611 ( .A(n1428), .Z(n317) );
  HS65_LH_BFX9 U612 ( .A(n1429), .Z(n312) );
  HS65_LH_BFX9 U613 ( .A(n1430), .Z(n307) );
  HS65_LH_BFX9 U614 ( .A(n1431), .Z(n302) );
  HS65_LH_BFX9 U615 ( .A(rst_n), .Z(n2764) );
  HS65_LH_NAND2X7 U616 ( .A(n846), .B(n857), .Z(n372) );
  HS65_LH_NOR2X6 U617 ( .A(n2900), .B(n2899), .Z(n841) );
  HS65_LH_NOR2X6 U618 ( .A(n2905), .B(n2904), .Z(n1369) );
  HS65_LH_AND2X4 U619 ( .A(n859), .B(n2898), .Z(n857) );
  HS65_LH_AND2X4 U620 ( .A(n862), .B(n2898), .Z(n861) );
  HS65_LH_AND2X4 U621 ( .A(n1390), .B(n2903), .Z(n1389) );
  HS65_LH_NOR2X6 U622 ( .A(n2902), .B(n2901), .Z(n859) );
  HS65_LH_NOR2X6 U623 ( .A(n2907), .B(n2906), .Z(n1387) );
  HS65_LH_AND2X4 U624 ( .A(n850), .B(n2898), .Z(n849) );
  HS65_LH_AND2X4 U625 ( .A(n1378), .B(n2903), .Z(n1377) );
  HS65_LH_BFX9 U626 ( .A(n2893), .Z(n280) );
  HS65_LH_BFX9 U627 ( .A(n2894), .Z(n285) );
  HS65_LH_BFX9 U628 ( .A(n2893), .Z(n278) );
  HS65_LH_BFX9 U629 ( .A(n2893), .Z(n279) );
  HS65_LH_BFX9 U630 ( .A(n2894), .Z(n283) );
  HS65_LH_BFX9 U631 ( .A(n2894), .Z(n284) );
  HS65_LH_NAND2X7 U632 ( .A(n840), .B(n841), .Z(n346) );
  HS65_LH_NAND2X7 U633 ( .A(n1368), .B(n1369), .Z(n874) );
  HS65_LH_NAND2X7 U634 ( .A(n842), .B(n845), .Z(n350) );
  HS65_LH_NAND2X7 U635 ( .A(n840), .B(n845), .Z(n351) );
  HS65_LH_NAND2X7 U636 ( .A(n1370), .B(n1373), .Z(n878) );
  HS65_LH_NAND2X7 U637 ( .A(n1368), .B(n1373), .Z(n879) );
  HS65_LH_NAND2X7 U638 ( .A(n843), .B(n857), .Z(n367) );
  HS65_LH_NAND2X7 U639 ( .A(n843), .B(n856), .Z(n368) );
  HS65_LH_NAND2X7 U640 ( .A(n1371), .B(n1385), .Z(n895) );
  HS65_LH_NAND2X7 U641 ( .A(n1371), .B(n1384), .Z(n896) );
  HS65_LH_NAND2X7 U642 ( .A(n846), .B(n856), .Z(n373) );
  HS65_LH_NAND2X7 U643 ( .A(n1374), .B(n1385), .Z(n900) );
  HS65_LH_NAND2X7 U644 ( .A(n1374), .B(n1384), .Z(n901) );
  HS65_LH_AND2X4 U645 ( .A(n847), .B(n2898), .Z(n842) );
  HS65_LH_AND2X4 U646 ( .A(n1375), .B(n2903), .Z(n1370) );
  HS65_LH_AND2X4 U647 ( .A(n1387), .B(n2903), .Z(n1385) );
  HS65_LH_BFX9 U648 ( .A(n2893), .Z(n281) );
  HS65_LH_BFX9 U649 ( .A(n2894), .Z(n287) );
  HS65_LH_BFX9 U650 ( .A(n2894), .Z(n286) );
  HS65_LH_BFX9 U651 ( .A(n2893), .Z(n282) );
  HS65_LH_NAND2X7 U652 ( .A(n1408), .B(n1391), .Z(n1407) );
  HS65_LH_NAND2X7 U653 ( .A(n1408), .B(n1393), .Z(n1409) );
  HS65_LH_NAND2X7 U654 ( .A(n1408), .B(n1404), .Z(n1414) );
  HS65_LH_NAND2X7 U655 ( .A(n1408), .B(n1406), .Z(n1415) );
  HS65_LH_NAND2X7 U656 ( .A(n1426), .B(n1402), .Z(n1431) );
  HS65_LH_NAND2X7 U657 ( .A(n1417), .B(n1391), .Z(n1416) );
  HS65_LH_NAND2X7 U658 ( .A(n1426), .B(n1391), .Z(n1425) );
  HS65_LH_NAND2X7 U659 ( .A(n1426), .B(n1400), .Z(n1430) );
  HS65_LH_NAND2X7 U660 ( .A(n1426), .B(n1396), .Z(n1428) );
  HS65_LH_NAND2X7 U661 ( .A(n1426), .B(n1398), .Z(n1429) );
  HS65_LH_IVX9 U662 ( .A(\regfile_i[FORWARD_B] ), .Z(n2894) );
  HS65_LH_NOR2X6 U663 ( .A(n2900), .B(\regfile_i[ADRREAD1][1] ), .Z(n843) );
  HS65_LH_NOR2X6 U664 ( .A(n2905), .B(\regfile_i[ADRREAD0][1] ), .Z(n1371) );
  HS65_LH_NOR2X6 U665 ( .A(n2899), .B(\regfile_i[ADRREAD1][2] ), .Z(n846) );
  HS65_LH_NOR2X6 U666 ( .A(n2904), .B(\regfile_i[ADRREAD0][2] ), .Z(n1374) );
  HS65_LH_NOR2X6 U667 ( .A(\regfile_i[ADRREAD1][1] ), .B(
        \regfile_i[ADRREAD1][2] ), .Z(n845) );
  HS65_LH_NOR2X6 U668 ( .A(\regfile_i[ADRREAD0][1] ), .B(
        \regfile_i[ADRREAD0][2] ), .Z(n1373) );
  HS65_LH_AOI212X4 U669 ( .A(\registers[11][0] ), .B(n2682), .C(
        \registers[10][0] ), .D(n2679), .E(n844), .Z(n837) );
  HS65_LH_OAI22X6 U670 ( .A(n2676), .B(n256), .C(n2673), .D(n224), .Z(n844) );
  HS65_LH_AOI212X4 U671 ( .A(\registers[11][1] ), .B(n2682), .C(
        \registers[10][1] ), .D(n2679), .E(n675), .Z(n672) );
  HS65_LH_OAI22X6 U672 ( .A(n2676), .B(n255), .C(n2673), .D(n223), .Z(n675) );
  HS65_LH_AOI212X4 U673 ( .A(\registers[11][2] ), .B(n2683), .C(
        \registers[10][2] ), .D(n2680), .E(n510), .Z(n507) );
  HS65_LH_OAI22X6 U674 ( .A(n2677), .B(n254), .C(n2674), .D(n222), .Z(n510) );
  HS65_LH_AOI212X4 U675 ( .A(\registers[11][11] ), .B(n2682), .C(
        \registers[10][11] ), .D(n2679), .E(n810), .Z(n807) );
  HS65_LH_OAI22X6 U676 ( .A(n2676), .B(n245), .C(n2673), .D(n213), .Z(n810) );
  HS65_LH_AOI212X4 U677 ( .A(\registers[11][12] ), .B(n2682), .C(
        \registers[10][12] ), .D(n2679), .E(n795), .Z(n792) );
  HS65_LH_OAI22X6 U678 ( .A(n2676), .B(n244), .C(n2673), .D(n212), .Z(n795) );
  HS65_LH_AOI212X4 U679 ( .A(\registers[11][13] ), .B(n2682), .C(
        \registers[10][13] ), .D(n2679), .E(n780), .Z(n777) );
  HS65_LH_OAI22X6 U680 ( .A(n2676), .B(n243), .C(n2673), .D(n211), .Z(n780) );
  HS65_LH_AOI212X4 U681 ( .A(\registers[11][14] ), .B(n2682), .C(
        \registers[10][14] ), .D(n2679), .E(n765), .Z(n762) );
  HS65_LH_OAI22X6 U682 ( .A(n2676), .B(n242), .C(n2673), .D(n210), .Z(n765) );
  HS65_LH_AOI212X4 U683 ( .A(\registers[11][15] ), .B(n2682), .C(
        \registers[10][15] ), .D(n2679), .E(n750), .Z(n747) );
  HS65_LH_OAI22X6 U684 ( .A(n2676), .B(n241), .C(n2673), .D(n209), .Z(n750) );
  HS65_LH_AOI212X4 U685 ( .A(\registers[11][16] ), .B(n2682), .C(
        \registers[10][16] ), .D(n2679), .E(n735), .Z(n732) );
  HS65_LH_OAI22X6 U686 ( .A(n2676), .B(n240), .C(n2673), .D(n208), .Z(n735) );
  HS65_LH_AOI212X4 U687 ( .A(\registers[11][17] ), .B(n2682), .C(
        \registers[10][17] ), .D(n2679), .E(n720), .Z(n717) );
  HS65_LH_OAI22X6 U688 ( .A(n2676), .B(n239), .C(n2673), .D(n207), .Z(n720) );
  HS65_LH_AOI212X4 U689 ( .A(\registers[11][18] ), .B(n2682), .C(
        \registers[10][18] ), .D(n2679), .E(n705), .Z(n702) );
  HS65_LH_OAI22X6 U690 ( .A(n2676), .B(n238), .C(n2673), .D(n206), .Z(n705) );
  HS65_LH_AOI212X4 U691 ( .A(\registers[11][19] ), .B(n2682), .C(
        \registers[10][19] ), .D(n2679), .E(n690), .Z(n687) );
  HS65_LH_OAI22X6 U692 ( .A(n2676), .B(n237), .C(n2673), .D(n205), .Z(n690) );
  HS65_LH_AOI212X4 U693 ( .A(\registers[11][20] ), .B(n2683), .C(
        \registers[10][20] ), .D(n2679), .E(n660), .Z(n657) );
  HS65_LH_OAI22X6 U694 ( .A(n2677), .B(n236), .C(n2673), .D(n204), .Z(n660) );
  HS65_LH_AOI212X4 U695 ( .A(\registers[11][21] ), .B(n2683), .C(
        \registers[10][21] ), .D(n2680), .E(n645), .Z(n642) );
  HS65_LH_OAI22X6 U696 ( .A(n2677), .B(n235), .C(n2674), .D(n203), .Z(n645) );
  HS65_LH_AOI212X4 U697 ( .A(\registers[11][22] ), .B(n2683), .C(
        \registers[10][22] ), .D(n2680), .E(n630), .Z(n627) );
  HS65_LH_OAI22X6 U698 ( .A(n2677), .B(n234), .C(n2674), .D(n202), .Z(n630) );
  HS65_LH_AOI212X4 U699 ( .A(\registers[11][23] ), .B(n2683), .C(
        \registers[10][23] ), .D(n2680), .E(n615), .Z(n612) );
  HS65_LH_OAI22X6 U700 ( .A(n2677), .B(n233), .C(n2674), .D(n201), .Z(n615) );
  HS65_LH_AOI212X4 U701 ( .A(\registers[11][24] ), .B(n2683), .C(
        \registers[10][24] ), .D(n2680), .E(n600), .Z(n597) );
  HS65_LH_OAI22X6 U702 ( .A(n2677), .B(n232), .C(n2674), .D(n200), .Z(n600) );
  HS65_LH_AOI212X4 U703 ( .A(\registers[11][25] ), .B(n2683), .C(
        \registers[10][25] ), .D(n2680), .E(n585), .Z(n582) );
  HS65_LH_OAI22X6 U704 ( .A(n2677), .B(n231), .C(n2674), .D(n199), .Z(n585) );
  HS65_LH_AOI212X4 U705 ( .A(\registers[11][26] ), .B(n2683), .C(
        \registers[10][26] ), .D(n2680), .E(n570), .Z(n567) );
  HS65_LH_OAI22X6 U706 ( .A(n2677), .B(n230), .C(n2674), .D(n198), .Z(n570) );
  HS65_LH_AOI212X4 U707 ( .A(\registers[11][27] ), .B(n2683), .C(
        \registers[10][27] ), .D(n2680), .E(n555), .Z(n552) );
  HS65_LH_OAI22X6 U708 ( .A(n2677), .B(n229), .C(n2674), .D(n197), .Z(n555) );
  HS65_LH_AOI212X4 U709 ( .A(\registers[11][28] ), .B(n2683), .C(
        \registers[10][28] ), .D(n2680), .E(n540), .Z(n537) );
  HS65_LH_OAI22X6 U710 ( .A(n2677), .B(n228), .C(n2674), .D(n196), .Z(n540) );
  HS65_LH_AOI212X4 U711 ( .A(\registers[11][29] ), .B(n2683), .C(
        \registers[10][29] ), .D(n2680), .E(n525), .Z(n522) );
  HS65_LH_OAI22X6 U712 ( .A(n2677), .B(n227), .C(n2674), .D(n195), .Z(n525) );
  HS65_LH_AOI212X4 U713 ( .A(\registers[11][30] ), .B(n2683), .C(
        \registers[10][30] ), .D(n2680), .E(n495), .Z(n492) );
  HS65_LH_OAI22X6 U714 ( .A(n2677), .B(n226), .C(n2674), .D(n194), .Z(n495) );
  HS65_LH_AOI212X4 U715 ( .A(n2589), .B(\registers[11][0] ), .C(n2586), .D(
        \registers[10][0] ), .E(n1372), .Z(n1365) );
  HS65_LH_OAI22X6 U716 ( .A(n256), .B(n2583), .C(n224), .D(n2580), .Z(n1372)
         );
  HS65_LH_AOI212X4 U717 ( .A(n2589), .B(\registers[11][1] ), .C(n2586), .D(
        \registers[10][1] ), .E(n1203), .Z(n1200) );
  HS65_LH_OAI22X6 U718 ( .A(n255), .B(n2583), .C(n223), .D(n2580), .Z(n1203)
         );
  HS65_LH_AOI212X4 U719 ( .A(n2590), .B(\registers[11][2] ), .C(n2587), .D(
        \registers[10][2] ), .E(n1038), .Z(n1035) );
  HS65_LH_OAI22X6 U720 ( .A(n254), .B(n2584), .C(n222), .D(n2581), .Z(n1038)
         );
  HS65_LH_AOI212X4 U721 ( .A(n2590), .B(\registers[11][3] ), .C(n2587), .D(
        \registers[10][3] ), .E(n993), .Z(n990) );
  HS65_LH_OAI22X6 U722 ( .A(n253), .B(n2585), .C(n221), .D(n2581), .Z(n993) );
  HS65_LH_AOI212X4 U723 ( .A(n2591), .B(\registers[11][4] ), .C(n2588), .D(
        \registers[10][4] ), .E(n978), .Z(n975) );
  HS65_LH_OAI22X6 U724 ( .A(n252), .B(n2585), .C(n220), .D(n2582), .Z(n978) );
  HS65_LH_AOI212X4 U725 ( .A(n2591), .B(\registers[11][5] ), .C(n2588), .D(
        \registers[10][5] ), .E(n963), .Z(n960) );
  HS65_LH_OAI22X6 U726 ( .A(n251), .B(n2585), .C(n219), .D(n2582), .Z(n963) );
  HS65_LH_AOI212X4 U727 ( .A(n2591), .B(\registers[11][6] ), .C(n2588), .D(
        \registers[10][6] ), .E(n948), .Z(n945) );
  HS65_LH_OAI22X6 U728 ( .A(n250), .B(n2585), .C(n218), .D(n2582), .Z(n948) );
  HS65_LH_AOI212X4 U729 ( .A(n2591), .B(\registers[11][7] ), .C(n2588), .D(
        \registers[10][7] ), .E(n933), .Z(n930) );
  HS65_LH_OAI22X6 U730 ( .A(n249), .B(n2585), .C(n217), .D(n2582), .Z(n933) );
  HS65_LH_AOI212X4 U731 ( .A(n2591), .B(\registers[11][8] ), .C(n2588), .D(
        \registers[10][8] ), .E(n918), .Z(n915) );
  HS65_LH_OAI22X6 U732 ( .A(n248), .B(n2585), .C(n216), .D(n2582), .Z(n918) );
  HS65_LH_AOI212X4 U733 ( .A(n2591), .B(\registers[11][9] ), .C(n2588), .D(
        \registers[10][9] ), .E(n877), .Z(n868) );
  HS65_LH_OAI22X6 U734 ( .A(n247), .B(n2585), .C(n215), .D(n2582), .Z(n877) );
  HS65_LH_AOI212X4 U735 ( .A(n2589), .B(\registers[11][10] ), .C(n2586), .D(
        \registers[10][10] ), .E(n1353), .Z(n1350) );
  HS65_LH_OAI22X6 U736 ( .A(n246), .B(n2583), .C(n214), .D(n2580), .Z(n1353)
         );
  HS65_LH_AOI212X4 U737 ( .A(n2589), .B(\registers[11][11] ), .C(n2586), .D(
        \registers[10][11] ), .E(n1338), .Z(n1335) );
  HS65_LH_OAI22X6 U738 ( .A(n245), .B(n2583), .C(n213), .D(n2580), .Z(n1338)
         );
  HS65_LH_AOI212X4 U739 ( .A(n2589), .B(\registers[11][12] ), .C(n2586), .D(
        \registers[10][12] ), .E(n1323), .Z(n1320) );
  HS65_LH_OAI22X6 U740 ( .A(n244), .B(n2583), .C(n212), .D(n2580), .Z(n1323)
         );
  HS65_LH_AOI212X4 U741 ( .A(n2589), .B(\registers[11][13] ), .C(n2586), .D(
        \registers[10][13] ), .E(n1308), .Z(n1305) );
  HS65_LH_OAI22X6 U742 ( .A(n243), .B(n2583), .C(n211), .D(n2580), .Z(n1308)
         );
  HS65_LH_AOI212X4 U743 ( .A(n2589), .B(\registers[11][14] ), .C(n2586), .D(
        \registers[10][14] ), .E(n1293), .Z(n1290) );
  HS65_LH_OAI22X6 U744 ( .A(n242), .B(n2583), .C(n210), .D(n2580), .Z(n1293)
         );
  HS65_LH_AOI212X4 U745 ( .A(n2589), .B(\registers[11][15] ), .C(n2586), .D(
        \registers[10][15] ), .E(n1278), .Z(n1275) );
  HS65_LH_OAI22X6 U746 ( .A(n241), .B(n2583), .C(n209), .D(n2580), .Z(n1278)
         );
  HS65_LH_AOI212X4 U747 ( .A(n2589), .B(\registers[11][16] ), .C(n2586), .D(
        \registers[10][16] ), .E(n1263), .Z(n1260) );
  HS65_LH_OAI22X6 U748 ( .A(n240), .B(n2583), .C(n208), .D(n2580), .Z(n1263)
         );
  HS65_LH_AOI212X4 U749 ( .A(n2589), .B(\registers[11][17] ), .C(n2586), .D(
        \registers[10][17] ), .E(n1248), .Z(n1245) );
  HS65_LH_OAI22X6 U750 ( .A(n239), .B(n2583), .C(n207), .D(n2580), .Z(n1248)
         );
  HS65_LH_AOI212X4 U751 ( .A(n2589), .B(\registers[11][18] ), .C(n2586), .D(
        \registers[10][18] ), .E(n1233), .Z(n1230) );
  HS65_LH_OAI22X6 U752 ( .A(n238), .B(n2583), .C(n206), .D(n2580), .Z(n1233)
         );
  HS65_LH_AOI212X4 U753 ( .A(n2589), .B(\registers[11][19] ), .C(n2586), .D(
        \registers[10][19] ), .E(n1218), .Z(n1215) );
  HS65_LH_OAI22X6 U754 ( .A(n237), .B(n2583), .C(n205), .D(n2580), .Z(n1218)
         );
  HS65_LH_AOI212X4 U755 ( .A(n2589), .B(\registers[11][20] ), .C(n2586), .D(
        \registers[10][20] ), .E(n1188), .Z(n1185) );
  HS65_LH_OAI22X6 U756 ( .A(n236), .B(n2584), .C(n204), .D(n2580), .Z(n1188)
         );
  HS65_LH_AOI212X4 U757 ( .A(n2590), .B(\registers[11][21] ), .C(n2587), .D(
        \registers[10][21] ), .E(n1173), .Z(n1170) );
  HS65_LH_OAI22X6 U758 ( .A(n235), .B(n2584), .C(n203), .D(n2581), .Z(n1173)
         );
  HS65_LH_AOI212X4 U759 ( .A(n2590), .B(\registers[11][22] ), .C(n2587), .D(
        \registers[10][22] ), .E(n1158), .Z(n1155) );
  HS65_LH_OAI22X6 U760 ( .A(n234), .B(n2584), .C(n202), .D(n2581), .Z(n1158)
         );
  HS65_LH_AOI212X4 U761 ( .A(n2590), .B(\registers[11][23] ), .C(n2587), .D(
        \registers[10][23] ), .E(n1143), .Z(n1140) );
  HS65_LH_OAI22X6 U762 ( .A(n233), .B(n2584), .C(n201), .D(n2581), .Z(n1143)
         );
  HS65_LH_AOI212X4 U763 ( .A(n2590), .B(\registers[11][24] ), .C(n2587), .D(
        \registers[10][24] ), .E(n1128), .Z(n1125) );
  HS65_LH_OAI22X6 U764 ( .A(n232), .B(n2584), .C(n200), .D(n2581), .Z(n1128)
         );
  HS65_LH_AOI212X4 U765 ( .A(n2590), .B(\registers[11][25] ), .C(n2587), .D(
        \registers[10][25] ), .E(n1113), .Z(n1110) );
  HS65_LH_OAI22X6 U766 ( .A(n231), .B(n2584), .C(n199), .D(n2581), .Z(n1113)
         );
  HS65_LH_AOI212X4 U767 ( .A(n2590), .B(\registers[11][26] ), .C(n2587), .D(
        \registers[10][26] ), .E(n1098), .Z(n1095) );
  HS65_LH_OAI22X6 U768 ( .A(n230), .B(n2584), .C(n198), .D(n2581), .Z(n1098)
         );
  HS65_LH_AOI212X4 U769 ( .A(n2590), .B(\registers[11][27] ), .C(n2587), .D(
        \registers[10][27] ), .E(n1083), .Z(n1080) );
  HS65_LH_OAI22X6 U770 ( .A(n229), .B(n2584), .C(n197), .D(n2581), .Z(n1083)
         );
  HS65_LH_AOI212X4 U771 ( .A(n2590), .B(\registers[11][28] ), .C(n2587), .D(
        \registers[10][28] ), .E(n1068), .Z(n1065) );
  HS65_LH_OAI22X6 U772 ( .A(n228), .B(n2584), .C(n196), .D(n2581), .Z(n1068)
         );
  HS65_LH_AOI212X4 U773 ( .A(n2590), .B(\registers[11][29] ), .C(n2587), .D(
        \registers[10][29] ), .E(n1053), .Z(n1050) );
  HS65_LH_OAI22X6 U774 ( .A(n227), .B(n2584), .C(n195), .D(n2581), .Z(n1053)
         );
  HS65_LH_AOI212X4 U775 ( .A(n2590), .B(\registers[11][30] ), .C(n2587), .D(
        \registers[10][30] ), .E(n1023), .Z(n1020) );
  HS65_LH_OAI22X6 U776 ( .A(n226), .B(n2584), .C(n194), .D(n2581), .Z(n1023)
         );
  HS65_LH_AOI212X4 U777 ( .A(n2590), .B(\registers[11][31] ), .C(n2587), .D(
        \registers[10][31] ), .E(n1008), .Z(n1005) );
  HS65_LH_OAI22X6 U778 ( .A(n225), .B(n2585), .C(n193), .D(n2581), .Z(n1008)
         );
  HS65_LH_AOI212X4 U779 ( .A(n2601), .B(\registers[13][0] ), .C(n2598), .D(
        \registers[12][0] ), .E(n1367), .Z(n1366) );
  HS65_LH_OAI22X6 U780 ( .A(n192), .B(n2595), .C(n160), .D(n2592), .Z(n1367)
         );
  HS65_LH_AOI212X4 U781 ( .A(n2601), .B(\registers[13][1] ), .C(n2598), .D(
        \registers[12][1] ), .E(n1202), .Z(n1201) );
  HS65_LH_OAI22X6 U782 ( .A(n191), .B(n2595), .C(n159), .D(n2592), .Z(n1202)
         );
  HS65_LH_AOI212X4 U783 ( .A(n2602), .B(\registers[13][2] ), .C(n2599), .D(
        \registers[12][2] ), .E(n1037), .Z(n1036) );
  HS65_LH_OAI22X6 U784 ( .A(n190), .B(n2596), .C(n158), .D(n2593), .Z(n1037)
         );
  HS65_LH_AOI212X4 U785 ( .A(n2602), .B(\registers[13][3] ), .C(n2599), .D(
        \registers[12][3] ), .E(n992), .Z(n991) );
  HS65_LH_OAI22X6 U786 ( .A(n189), .B(n2597), .C(n157), .D(n2593), .Z(n992) );
  HS65_LH_AOI212X4 U787 ( .A(n2601), .B(\registers[13][10] ), .C(n2598), .D(
        \registers[12][10] ), .E(n1352), .Z(n1351) );
  HS65_LH_OAI22X6 U788 ( .A(n182), .B(n2595), .C(n150), .D(n2592), .Z(n1352)
         );
  HS65_LH_AOI212X4 U789 ( .A(n2601), .B(\registers[13][11] ), .C(n2598), .D(
        \registers[12][11] ), .E(n1337), .Z(n1336) );
  HS65_LH_OAI22X6 U790 ( .A(n181), .B(n2595), .C(n149), .D(n2592), .Z(n1337)
         );
  HS65_LH_AOI212X4 U791 ( .A(n2601), .B(\registers[13][12] ), .C(n2598), .D(
        \registers[12][12] ), .E(n1322), .Z(n1321) );
  HS65_LH_OAI22X6 U792 ( .A(n180), .B(n2595), .C(n148), .D(n2592), .Z(n1322)
         );
  HS65_LH_AOI212X4 U793 ( .A(n2601), .B(\registers[13][13] ), .C(n2598), .D(
        \registers[12][13] ), .E(n1307), .Z(n1306) );
  HS65_LH_OAI22X6 U794 ( .A(n179), .B(n2595), .C(n147), .D(n2592), .Z(n1307)
         );
  HS65_LH_AOI212X4 U795 ( .A(n2601), .B(\registers[13][14] ), .C(n2598), .D(
        \registers[12][14] ), .E(n1292), .Z(n1291) );
  HS65_LH_OAI22X6 U796 ( .A(n178), .B(n2595), .C(n146), .D(n2592), .Z(n1292)
         );
  HS65_LH_AOI212X4 U797 ( .A(n2601), .B(\registers[13][15] ), .C(n2598), .D(
        \registers[12][15] ), .E(n1277), .Z(n1276) );
  HS65_LH_OAI22X6 U798 ( .A(n177), .B(n2595), .C(n145), .D(n2592), .Z(n1277)
         );
  HS65_LH_AOI212X4 U799 ( .A(n2601), .B(\registers[13][16] ), .C(n2598), .D(
        \registers[12][16] ), .E(n1262), .Z(n1261) );
  HS65_LH_OAI22X6 U800 ( .A(n176), .B(n2595), .C(n144), .D(n2592), .Z(n1262)
         );
  HS65_LH_AOI212X4 U801 ( .A(n2601), .B(\registers[13][17] ), .C(n2598), .D(
        \registers[12][17] ), .E(n1247), .Z(n1246) );
  HS65_LH_OAI22X6 U802 ( .A(n175), .B(n2595), .C(n143), .D(n2592), .Z(n1247)
         );
  HS65_LH_AOI212X4 U803 ( .A(n2601), .B(\registers[13][18] ), .C(n2598), .D(
        \registers[12][18] ), .E(n1232), .Z(n1231) );
  HS65_LH_OAI22X6 U804 ( .A(n174), .B(n2595), .C(n142), .D(n2592), .Z(n1232)
         );
  HS65_LH_AOI212X4 U805 ( .A(n2601), .B(\registers[13][19] ), .C(n2598), .D(
        \registers[12][19] ), .E(n1217), .Z(n1216) );
  HS65_LH_OAI22X6 U806 ( .A(n173), .B(n2595), .C(n141), .D(n2592), .Z(n1217)
         );
  HS65_LH_AOI212X4 U807 ( .A(n2601), .B(\registers[13][20] ), .C(n2598), .D(
        \registers[12][20] ), .E(n1187), .Z(n1186) );
  HS65_LH_OAI22X6 U808 ( .A(n172), .B(n2596), .C(n140), .D(n2592), .Z(n1187)
         );
  HS65_LH_AOI212X4 U809 ( .A(n2602), .B(\registers[13][21] ), .C(n2599), .D(
        \registers[12][21] ), .E(n1172), .Z(n1171) );
  HS65_LH_OAI22X6 U810 ( .A(n171), .B(n2596), .C(n139), .D(n2593), .Z(n1172)
         );
  HS65_LH_AOI212X4 U811 ( .A(n2602), .B(\registers[13][22] ), .C(n2599), .D(
        \registers[12][22] ), .E(n1157), .Z(n1156) );
  HS65_LH_OAI22X6 U812 ( .A(n170), .B(n2596), .C(n138), .D(n2593), .Z(n1157)
         );
  HS65_LH_AOI212X4 U813 ( .A(n2602), .B(\registers[13][23] ), .C(n2599), .D(
        \registers[12][23] ), .E(n1142), .Z(n1141) );
  HS65_LH_OAI22X6 U814 ( .A(n169), .B(n2596), .C(n137), .D(n2593), .Z(n1142)
         );
  HS65_LH_AOI212X4 U815 ( .A(n2602), .B(\registers[13][24] ), .C(n2599), .D(
        \registers[12][24] ), .E(n1127), .Z(n1126) );
  HS65_LH_OAI22X6 U816 ( .A(n168), .B(n2596), .C(n136), .D(n2593), .Z(n1127)
         );
  HS65_LH_AOI212X4 U817 ( .A(n2602), .B(\registers[13][25] ), .C(n2599), .D(
        \registers[12][25] ), .E(n1112), .Z(n1111) );
  HS65_LH_OAI22X6 U818 ( .A(n167), .B(n2596), .C(n135), .D(n2593), .Z(n1112)
         );
  HS65_LH_AOI212X4 U819 ( .A(n2602), .B(\registers[13][26] ), .C(n2599), .D(
        \registers[12][26] ), .E(n1097), .Z(n1096) );
  HS65_LH_OAI22X6 U820 ( .A(n166), .B(n2596), .C(n134), .D(n2593), .Z(n1097)
         );
  HS65_LH_AOI212X4 U821 ( .A(n2602), .B(\registers[13][27] ), .C(n2599), .D(
        \registers[12][27] ), .E(n1082), .Z(n1081) );
  HS65_LH_OAI22X6 U822 ( .A(n165), .B(n2596), .C(n133), .D(n2593), .Z(n1082)
         );
  HS65_LH_AOI212X4 U823 ( .A(n2602), .B(\registers[13][28] ), .C(n2599), .D(
        \registers[12][28] ), .E(n1067), .Z(n1066) );
  HS65_LH_OAI22X6 U824 ( .A(n164), .B(n2596), .C(n132), .D(n2593), .Z(n1067)
         );
  HS65_LH_AOI212X4 U825 ( .A(n2602), .B(\registers[13][29] ), .C(n2599), .D(
        \registers[12][29] ), .E(n1052), .Z(n1051) );
  HS65_LH_OAI22X6 U826 ( .A(n163), .B(n2596), .C(n131), .D(n2593), .Z(n1052)
         );
  HS65_LH_AOI212X4 U827 ( .A(n2602), .B(\registers[13][30] ), .C(n2599), .D(
        \registers[12][30] ), .E(n1022), .Z(n1021) );
  HS65_LH_OAI22X6 U828 ( .A(n162), .B(n2596), .C(n130), .D(n2593), .Z(n1022)
         );
  HS65_LH_AOI212X4 U829 ( .A(n2602), .B(\registers[13][31] ), .C(n2599), .D(
        \registers[12][31] ), .E(n1007), .Z(n1006) );
  HS65_LH_OAI22X6 U830 ( .A(n161), .B(n2597), .C(n129), .D(n2593), .Z(n1007)
         );
  HS65_LH_OAI22X6 U831 ( .A(n2631), .B(n128), .C(n2628), .D(n96), .Z(n858) );
  HS65_LH_OAI22X6 U832 ( .A(n2631), .B(n127), .C(n2628), .D(n95), .Z(n681) );
  HS65_LH_OAI22X6 U833 ( .A(n2632), .B(n126), .C(n2629), .D(n94), .Z(n516) );
  HS65_LH_OAI22X6 U834 ( .A(n2631), .B(n118), .C(n2628), .D(n86), .Z(n831) );
  HS65_LH_OAI22X6 U835 ( .A(n2631), .B(n117), .C(n2628), .D(n85), .Z(n816) );
  HS65_LH_OAI22X6 U836 ( .A(n2631), .B(n116), .C(n2628), .D(n84), .Z(n801) );
  HS65_LH_OAI22X6 U837 ( .A(n2631), .B(n115), .C(n2628), .D(n83), .Z(n786) );
  HS65_LH_OAI22X6 U838 ( .A(n2631), .B(n114), .C(n2628), .D(n82), .Z(n771) );
  HS65_LH_OAI22X6 U839 ( .A(n2631), .B(n113), .C(n2628), .D(n81), .Z(n756) );
  HS65_LH_OAI22X6 U840 ( .A(n2631), .B(n112), .C(n2628), .D(n80), .Z(n741) );
  HS65_LH_OAI22X6 U841 ( .A(n2631), .B(n111), .C(n2628), .D(n79), .Z(n726) );
  HS65_LH_OAI22X6 U842 ( .A(n2631), .B(n110), .C(n2628), .D(n78), .Z(n711) );
  HS65_LH_OAI22X6 U843 ( .A(n2631), .B(n109), .C(n2628), .D(n77), .Z(n696) );
  HS65_LH_OAI22X6 U844 ( .A(n2632), .B(n108), .C(n2628), .D(n76), .Z(n666) );
  HS65_LH_OAI22X6 U845 ( .A(n2632), .B(n107), .C(n2629), .D(n75), .Z(n651) );
  HS65_LH_OAI22X6 U846 ( .A(n2632), .B(n106), .C(n2629), .D(n74), .Z(n636) );
  HS65_LH_OAI22X6 U847 ( .A(n2632), .B(n105), .C(n2629), .D(n73), .Z(n621) );
  HS65_LH_OAI22X6 U848 ( .A(n2632), .B(n104), .C(n2629), .D(n72), .Z(n606) );
  HS65_LH_OAI22X6 U849 ( .A(n2632), .B(n103), .C(n2629), .D(n71), .Z(n591) );
  HS65_LH_OAI22X6 U850 ( .A(n2632), .B(n102), .C(n2629), .D(n70), .Z(n576) );
  HS65_LH_OAI22X6 U851 ( .A(n2632), .B(n101), .C(n2629), .D(n69), .Z(n561) );
  HS65_LH_OAI22X6 U852 ( .A(n2632), .B(n100), .C(n2629), .D(n68), .Z(n546) );
  HS65_LH_OAI22X6 U853 ( .A(n2632), .B(n99), .C(n2629), .D(n67), .Z(n531) );
  HS65_LH_OAI22X6 U854 ( .A(n2632), .B(n98), .C(n2629), .D(n66), .Z(n501) );
  HS65_LH_NAND4ABX3 U855 ( .A(n851), .B(n852), .C(n853), .D(n854), .Z(n833) );
  HS65_LH_AOI212X4 U856 ( .A(\registers[31][0] ), .B(n2649), .C(
        \registers[30][0] ), .D(n2646), .E(n855), .Z(n854) );
  HS65_LH_AOI212X4 U857 ( .A(\registers[25][0] ), .B(n2637), .C(
        \registers[24][0] ), .D(n2634), .E(n858), .Z(n853) );
  HS65_LH_MX41X7 U858 ( .D0(\registers[16][0] ), .S0(n2625), .D1(
        \registers[17][0] ), .S1(n2622), .D2(\registers[18][0] ), .S2(n2619), 
        .D3(\registers[19][0] ), .S3(n2616), .Z(n852) );
  HS65_LH_NAND4ABX3 U859 ( .A(n676), .B(n677), .C(n678), .D(n679), .Z(n668) );
  HS65_LH_AOI212X4 U860 ( .A(\registers[31][1] ), .B(n2649), .C(
        \registers[30][1] ), .D(n2646), .E(n680), .Z(n679) );
  HS65_LH_AOI212X4 U861 ( .A(\registers[25][1] ), .B(n2637), .C(
        \registers[24][1] ), .D(n2634), .E(n681), .Z(n678) );
  HS65_LH_MX41X7 U862 ( .D0(\registers[16][1] ), .S0(n2625), .D1(
        \registers[17][1] ), .S1(n2622), .D2(\registers[18][1] ), .S2(n2619), 
        .D3(\registers[19][1] ), .S3(n2616), .Z(n677) );
  HS65_LH_NAND4ABX3 U863 ( .A(n511), .B(n512), .C(n513), .D(n514), .Z(n503) );
  HS65_LH_AOI212X4 U864 ( .A(\registers[31][2] ), .B(n2650), .C(
        \registers[30][2] ), .D(n2647), .E(n515), .Z(n514) );
  HS65_LH_AOI212X4 U865 ( .A(\registers[25][2] ), .B(n2638), .C(
        \registers[24][2] ), .D(n2635), .E(n516), .Z(n513) );
  HS65_LH_MX41X7 U866 ( .D0(\registers[16][2] ), .S0(n2626), .D1(
        \registers[17][2] ), .S1(n2623), .D2(\registers[18][2] ), .S2(n2620), 
        .D3(\registers[19][2] ), .S3(n2617), .Z(n512) );
  HS65_LH_NAND4ABX3 U867 ( .A(n466), .B(n467), .C(n468), .D(n469), .Z(n458) );
  HS65_LH_AOI212X4 U868 ( .A(\registers[31][3] ), .B(n2651), .C(
        \registers[30][3] ), .D(n2647), .E(n470), .Z(n469) );
  HS65_LH_AOI212X4 U869 ( .A(\registers[25][3] ), .B(n2639), .C(
        \registers[24][3] ), .D(n2635), .E(n471), .Z(n468) );
  HS65_LH_MX41X7 U870 ( .D0(\registers[16][3] ), .S0(n2627), .D1(
        \registers[17][3] ), .S1(n2624), .D2(\registers[18][3] ), .S2(n2621), 
        .D3(\registers[19][3] ), .S3(n2618), .Z(n467) );
  HS65_LH_NAND4ABX3 U871 ( .A(n451), .B(n452), .C(n453), .D(n454), .Z(n443) );
  HS65_LH_AOI212X4 U872 ( .A(\registers[31][4] ), .B(n2651), .C(
        \registers[30][4] ), .D(n2648), .E(n455), .Z(n454) );
  HS65_LH_AOI212X4 U873 ( .A(\registers[25][4] ), .B(n2639), .C(
        \registers[24][4] ), .D(n2636), .E(n456), .Z(n453) );
  HS65_LH_MX41X7 U874 ( .D0(\registers[16][4] ), .S0(n2627), .D1(
        \registers[17][4] ), .S1(n2624), .D2(\registers[18][4] ), .S2(n2621), 
        .D3(\registers[19][4] ), .S3(n2618), .Z(n452) );
  HS65_LH_NAND4ABX3 U875 ( .A(n436), .B(n437), .C(n438), .D(n439), .Z(n428) );
  HS65_LH_AOI212X4 U876 ( .A(\registers[31][5] ), .B(n2651), .C(
        \registers[30][5] ), .D(n2648), .E(n440), .Z(n439) );
  HS65_LH_AOI212X4 U877 ( .A(\registers[25][5] ), .B(n2639), .C(
        \registers[24][5] ), .D(n2636), .E(n441), .Z(n438) );
  HS65_LH_MX41X7 U878 ( .D0(\registers[16][5] ), .S0(n2627), .D1(
        \registers[17][5] ), .S1(n2624), .D2(\registers[18][5] ), .S2(n2621), 
        .D3(\registers[19][5] ), .S3(n2618), .Z(n437) );
  HS65_LH_NAND4ABX3 U879 ( .A(n421), .B(n422), .C(n423), .D(n424), .Z(n413) );
  HS65_LH_AOI212X4 U880 ( .A(\registers[31][6] ), .B(n2651), .C(
        \registers[30][6] ), .D(n2648), .E(n425), .Z(n424) );
  HS65_LH_AOI212X4 U881 ( .A(\registers[25][6] ), .B(n2639), .C(
        \registers[24][6] ), .D(n2636), .E(n426), .Z(n423) );
  HS65_LH_MX41X7 U882 ( .D0(\registers[16][6] ), .S0(n2627), .D1(
        \registers[17][6] ), .S1(n2624), .D2(\registers[18][6] ), .S2(n2621), 
        .D3(\registers[19][6] ), .S3(n2618), .Z(n422) );
  HS65_LH_NAND4ABX3 U883 ( .A(n406), .B(n407), .C(n408), .D(n409), .Z(n398) );
  HS65_LH_AOI212X4 U884 ( .A(\registers[31][7] ), .B(n2651), .C(
        \registers[30][7] ), .D(n2648), .E(n410), .Z(n409) );
  HS65_LH_AOI212X4 U885 ( .A(\registers[25][7] ), .B(n2639), .C(
        \registers[24][7] ), .D(n2636), .E(n411), .Z(n408) );
  HS65_LH_MX41X7 U886 ( .D0(\registers[16][7] ), .S0(n2627), .D1(
        \registers[17][7] ), .S1(n2624), .D2(\registers[18][7] ), .S2(n2621), 
        .D3(\registers[19][7] ), .S3(n2618), .Z(n407) );
  HS65_LH_NAND4ABX3 U887 ( .A(n391), .B(n392), .C(n393), .D(n394), .Z(n383) );
  HS65_LH_AOI212X4 U888 ( .A(\registers[31][8] ), .B(n2651), .C(
        \registers[30][8] ), .D(n2648), .E(n395), .Z(n394) );
  HS65_LH_AOI212X4 U889 ( .A(\registers[25][8] ), .B(n2639), .C(
        \registers[24][8] ), .D(n2636), .E(n396), .Z(n393) );
  HS65_LH_MX41X7 U890 ( .D0(\registers[16][8] ), .S0(n2627), .D1(
        \registers[17][8] ), .S1(n2624), .D2(\registers[18][8] ), .S2(n2621), 
        .D3(\registers[19][8] ), .S3(n2618), .Z(n392) );
  HS65_LH_NAND4ABX3 U891 ( .A(n360), .B(n361), .C(n362), .D(n363), .Z(n336) );
  HS65_LH_AOI212X4 U892 ( .A(\registers[31][9] ), .B(n2651), .C(
        \registers[30][9] ), .D(n2648), .E(n366), .Z(n363) );
  HS65_LH_AOI212X4 U893 ( .A(\registers[25][9] ), .B(n2639), .C(
        \registers[24][9] ), .D(n2636), .E(n371), .Z(n362) );
  HS65_LH_MX41X7 U894 ( .D0(\registers[16][9] ), .S0(n2627), .D1(
        \registers[17][9] ), .S1(n2624), .D2(\registers[18][9] ), .S2(n2621), 
        .D3(\registers[19][9] ), .S3(n2618), .Z(n361) );
  HS65_LH_NAND4ABX3 U895 ( .A(n826), .B(n827), .C(n828), .D(n829), .Z(n818) );
  HS65_LH_AOI212X4 U896 ( .A(\registers[31][10] ), .B(n2649), .C(
        \registers[30][10] ), .D(n2646), .E(n830), .Z(n829) );
  HS65_LH_AOI212X4 U897 ( .A(\registers[25][10] ), .B(n2637), .C(
        \registers[24][10] ), .D(n2634), .E(n831), .Z(n828) );
  HS65_LH_MX41X7 U898 ( .D0(\registers[16][10] ), .S0(n2625), .D1(
        \registers[17][10] ), .S1(n2622), .D2(\registers[18][10] ), .S2(n2619), 
        .D3(\registers[19][10] ), .S3(n2616), .Z(n827) );
  HS65_LH_NAND4ABX3 U899 ( .A(n811), .B(n812), .C(n813), .D(n814), .Z(n803) );
  HS65_LH_AOI212X4 U900 ( .A(\registers[31][11] ), .B(n2649), .C(
        \registers[30][11] ), .D(n2646), .E(n815), .Z(n814) );
  HS65_LH_AOI212X4 U901 ( .A(\registers[25][11] ), .B(n2637), .C(
        \registers[24][11] ), .D(n2634), .E(n816), .Z(n813) );
  HS65_LH_MX41X7 U902 ( .D0(\registers[16][11] ), .S0(n2625), .D1(
        \registers[17][11] ), .S1(n2622), .D2(\registers[18][11] ), .S2(n2619), 
        .D3(\registers[19][11] ), .S3(n2616), .Z(n812) );
  HS65_LH_NAND4ABX3 U903 ( .A(n796), .B(n797), .C(n798), .D(n799), .Z(n788) );
  HS65_LH_AOI212X4 U904 ( .A(\registers[31][12] ), .B(n2649), .C(
        \registers[30][12] ), .D(n2646), .E(n800), .Z(n799) );
  HS65_LH_AOI212X4 U905 ( .A(\registers[25][12] ), .B(n2637), .C(
        \registers[24][12] ), .D(n2634), .E(n801), .Z(n798) );
  HS65_LH_MX41X7 U906 ( .D0(\registers[16][12] ), .S0(n2625), .D1(
        \registers[17][12] ), .S1(n2622), .D2(\registers[18][12] ), .S2(n2619), 
        .D3(\registers[19][12] ), .S3(n2616), .Z(n797) );
  HS65_LH_NAND4ABX3 U907 ( .A(n781), .B(n782), .C(n783), .D(n784), .Z(n773) );
  HS65_LH_AOI212X4 U908 ( .A(\registers[31][13] ), .B(n2649), .C(
        \registers[30][13] ), .D(n2646), .E(n785), .Z(n784) );
  HS65_LH_AOI212X4 U909 ( .A(\registers[25][13] ), .B(n2637), .C(
        \registers[24][13] ), .D(n2634), .E(n786), .Z(n783) );
  HS65_LH_MX41X7 U910 ( .D0(\registers[16][13] ), .S0(n2625), .D1(
        \registers[17][13] ), .S1(n2622), .D2(\registers[18][13] ), .S2(n2619), 
        .D3(\registers[19][13] ), .S3(n2616), .Z(n782) );
  HS65_LH_NAND4ABX3 U911 ( .A(n766), .B(n767), .C(n768), .D(n769), .Z(n758) );
  HS65_LH_AOI212X4 U912 ( .A(\registers[31][14] ), .B(n2649), .C(
        \registers[30][14] ), .D(n2646), .E(n770), .Z(n769) );
  HS65_LH_AOI212X4 U913 ( .A(\registers[25][14] ), .B(n2637), .C(
        \registers[24][14] ), .D(n2634), .E(n771), .Z(n768) );
  HS65_LH_MX41X7 U914 ( .D0(\registers[16][14] ), .S0(n2625), .D1(
        \registers[17][14] ), .S1(n2622), .D2(\registers[18][14] ), .S2(n2619), 
        .D3(\registers[19][14] ), .S3(n2616), .Z(n767) );
  HS65_LH_NAND4ABX3 U915 ( .A(n751), .B(n752), .C(n753), .D(n754), .Z(n743) );
  HS65_LH_AOI212X4 U916 ( .A(\registers[31][15] ), .B(n2649), .C(
        \registers[30][15] ), .D(n2646), .E(n755), .Z(n754) );
  HS65_LH_AOI212X4 U917 ( .A(\registers[25][15] ), .B(n2637), .C(
        \registers[24][15] ), .D(n2634), .E(n756), .Z(n753) );
  HS65_LH_MX41X7 U918 ( .D0(\registers[16][15] ), .S0(n2625), .D1(
        \registers[17][15] ), .S1(n2622), .D2(\registers[18][15] ), .S2(n2619), 
        .D3(\registers[19][15] ), .S3(n2616), .Z(n752) );
  HS65_LH_NAND4ABX3 U919 ( .A(n736), .B(n737), .C(n738), .D(n739), .Z(n728) );
  HS65_LH_AOI212X4 U920 ( .A(\registers[31][16] ), .B(n2649), .C(
        \registers[30][16] ), .D(n2646), .E(n740), .Z(n739) );
  HS65_LH_AOI212X4 U921 ( .A(\registers[25][16] ), .B(n2637), .C(
        \registers[24][16] ), .D(n2634), .E(n741), .Z(n738) );
  HS65_LH_MX41X7 U922 ( .D0(\registers[16][16] ), .S0(n2625), .D1(
        \registers[17][16] ), .S1(n2622), .D2(\registers[18][16] ), .S2(n2619), 
        .D3(\registers[19][16] ), .S3(n2616), .Z(n737) );
  HS65_LH_NAND4ABX3 U923 ( .A(n721), .B(n722), .C(n723), .D(n724), .Z(n713) );
  HS65_LH_AOI212X4 U924 ( .A(\registers[31][17] ), .B(n2649), .C(
        \registers[30][17] ), .D(n2646), .E(n725), .Z(n724) );
  HS65_LH_AOI212X4 U925 ( .A(\registers[25][17] ), .B(n2637), .C(
        \registers[24][17] ), .D(n2634), .E(n726), .Z(n723) );
  HS65_LH_MX41X7 U926 ( .D0(\registers[16][17] ), .S0(n2625), .D1(
        \registers[17][17] ), .S1(n2622), .D2(\registers[18][17] ), .S2(n2619), 
        .D3(\registers[19][17] ), .S3(n2616), .Z(n722) );
  HS65_LH_NAND4ABX3 U927 ( .A(n706), .B(n707), .C(n708), .D(n709), .Z(n698) );
  HS65_LH_AOI212X4 U928 ( .A(\registers[31][18] ), .B(n2649), .C(
        \registers[30][18] ), .D(n2646), .E(n710), .Z(n709) );
  HS65_LH_AOI212X4 U929 ( .A(\registers[25][18] ), .B(n2637), .C(
        \registers[24][18] ), .D(n2634), .E(n711), .Z(n708) );
  HS65_LH_MX41X7 U930 ( .D0(\registers[16][18] ), .S0(n2625), .D1(
        \registers[17][18] ), .S1(n2622), .D2(\registers[18][18] ), .S2(n2619), 
        .D3(\registers[19][18] ), .S3(n2616), .Z(n707) );
  HS65_LH_NAND4ABX3 U931 ( .A(n691), .B(n692), .C(n693), .D(n694), .Z(n683) );
  HS65_LH_AOI212X4 U932 ( .A(\registers[31][19] ), .B(n2649), .C(
        \registers[30][19] ), .D(n2646), .E(n695), .Z(n694) );
  HS65_LH_AOI212X4 U933 ( .A(\registers[25][19] ), .B(n2637), .C(
        \registers[24][19] ), .D(n2634), .E(n696), .Z(n693) );
  HS65_LH_MX41X7 U934 ( .D0(\registers[16][19] ), .S0(n2625), .D1(
        \registers[17][19] ), .S1(n2622), .D2(\registers[18][19] ), .S2(n2619), 
        .D3(\registers[19][19] ), .S3(n2616), .Z(n692) );
  HS65_LH_NAND4ABX3 U935 ( .A(n661), .B(n662), .C(n663), .D(n664), .Z(n653) );
  HS65_LH_AOI212X4 U936 ( .A(\registers[31][20] ), .B(n2650), .C(
        \registers[30][20] ), .D(n2646), .E(n665), .Z(n664) );
  HS65_LH_AOI212X4 U937 ( .A(\registers[25][20] ), .B(n2638), .C(
        \registers[24][20] ), .D(n2634), .E(n666), .Z(n663) );
  HS65_LH_MX41X7 U938 ( .D0(\registers[16][20] ), .S0(n2626), .D1(
        \registers[17][20] ), .S1(n2623), .D2(\registers[18][20] ), .S2(n2620), 
        .D3(\registers[19][20] ), .S3(n2617), .Z(n662) );
  HS65_LH_NAND4ABX3 U939 ( .A(n646), .B(n647), .C(n648), .D(n649), .Z(n638) );
  HS65_LH_AOI212X4 U940 ( .A(\registers[31][21] ), .B(n2650), .C(
        \registers[30][21] ), .D(n2647), .E(n650), .Z(n649) );
  HS65_LH_AOI212X4 U941 ( .A(\registers[25][21] ), .B(n2638), .C(
        \registers[24][21] ), .D(n2635), .E(n651), .Z(n648) );
  HS65_LH_MX41X7 U942 ( .D0(\registers[16][21] ), .S0(n2626), .D1(
        \registers[17][21] ), .S1(n2623), .D2(\registers[18][21] ), .S2(n2620), 
        .D3(\registers[19][21] ), .S3(n2617), .Z(n647) );
  HS65_LH_NAND4ABX3 U943 ( .A(n631), .B(n632), .C(n633), .D(n634), .Z(n623) );
  HS65_LH_AOI212X4 U944 ( .A(\registers[31][22] ), .B(n2650), .C(
        \registers[30][22] ), .D(n2647), .E(n635), .Z(n634) );
  HS65_LH_AOI212X4 U945 ( .A(\registers[25][22] ), .B(n2638), .C(
        \registers[24][22] ), .D(n2635), .E(n636), .Z(n633) );
  HS65_LH_MX41X7 U946 ( .D0(\registers[16][22] ), .S0(n2626), .D1(
        \registers[17][22] ), .S1(n2623), .D2(\registers[18][22] ), .S2(n2620), 
        .D3(\registers[19][22] ), .S3(n2617), .Z(n632) );
  HS65_LH_NAND4ABX3 U947 ( .A(n616), .B(n617), .C(n618), .D(n619), .Z(n608) );
  HS65_LH_AOI212X4 U948 ( .A(\registers[31][23] ), .B(n2650), .C(
        \registers[30][23] ), .D(n2647), .E(n620), .Z(n619) );
  HS65_LH_AOI212X4 U949 ( .A(\registers[25][23] ), .B(n2638), .C(
        \registers[24][23] ), .D(n2635), .E(n621), .Z(n618) );
  HS65_LH_MX41X7 U950 ( .D0(\registers[16][23] ), .S0(n2626), .D1(
        \registers[17][23] ), .S1(n2623), .D2(\registers[18][23] ), .S2(n2620), 
        .D3(\registers[19][23] ), .S3(n2617), .Z(n617) );
  HS65_LH_NAND4ABX3 U951 ( .A(n601), .B(n602), .C(n603), .D(n604), .Z(n593) );
  HS65_LH_AOI212X4 U952 ( .A(\registers[31][24] ), .B(n2650), .C(
        \registers[30][24] ), .D(n2647), .E(n605), .Z(n604) );
  HS65_LH_AOI212X4 U953 ( .A(\registers[25][24] ), .B(n2638), .C(
        \registers[24][24] ), .D(n2635), .E(n606), .Z(n603) );
  HS65_LH_MX41X7 U954 ( .D0(\registers[16][24] ), .S0(n2626), .D1(
        \registers[17][24] ), .S1(n2623), .D2(\registers[18][24] ), .S2(n2620), 
        .D3(\registers[19][24] ), .S3(n2617), .Z(n602) );
  HS65_LH_NAND4ABX3 U955 ( .A(n586), .B(n587), .C(n588), .D(n589), .Z(n578) );
  HS65_LH_AOI212X4 U956 ( .A(\registers[31][25] ), .B(n2650), .C(
        \registers[30][25] ), .D(n2647), .E(n590), .Z(n589) );
  HS65_LH_AOI212X4 U957 ( .A(\registers[25][25] ), .B(n2638), .C(
        \registers[24][25] ), .D(n2635), .E(n591), .Z(n588) );
  HS65_LH_MX41X7 U958 ( .D0(\registers[16][25] ), .S0(n2626), .D1(
        \registers[17][25] ), .S1(n2623), .D2(\registers[18][25] ), .S2(n2620), 
        .D3(\registers[19][25] ), .S3(n2617), .Z(n587) );
  HS65_LH_NAND4ABX3 U959 ( .A(n571), .B(n572), .C(n573), .D(n574), .Z(n563) );
  HS65_LH_AOI212X4 U960 ( .A(\registers[31][26] ), .B(n2650), .C(
        \registers[30][26] ), .D(n2647), .E(n575), .Z(n574) );
  HS65_LH_AOI212X4 U961 ( .A(\registers[25][26] ), .B(n2638), .C(
        \registers[24][26] ), .D(n2635), .E(n576), .Z(n573) );
  HS65_LH_MX41X7 U962 ( .D0(\registers[16][26] ), .S0(n2626), .D1(
        \registers[17][26] ), .S1(n2623), .D2(\registers[18][26] ), .S2(n2620), 
        .D3(\registers[19][26] ), .S3(n2617), .Z(n572) );
  HS65_LH_NAND4ABX3 U963 ( .A(n556), .B(n557), .C(n558), .D(n559), .Z(n548) );
  HS65_LH_AOI212X4 U964 ( .A(\registers[31][27] ), .B(n2650), .C(
        \registers[30][27] ), .D(n2647), .E(n560), .Z(n559) );
  HS65_LH_AOI212X4 U965 ( .A(\registers[25][27] ), .B(n2638), .C(
        \registers[24][27] ), .D(n2635), .E(n561), .Z(n558) );
  HS65_LH_MX41X7 U966 ( .D0(\registers[16][27] ), .S0(n2626), .D1(
        \registers[17][27] ), .S1(n2623), .D2(\registers[18][27] ), .S2(n2620), 
        .D3(\registers[19][27] ), .S3(n2617), .Z(n557) );
  HS65_LH_NAND4ABX3 U967 ( .A(n541), .B(n542), .C(n543), .D(n544), .Z(n533) );
  HS65_LH_AOI212X4 U968 ( .A(\registers[31][28] ), .B(n2650), .C(
        \registers[30][28] ), .D(n2647), .E(n545), .Z(n544) );
  HS65_LH_AOI212X4 U969 ( .A(\registers[25][28] ), .B(n2638), .C(
        \registers[24][28] ), .D(n2635), .E(n546), .Z(n543) );
  HS65_LH_MX41X7 U970 ( .D0(\registers[16][28] ), .S0(n2626), .D1(
        \registers[17][28] ), .S1(n2623), .D2(\registers[18][28] ), .S2(n2620), 
        .D3(\registers[19][28] ), .S3(n2617), .Z(n542) );
  HS65_LH_NAND4ABX3 U971 ( .A(n526), .B(n527), .C(n528), .D(n529), .Z(n518) );
  HS65_LH_AOI212X4 U972 ( .A(\registers[31][29] ), .B(n2650), .C(
        \registers[30][29] ), .D(n2647), .E(n530), .Z(n529) );
  HS65_LH_AOI212X4 U973 ( .A(\registers[25][29] ), .B(n2638), .C(
        \registers[24][29] ), .D(n2635), .E(n531), .Z(n528) );
  HS65_LH_MX41X7 U974 ( .D0(\registers[16][29] ), .S0(n2626), .D1(
        \registers[17][29] ), .S1(n2623), .D2(\registers[18][29] ), .S2(n2620), 
        .D3(\registers[19][29] ), .S3(n2617), .Z(n527) );
  HS65_LH_NAND4ABX3 U975 ( .A(n496), .B(n497), .C(n498), .D(n499), .Z(n488) );
  HS65_LH_AOI212X4 U976 ( .A(\registers[31][30] ), .B(n2650), .C(
        \registers[30][30] ), .D(n2647), .E(n500), .Z(n499) );
  HS65_LH_AOI212X4 U977 ( .A(\registers[25][30] ), .B(n2638), .C(
        \registers[24][30] ), .D(n2635), .E(n501), .Z(n498) );
  HS65_LH_MX41X7 U978 ( .D0(\registers[16][30] ), .S0(n2626), .D1(
        \registers[17][30] ), .S1(n2623), .D2(\registers[18][30] ), .S2(n2620), 
        .D3(\registers[19][30] ), .S3(n2617), .Z(n497) );
  HS65_LH_NAND4ABX3 U979 ( .A(n481), .B(n482), .C(n483), .D(n484), .Z(n473) );
  HS65_LH_AOI212X4 U980 ( .A(\registers[31][31] ), .B(n2651), .C(
        \registers[30][31] ), .D(n2647), .E(n485), .Z(n484) );
  HS65_LH_AOI212X4 U981 ( .A(\registers[25][31] ), .B(n2639), .C(
        \registers[24][31] ), .D(n2635), .E(n486), .Z(n483) );
  HS65_LH_MX41X7 U982 ( .D0(\registers[16][31] ), .S0(n2627), .D1(
        \registers[17][31] ), .S1(n2624), .D2(\registers[18][31] ), .S2(n2621), 
        .D3(\registers[19][31] ), .S3(n2618), .Z(n482) );
  HS65_LH_NAND4ABX3 U983 ( .A(n1379), .B(n1380), .C(n1381), .D(n1382), .Z(
        n1361) );
  HS65_LH_AOI212X4 U984 ( .A(n2556), .B(\registers[31][0] ), .C(n2553), .D(
        \registers[30][0] ), .E(n1383), .Z(n1382) );
  HS65_LH_AOI212X4 U985 ( .A(n2544), .B(\registers[25][0] ), .C(n2541), .D(
        \registers[24][0] ), .E(n1386), .Z(n1381) );
  HS65_LH_MX41X7 U986 ( .D0(n2532), .S0(\registers[16][0] ), .D1(n2529), .S1(
        \registers[17][0] ), .D2(n2526), .S2(\registers[18][0] ), .D3(n2523), 
        .S3(\registers[19][0] ), .Z(n1380) );
  HS65_LH_NAND4ABX3 U987 ( .A(n1204), .B(n1205), .C(n1206), .D(n1207), .Z(
        n1196) );
  HS65_LH_AOI212X4 U988 ( .A(n2556), .B(\registers[31][1] ), .C(n2553), .D(
        \registers[30][1] ), .E(n1208), .Z(n1207) );
  HS65_LH_AOI212X4 U989 ( .A(n2544), .B(\registers[25][1] ), .C(n2541), .D(
        \registers[24][1] ), .E(n1209), .Z(n1206) );
  HS65_LH_MX41X7 U990 ( .D0(n2532), .S0(\registers[16][1] ), .D1(n2529), .S1(
        \registers[17][1] ), .D2(n2526), .S2(\registers[18][1] ), .D3(n2523), 
        .S3(\registers[19][1] ), .Z(n1205) );
  HS65_LH_NAND4ABX3 U991 ( .A(n1039), .B(n1040), .C(n1041), .D(n1042), .Z(
        n1031) );
  HS65_LH_AOI212X4 U992 ( .A(n2557), .B(\registers[31][2] ), .C(n2554), .D(
        \registers[30][2] ), .E(n1043), .Z(n1042) );
  HS65_LH_AOI212X4 U993 ( .A(n2545), .B(\registers[25][2] ), .C(n2542), .D(
        \registers[24][2] ), .E(n1044), .Z(n1041) );
  HS65_LH_MX41X7 U994 ( .D0(n2533), .S0(\registers[16][2] ), .D1(n2530), .S1(
        \registers[17][2] ), .D2(n2527), .S2(\registers[18][2] ), .D3(n2524), 
        .S3(\registers[19][2] ), .Z(n1040) );
  HS65_LH_NAND4ABX3 U995 ( .A(n994), .B(n995), .C(n996), .D(n997), .Z(n986) );
  HS65_LH_AOI212X4 U996 ( .A(n2557), .B(\registers[31][3] ), .C(n2554), .D(
        \registers[30][3] ), .E(n998), .Z(n997) );
  HS65_LH_AOI212X4 U997 ( .A(n2545), .B(\registers[25][3] ), .C(n2542), .D(
        \registers[24][3] ), .E(n999), .Z(n996) );
  HS65_LH_MX41X7 U998 ( .D0(n2533), .S0(\registers[16][3] ), .D1(n2531), .S1(
        \registers[17][3] ), .D2(n2527), .S2(\registers[18][3] ), .D3(n2525), 
        .S3(\registers[19][3] ), .Z(n995) );
  HS65_LH_NAND4ABX3 U999 ( .A(n979), .B(n980), .C(n981), .D(n982), .Z(n971) );
  HS65_LH_AOI212X4 U1000 ( .A(n2558), .B(\registers[31][4] ), .C(n2555), .D(
        \registers[30][4] ), .E(n983), .Z(n982) );
  HS65_LH_AOI212X4 U1001 ( .A(n2546), .B(\registers[25][4] ), .C(n2543), .D(
        \registers[24][4] ), .E(n984), .Z(n981) );
  HS65_LH_MX41X7 U1002 ( .D0(n2534), .S0(\registers[16][4] ), .D1(n2531), .S1(
        \registers[17][4] ), .D2(n2528), .S2(\registers[18][4] ), .D3(n2525), 
        .S3(\registers[19][4] ), .Z(n980) );
  HS65_LH_NAND4ABX3 U1003 ( .A(n964), .B(n965), .C(n966), .D(n967), .Z(n956)
         );
  HS65_LH_AOI212X4 U1004 ( .A(n2558), .B(\registers[31][5] ), .C(n2555), .D(
        \registers[30][5] ), .E(n968), .Z(n967) );
  HS65_LH_AOI212X4 U1005 ( .A(n2546), .B(\registers[25][5] ), .C(n2543), .D(
        \registers[24][5] ), .E(n969), .Z(n966) );
  HS65_LH_MX41X7 U1006 ( .D0(n2534), .S0(\registers[16][5] ), .D1(n2531), .S1(
        \registers[17][5] ), .D2(n2528), .S2(\registers[18][5] ), .D3(n2525), 
        .S3(\registers[19][5] ), .Z(n965) );
  HS65_LH_NAND4ABX3 U1007 ( .A(n949), .B(n950), .C(n951), .D(n952), .Z(n941)
         );
  HS65_LH_AOI212X4 U1008 ( .A(n2558), .B(\registers[31][6] ), .C(n2555), .D(
        \registers[30][6] ), .E(n953), .Z(n952) );
  HS65_LH_AOI212X4 U1009 ( .A(n2546), .B(\registers[25][6] ), .C(n2543), .D(
        \registers[24][6] ), .E(n954), .Z(n951) );
  HS65_LH_MX41X7 U1010 ( .D0(n2534), .S0(\registers[16][6] ), .D1(n2531), .S1(
        \registers[17][6] ), .D2(n2528), .S2(\registers[18][6] ), .D3(n2525), 
        .S3(\registers[19][6] ), .Z(n950) );
  HS65_LH_NAND4ABX3 U1011 ( .A(n934), .B(n935), .C(n936), .D(n937), .Z(n926)
         );
  HS65_LH_AOI212X4 U1012 ( .A(n2558), .B(\registers[31][7] ), .C(n2555), .D(
        \registers[30][7] ), .E(n938), .Z(n937) );
  HS65_LH_AOI212X4 U1013 ( .A(n2546), .B(\registers[25][7] ), .C(n2543), .D(
        \registers[24][7] ), .E(n939), .Z(n936) );
  HS65_LH_MX41X7 U1014 ( .D0(n2534), .S0(\registers[16][7] ), .D1(n2531), .S1(
        \registers[17][7] ), .D2(n2528), .S2(\registers[18][7] ), .D3(n2525), 
        .S3(\registers[19][7] ), .Z(n935) );
  HS65_LH_NAND4ABX3 U1015 ( .A(n919), .B(n920), .C(n921), .D(n922), .Z(n911)
         );
  HS65_LH_AOI212X4 U1016 ( .A(n2558), .B(\registers[31][8] ), .C(n2555), .D(
        \registers[30][8] ), .E(n923), .Z(n922) );
  HS65_LH_AOI212X4 U1017 ( .A(n2546), .B(\registers[25][8] ), .C(n2543), .D(
        \registers[24][8] ), .E(n924), .Z(n921) );
  HS65_LH_MX41X7 U1018 ( .D0(n2534), .S0(\registers[16][8] ), .D1(n2531), .S1(
        \registers[17][8] ), .D2(n2528), .S2(\registers[18][8] ), .D3(n2525), 
        .S3(\registers[19][8] ), .Z(n920) );
  HS65_LH_NAND4ABX3 U1019 ( .A(n888), .B(n889), .C(n890), .D(n891), .Z(n864)
         );
  HS65_LH_AOI212X4 U1020 ( .A(n2558), .B(\registers[31][9] ), .C(n2555), .D(
        \registers[30][9] ), .E(n894), .Z(n891) );
  HS65_LH_AOI212X4 U1021 ( .A(n2546), .B(\registers[25][9] ), .C(n2543), .D(
        \registers[24][9] ), .E(n899), .Z(n890) );
  HS65_LH_MX41X7 U1022 ( .D0(n2534), .S0(\registers[16][9] ), .D1(n2531), .S1(
        \registers[17][9] ), .D2(n2528), .S2(\registers[18][9] ), .D3(n2525), 
        .S3(\registers[19][9] ), .Z(n889) );
  HS65_LH_NAND4ABX3 U1023 ( .A(n1354), .B(n1355), .C(n1356), .D(n1357), .Z(
        n1346) );
  HS65_LH_AOI212X4 U1024 ( .A(n2556), .B(\registers[31][10] ), .C(n2553), .D(
        \registers[30][10] ), .E(n1358), .Z(n1357) );
  HS65_LH_AOI212X4 U1025 ( .A(n2544), .B(\registers[25][10] ), .C(n2541), .D(
        \registers[24][10] ), .E(n1359), .Z(n1356) );
  HS65_LH_MX41X7 U1026 ( .D0(n2532), .S0(\registers[16][10] ), .D1(n2529), 
        .S1(\registers[17][10] ), .D2(n2526), .S2(\registers[18][10] ), .D3(
        n2523), .S3(\registers[19][10] ), .Z(n1355) );
  HS65_LH_NAND4ABX3 U1027 ( .A(n1339), .B(n1340), .C(n1341), .D(n1342), .Z(
        n1331) );
  HS65_LH_AOI212X4 U1028 ( .A(n2556), .B(\registers[31][11] ), .C(n2553), .D(
        \registers[30][11] ), .E(n1343), .Z(n1342) );
  HS65_LH_AOI212X4 U1029 ( .A(n2544), .B(\registers[25][11] ), .C(n2541), .D(
        \registers[24][11] ), .E(n1344), .Z(n1341) );
  HS65_LH_MX41X7 U1030 ( .D0(n2532), .S0(\registers[16][11] ), .D1(n2529), 
        .S1(\registers[17][11] ), .D2(n2526), .S2(\registers[18][11] ), .D3(
        n2523), .S3(\registers[19][11] ), .Z(n1340) );
  HS65_LH_NAND4ABX3 U1031 ( .A(n1324), .B(n1325), .C(n1326), .D(n1327), .Z(
        n1316) );
  HS65_LH_AOI212X4 U1032 ( .A(n2556), .B(\registers[31][12] ), .C(n2553), .D(
        \registers[30][12] ), .E(n1328), .Z(n1327) );
  HS65_LH_AOI212X4 U1033 ( .A(n2544), .B(\registers[25][12] ), .C(n2541), .D(
        \registers[24][12] ), .E(n1329), .Z(n1326) );
  HS65_LH_MX41X7 U1034 ( .D0(n2532), .S0(\registers[16][12] ), .D1(n2529), 
        .S1(\registers[17][12] ), .D2(n2526), .S2(\registers[18][12] ), .D3(
        n2523), .S3(\registers[19][12] ), .Z(n1325) );
  HS65_LH_NAND4ABX3 U1035 ( .A(n1309), .B(n1310), .C(n1311), .D(n1312), .Z(
        n1301) );
  HS65_LH_AOI212X4 U1036 ( .A(n2556), .B(\registers[31][13] ), .C(n2553), .D(
        \registers[30][13] ), .E(n1313), .Z(n1312) );
  HS65_LH_AOI212X4 U1037 ( .A(n2544), .B(\registers[25][13] ), .C(n2541), .D(
        \registers[24][13] ), .E(n1314), .Z(n1311) );
  HS65_LH_MX41X7 U1038 ( .D0(n2532), .S0(\registers[16][13] ), .D1(n2529), 
        .S1(\registers[17][13] ), .D2(n2526), .S2(\registers[18][13] ), .D3(
        n2523), .S3(\registers[19][13] ), .Z(n1310) );
  HS65_LH_NAND4ABX3 U1039 ( .A(n1294), .B(n1295), .C(n1296), .D(n1297), .Z(
        n1286) );
  HS65_LH_AOI212X4 U1040 ( .A(n2556), .B(\registers[31][14] ), .C(n2553), .D(
        \registers[30][14] ), .E(n1298), .Z(n1297) );
  HS65_LH_AOI212X4 U1041 ( .A(n2544), .B(\registers[25][14] ), .C(n2541), .D(
        \registers[24][14] ), .E(n1299), .Z(n1296) );
  HS65_LH_MX41X7 U1042 ( .D0(n2532), .S0(\registers[16][14] ), .D1(n2529), 
        .S1(\registers[17][14] ), .D2(n2526), .S2(\registers[18][14] ), .D3(
        n2523), .S3(\registers[19][14] ), .Z(n1295) );
  HS65_LH_NAND4ABX3 U1043 ( .A(n1279), .B(n1280), .C(n1281), .D(n1282), .Z(
        n1271) );
  HS65_LH_AOI212X4 U1044 ( .A(n2556), .B(\registers[31][15] ), .C(n2553), .D(
        \registers[30][15] ), .E(n1283), .Z(n1282) );
  HS65_LH_AOI212X4 U1045 ( .A(n2544), .B(\registers[25][15] ), .C(n2541), .D(
        \registers[24][15] ), .E(n1284), .Z(n1281) );
  HS65_LH_MX41X7 U1046 ( .D0(n2532), .S0(\registers[16][15] ), .D1(n2529), 
        .S1(\registers[17][15] ), .D2(n2526), .S2(\registers[18][15] ), .D3(
        n2523), .S3(\registers[19][15] ), .Z(n1280) );
  HS65_LH_NAND4ABX3 U1047 ( .A(n1264), .B(n1265), .C(n1266), .D(n1267), .Z(
        n1256) );
  HS65_LH_AOI212X4 U1048 ( .A(n2556), .B(\registers[31][16] ), .C(n2553), .D(
        \registers[30][16] ), .E(n1268), .Z(n1267) );
  HS65_LH_AOI212X4 U1049 ( .A(n2544), .B(\registers[25][16] ), .C(n2541), .D(
        \registers[24][16] ), .E(n1269), .Z(n1266) );
  HS65_LH_MX41X7 U1050 ( .D0(n2532), .S0(\registers[16][16] ), .D1(n2529), 
        .S1(\registers[17][16] ), .D2(n2526), .S2(\registers[18][16] ), .D3(
        n2523), .S3(\registers[19][16] ), .Z(n1265) );
  HS65_LH_NAND4ABX3 U1051 ( .A(n1249), .B(n1250), .C(n1251), .D(n1252), .Z(
        n1241) );
  HS65_LH_AOI212X4 U1052 ( .A(n2556), .B(\registers[31][17] ), .C(n2553), .D(
        \registers[30][17] ), .E(n1253), .Z(n1252) );
  HS65_LH_AOI212X4 U1053 ( .A(n2544), .B(\registers[25][17] ), .C(n2541), .D(
        \registers[24][17] ), .E(n1254), .Z(n1251) );
  HS65_LH_MX41X7 U1054 ( .D0(n2532), .S0(\registers[16][17] ), .D1(n2529), 
        .S1(\registers[17][17] ), .D2(n2526), .S2(\registers[18][17] ), .D3(
        n2523), .S3(\registers[19][17] ), .Z(n1250) );
  HS65_LH_NAND4ABX3 U1055 ( .A(n1234), .B(n1235), .C(n1236), .D(n1237), .Z(
        n1226) );
  HS65_LH_AOI212X4 U1056 ( .A(n2556), .B(\registers[31][18] ), .C(n2553), .D(
        \registers[30][18] ), .E(n1238), .Z(n1237) );
  HS65_LH_AOI212X4 U1057 ( .A(n2544), .B(\registers[25][18] ), .C(n2541), .D(
        \registers[24][18] ), .E(n1239), .Z(n1236) );
  HS65_LH_MX41X7 U1058 ( .D0(n2532), .S0(\registers[16][18] ), .D1(n2529), 
        .S1(\registers[17][18] ), .D2(n2526), .S2(\registers[18][18] ), .D3(
        n2523), .S3(\registers[19][18] ), .Z(n1235) );
  HS65_LH_NAND4ABX3 U1059 ( .A(n1219), .B(n1220), .C(n1221), .D(n1222), .Z(
        n1211) );
  HS65_LH_AOI212X4 U1060 ( .A(n2556), .B(\registers[31][19] ), .C(n2553), .D(
        \registers[30][19] ), .E(n1223), .Z(n1222) );
  HS65_LH_AOI212X4 U1061 ( .A(n2544), .B(\registers[25][19] ), .C(n2541), .D(
        \registers[24][19] ), .E(n1224), .Z(n1221) );
  HS65_LH_MX41X7 U1062 ( .D0(n2532), .S0(\registers[16][19] ), .D1(n2529), 
        .S1(\registers[17][19] ), .D2(n2526), .S2(\registers[18][19] ), .D3(
        n2523), .S3(\registers[19][19] ), .Z(n1220) );
  HS65_LH_NAND4ABX3 U1063 ( .A(n1189), .B(n1190), .C(n1191), .D(n1192), .Z(
        n1181) );
  HS65_LH_AOI212X4 U1064 ( .A(n2556), .B(\registers[31][20] ), .C(n2553), .D(
        \registers[30][20] ), .E(n1193), .Z(n1192) );
  HS65_LH_AOI212X4 U1065 ( .A(n2544), .B(\registers[25][20] ), .C(n2541), .D(
        \registers[24][20] ), .E(n1194), .Z(n1191) );
  HS65_LH_MX41X7 U1066 ( .D0(n2532), .S0(\registers[16][20] ), .D1(n2530), 
        .S1(\registers[17][20] ), .D2(n2526), .S2(\registers[18][20] ), .D3(
        n2524), .S3(\registers[19][20] ), .Z(n1190) );
  HS65_LH_NAND4ABX3 U1067 ( .A(n1174), .B(n1175), .C(n1176), .D(n1177), .Z(
        n1166) );
  HS65_LH_AOI212X4 U1068 ( .A(n2557), .B(\registers[31][21] ), .C(n2554), .D(
        \registers[30][21] ), .E(n1178), .Z(n1177) );
  HS65_LH_AOI212X4 U1069 ( .A(n2545), .B(\registers[25][21] ), .C(n2542), .D(
        \registers[24][21] ), .E(n1179), .Z(n1176) );
  HS65_LH_MX41X7 U1070 ( .D0(n2533), .S0(\registers[16][21] ), .D1(n2530), 
        .S1(\registers[17][21] ), .D2(n2527), .S2(\registers[18][21] ), .D3(
        n2524), .S3(\registers[19][21] ), .Z(n1175) );
  HS65_LH_NAND4ABX3 U1071 ( .A(n1159), .B(n1160), .C(n1161), .D(n1162), .Z(
        n1151) );
  HS65_LH_AOI212X4 U1072 ( .A(n2557), .B(\registers[31][22] ), .C(n2554), .D(
        \registers[30][22] ), .E(n1163), .Z(n1162) );
  HS65_LH_AOI212X4 U1073 ( .A(n2545), .B(\registers[25][22] ), .C(n2542), .D(
        \registers[24][22] ), .E(n1164), .Z(n1161) );
  HS65_LH_MX41X7 U1074 ( .D0(n2533), .S0(\registers[16][22] ), .D1(n2530), 
        .S1(\registers[17][22] ), .D2(n2527), .S2(\registers[18][22] ), .D3(
        n2524), .S3(\registers[19][22] ), .Z(n1160) );
  HS65_LH_NAND4ABX3 U1075 ( .A(n1144), .B(n1145), .C(n1146), .D(n1147), .Z(
        n1136) );
  HS65_LH_AOI212X4 U1076 ( .A(n2557), .B(\registers[31][23] ), .C(n2554), .D(
        \registers[30][23] ), .E(n1148), .Z(n1147) );
  HS65_LH_AOI212X4 U1077 ( .A(n2545), .B(\registers[25][23] ), .C(n2542), .D(
        \registers[24][23] ), .E(n1149), .Z(n1146) );
  HS65_LH_MX41X7 U1078 ( .D0(n2533), .S0(\registers[16][23] ), .D1(n2530), 
        .S1(\registers[17][23] ), .D2(n2527), .S2(\registers[18][23] ), .D3(
        n2524), .S3(\registers[19][23] ), .Z(n1145) );
  HS65_LH_NAND4ABX3 U1079 ( .A(n1129), .B(n1130), .C(n1131), .D(n1132), .Z(
        n1121) );
  HS65_LH_AOI212X4 U1080 ( .A(n2557), .B(\registers[31][24] ), .C(n2554), .D(
        \registers[30][24] ), .E(n1133), .Z(n1132) );
  HS65_LH_AOI212X4 U1081 ( .A(n2545), .B(\registers[25][24] ), .C(n2542), .D(
        \registers[24][24] ), .E(n1134), .Z(n1131) );
  HS65_LH_MX41X7 U1082 ( .D0(n2533), .S0(\registers[16][24] ), .D1(n2530), 
        .S1(\registers[17][24] ), .D2(n2527), .S2(\registers[18][24] ), .D3(
        n2524), .S3(\registers[19][24] ), .Z(n1130) );
  HS65_LH_NAND4ABX3 U1083 ( .A(n1114), .B(n1115), .C(n1116), .D(n1117), .Z(
        n1106) );
  HS65_LH_AOI212X4 U1084 ( .A(n2557), .B(\registers[31][25] ), .C(n2554), .D(
        \registers[30][25] ), .E(n1118), .Z(n1117) );
  HS65_LH_AOI212X4 U1085 ( .A(n2545), .B(\registers[25][25] ), .C(n2542), .D(
        \registers[24][25] ), .E(n1119), .Z(n1116) );
  HS65_LH_MX41X7 U1086 ( .D0(n2533), .S0(\registers[16][25] ), .D1(n2530), 
        .S1(\registers[17][25] ), .D2(n2527), .S2(\registers[18][25] ), .D3(
        n2524), .S3(\registers[19][25] ), .Z(n1115) );
  HS65_LH_NAND4ABX3 U1087 ( .A(n1099), .B(n1100), .C(n1101), .D(n1102), .Z(
        n1091) );
  HS65_LH_AOI212X4 U1088 ( .A(n2557), .B(\registers[31][26] ), .C(n2554), .D(
        \registers[30][26] ), .E(n1103), .Z(n1102) );
  HS65_LH_AOI212X4 U1089 ( .A(n2545), .B(\registers[25][26] ), .C(n2542), .D(
        \registers[24][26] ), .E(n1104), .Z(n1101) );
  HS65_LH_MX41X7 U1090 ( .D0(n2533), .S0(\registers[16][26] ), .D1(n2530), 
        .S1(\registers[17][26] ), .D2(n2527), .S2(\registers[18][26] ), .D3(
        n2524), .S3(\registers[19][26] ), .Z(n1100) );
  HS65_LH_NAND4ABX3 U1091 ( .A(n1084), .B(n1085), .C(n1086), .D(n1087), .Z(
        n1076) );
  HS65_LH_AOI212X4 U1092 ( .A(n2557), .B(\registers[31][27] ), .C(n2554), .D(
        \registers[30][27] ), .E(n1088), .Z(n1087) );
  HS65_LH_AOI212X4 U1093 ( .A(n2545), .B(\registers[25][27] ), .C(n2542), .D(
        \registers[24][27] ), .E(n1089), .Z(n1086) );
  HS65_LH_MX41X7 U1094 ( .D0(n2533), .S0(\registers[16][27] ), .D1(n2530), 
        .S1(\registers[17][27] ), .D2(n2527), .S2(\registers[18][27] ), .D3(
        n2524), .S3(\registers[19][27] ), .Z(n1085) );
  HS65_LH_NAND4ABX3 U1095 ( .A(n1069), .B(n1070), .C(n1071), .D(n1072), .Z(
        n1061) );
  HS65_LH_AOI212X4 U1096 ( .A(n2557), .B(\registers[31][28] ), .C(n2554), .D(
        \registers[30][28] ), .E(n1073), .Z(n1072) );
  HS65_LH_AOI212X4 U1097 ( .A(n2545), .B(\registers[25][28] ), .C(n2542), .D(
        \registers[24][28] ), .E(n1074), .Z(n1071) );
  HS65_LH_MX41X7 U1098 ( .D0(n2533), .S0(\registers[16][28] ), .D1(n2530), 
        .S1(\registers[17][28] ), .D2(n2527), .S2(\registers[18][28] ), .D3(
        n2524), .S3(\registers[19][28] ), .Z(n1070) );
  HS65_LH_NAND4ABX3 U1099 ( .A(n1054), .B(n1055), .C(n1056), .D(n1057), .Z(
        n1046) );
  HS65_LH_AOI212X4 U1100 ( .A(n2557), .B(\registers[31][29] ), .C(n2554), .D(
        \registers[30][29] ), .E(n1058), .Z(n1057) );
  HS65_LH_AOI212X4 U1101 ( .A(n2545), .B(\registers[25][29] ), .C(n2542), .D(
        \registers[24][29] ), .E(n1059), .Z(n1056) );
  HS65_LH_MX41X7 U1102 ( .D0(n2533), .S0(\registers[16][29] ), .D1(n2530), 
        .S1(\registers[17][29] ), .D2(n2527), .S2(\registers[18][29] ), .D3(
        n2524), .S3(\registers[19][29] ), .Z(n1055) );
  HS65_LH_NAND4ABX3 U1103 ( .A(n1024), .B(n1025), .C(n1026), .D(n1027), .Z(
        n1016) );
  HS65_LH_AOI212X4 U1104 ( .A(n2557), .B(\registers[31][30] ), .C(n2554), .D(
        \registers[30][30] ), .E(n1028), .Z(n1027) );
  HS65_LH_AOI212X4 U1105 ( .A(n2545), .B(\registers[25][30] ), .C(n2542), .D(
        \registers[24][30] ), .E(n1029), .Z(n1026) );
  HS65_LH_MX41X7 U1106 ( .D0(n2533), .S0(\registers[16][30] ), .D1(n2530), 
        .S1(\registers[17][30] ), .D2(n2527), .S2(\registers[18][30] ), .D3(
        n2524), .S3(\registers[19][30] ), .Z(n1025) );
  HS65_LH_NAND4ABX3 U1107 ( .A(n1009), .B(n1010), .C(n1011), .D(n1012), .Z(
        n1001) );
  HS65_LH_AOI212X4 U1108 ( .A(n2557), .B(\registers[31][31] ), .C(n2554), .D(
        \registers[30][31] ), .E(n1013), .Z(n1012) );
  HS65_LH_AOI212X4 U1109 ( .A(n2545), .B(\registers[25][31] ), .C(n2542), .D(
        \registers[24][31] ), .E(n1014), .Z(n1011) );
  HS65_LH_MX41X7 U1110 ( .D0(n2533), .S0(\registers[16][31] ), .D1(n2531), 
        .S1(\registers[17][31] ), .D2(n2527), .S2(\registers[18][31] ), .D3(
        n2525), .S3(\registers[19][31] ), .Z(n1010) );
  HS65_LH_NAND4ABX3 U1111 ( .A(n820), .B(n821), .C(n822), .D(n823), .Z(n819)
         );
  HS65_LH_NAND3X5 U1112 ( .A(n2968), .B(n2969), .C(n2970), .Z(n821) );
  HS65_LH_AOI212X4 U1113 ( .A(\registers[13][10] ), .B(n2694), .C(
        \registers[12][10] ), .D(n2691), .E(n824), .Z(n823) );
  HS65_LH_AOI212X4 U1114 ( .A(\registers[11][10] ), .B(n2682), .C(
        \registers[10][10] ), .D(n2679), .E(n825), .Z(n822) );
  HS65_LH_AND2X4 U1115 ( .A(n847), .B(\regfile_i[ADRREAD1][0] ), .Z(n840) );
  HS65_LH_AND2X4 U1116 ( .A(n1375), .B(\regfile_i[ADRREAD0][0] ), .Z(n1368) );
  HS65_LH_AND2X4 U1117 ( .A(n859), .B(\regfile_i[ADRREAD1][0] ), .Z(n856) );
  HS65_LH_AND2X4 U1118 ( .A(n1387), .B(\regfile_i[ADRREAD0][0] ), .Z(n1384) );
  HS65_LH_AND2X4 U1119 ( .A(n862), .B(\regfile_i[ADRREAD1][0] ), .Z(n860) );
  HS65_LH_AND2X4 U1120 ( .A(n850), .B(\regfile_i[ADRREAD1][0] ), .Z(n848) );
  HS65_LH_AND2X4 U1121 ( .A(n1390), .B(\regfile_i[ADRREAD0][0] ), .Z(n1388) );
  HS65_LH_AND2X4 U1122 ( .A(n1378), .B(\regfile_i[ADRREAD0][0] ), .Z(n1376) );
  HS65_LH_NOR2X6 U1123 ( .A(n2902), .B(\regfile_i[ADRREAD1][3] ), .Z(n862) );
  HS65_LH_NOR2X6 U1124 ( .A(n2907), .B(\regfile_i[ADRREAD0][3] ), .Z(n1390) );
  HS65_LH_NOR2X6 U1125 ( .A(\regfile_i[ADRREAD1][3] ), .B(
        \regfile_i[ADRREAD1][4] ), .Z(n850) );
  HS65_LH_NOR2X6 U1126 ( .A(n2901), .B(\regfile_i[ADRREAD1][4] ), .Z(n847) );
  HS65_LH_NOR2X6 U1127 ( .A(\regfile_i[ADRREAD0][3] ), .B(
        \regfile_i[ADRREAD0][4] ), .Z(n1378) );
  HS65_LH_NOR2X6 U1128 ( .A(n2906), .B(\regfile_i[ADRREAD0][4] ), .Z(n1375) );
  HS65_LH_MX41X7 U1129 ( .D0(\registers[20][0] ), .S0(n2613), .D1(
        \registers[21][0] ), .S1(n2610), .D2(\registers[22][0] ), .S2(n2607), 
        .D3(\registers[23][0] ), .S3(n2604), .Z(n851) );
  HS65_LH_MX41X7 U1130 ( .D0(\registers[4][0] ), .S0(n2661), .D1(
        \registers[5][0] ), .S1(n2658), .D2(\registers[6][0] ), .S2(n2655), 
        .D3(\registers[7][0] ), .S3(n2652), .Z(n835) );
  HS65_LH_MX41X7 U1131 ( .D0(\registers[20][1] ), .S0(n2613), .D1(
        \registers[21][1] ), .S1(n2610), .D2(\registers[22][1] ), .S2(n2607), 
        .D3(\registers[23][1] ), .S3(n2604), .Z(n676) );
  HS65_LH_MX41X7 U1132 ( .D0(\registers[4][1] ), .S0(n2661), .D1(
        \registers[5][1] ), .S1(n2658), .D2(\registers[6][1] ), .S2(n2655), 
        .D3(\registers[7][1] ), .S3(n2652), .Z(n670) );
  HS65_LH_MX41X7 U1133 ( .D0(\registers[20][2] ), .S0(n2614), .D1(
        \registers[21][2] ), .S1(n2611), .D2(\registers[22][2] ), .S2(n2608), 
        .D3(\registers[23][2] ), .S3(n2605), .Z(n511) );
  HS65_LH_MX41X7 U1134 ( .D0(\registers[4][2] ), .S0(n2662), .D1(
        \registers[5][2] ), .S1(n2659), .D2(\registers[6][2] ), .S2(n2656), 
        .D3(\registers[7][2] ), .S3(n2653), .Z(n505) );
  HS65_LH_MX41X7 U1135 ( .D0(\registers[20][3] ), .S0(n2615), .D1(
        \registers[21][3] ), .S1(n2612), .D2(\registers[22][3] ), .S2(n2609), 
        .D3(\registers[23][3] ), .S3(n2606), .Z(n466) );
  HS65_LH_MX41X7 U1136 ( .D0(\registers[4][3] ), .S0(n2663), .D1(
        \registers[5][3] ), .S1(n2660), .D2(\registers[6][3] ), .S2(n2657), 
        .D3(\registers[7][3] ), .S3(n2654), .Z(n460) );
  HS65_LH_MX41X7 U1137 ( .D0(\registers[20][4] ), .S0(n2615), .D1(
        \registers[21][4] ), .S1(n2612), .D2(\registers[22][4] ), .S2(n2609), 
        .D3(\registers[23][4] ), .S3(n2606), .Z(n451) );
  HS65_LH_MX41X7 U1138 ( .D0(\registers[4][4] ), .S0(n2663), .D1(
        \registers[5][4] ), .S1(n2660), .D2(\registers[6][4] ), .S2(n2657), 
        .D3(\registers[7][4] ), .S3(n2654), .Z(n445) );
  HS65_LH_MX41X7 U1139 ( .D0(\registers[20][5] ), .S0(n2615), .D1(
        \registers[21][5] ), .S1(n2612), .D2(\registers[22][5] ), .S2(n2609), 
        .D3(\registers[23][5] ), .S3(n2606), .Z(n436) );
  HS65_LH_MX41X7 U1140 ( .D0(\registers[4][5] ), .S0(n2663), .D1(
        \registers[5][5] ), .S1(n2660), .D2(\registers[6][5] ), .S2(n2657), 
        .D3(\registers[7][5] ), .S3(n2654), .Z(n430) );
  HS65_LH_MX41X7 U1141 ( .D0(\registers[20][6] ), .S0(n2615), .D1(
        \registers[21][6] ), .S1(n2612), .D2(\registers[22][6] ), .S2(n2609), 
        .D3(\registers[23][6] ), .S3(n2606), .Z(n421) );
  HS65_LH_MX41X7 U1142 ( .D0(\registers[4][6] ), .S0(n2663), .D1(
        \registers[5][6] ), .S1(n2660), .D2(\registers[6][6] ), .S2(n2657), 
        .D3(\registers[7][6] ), .S3(n2654), .Z(n415) );
  HS65_LH_MX41X7 U1143 ( .D0(\registers[20][7] ), .S0(n2615), .D1(
        \registers[21][7] ), .S1(n2612), .D2(\registers[22][7] ), .S2(n2609), 
        .D3(\registers[23][7] ), .S3(n2606), .Z(n406) );
  HS65_LH_MX41X7 U1144 ( .D0(\registers[4][7] ), .S0(n2663), .D1(
        \registers[5][7] ), .S1(n2660), .D2(\registers[6][7] ), .S2(n2657), 
        .D3(\registers[7][7] ), .S3(n2654), .Z(n400) );
  HS65_LH_MX41X7 U1145 ( .D0(\registers[20][8] ), .S0(n2615), .D1(
        \registers[21][8] ), .S1(n2612), .D2(\registers[22][8] ), .S2(n2609), 
        .D3(\registers[23][8] ), .S3(n2606), .Z(n391) );
  HS65_LH_MX41X7 U1146 ( .D0(\registers[4][8] ), .S0(n2663), .D1(
        \registers[5][8] ), .S1(n2660), .D2(\registers[6][8] ), .S2(n2657), 
        .D3(\registers[7][8] ), .S3(n2654), .Z(n385) );
  HS65_LH_MX41X7 U1147 ( .D0(\registers[20][9] ), .S0(n2615), .D1(
        \registers[21][9] ), .S1(n2612), .D2(\registers[22][9] ), .S2(n2609), 
        .D3(\registers[23][9] ), .S3(n2606), .Z(n360) );
  HS65_LH_MX41X7 U1148 ( .D0(\registers[4][9] ), .S0(n2663), .D1(
        \registers[5][9] ), .S1(n2660), .D2(\registers[6][9] ), .S2(n2657), 
        .D3(\registers[7][9] ), .S3(n2654), .Z(n338) );
  HS65_LH_MX41X7 U1149 ( .D0(\registers[20][10] ), .S0(n2613), .D1(
        \registers[21][10] ), .S1(n2610), .D2(\registers[22][10] ), .S2(n2607), 
        .D3(\registers[23][10] ), .S3(n2604), .Z(n826) );
  HS65_LH_MX41X7 U1150 ( .D0(\registers[4][10] ), .S0(n2661), .D1(
        \registers[5][10] ), .S1(n2658), .D2(\registers[6][10] ), .S2(n2655), 
        .D3(\registers[7][10] ), .S3(n2652), .Z(n820) );
  HS65_LH_MX41X7 U1151 ( .D0(\registers[20][11] ), .S0(n2613), .D1(
        \registers[21][11] ), .S1(n2610), .D2(\registers[22][11] ), .S2(n2607), 
        .D3(\registers[23][11] ), .S3(n2604), .Z(n811) );
  HS65_LH_MX41X7 U1152 ( .D0(\registers[4][11] ), .S0(n2661), .D1(
        \registers[5][11] ), .S1(n2658), .D2(\registers[6][11] ), .S2(n2655), 
        .D3(\registers[7][11] ), .S3(n2652), .Z(n805) );
  HS65_LH_MX41X7 U1153 ( .D0(\registers[20][12] ), .S0(n2613), .D1(
        \registers[21][12] ), .S1(n2610), .D2(\registers[22][12] ), .S2(n2607), 
        .D3(\registers[23][12] ), .S3(n2604), .Z(n796) );
  HS65_LH_MX41X7 U1154 ( .D0(\registers[4][12] ), .S0(n2661), .D1(
        \registers[5][12] ), .S1(n2658), .D2(\registers[6][12] ), .S2(n2655), 
        .D3(\registers[7][12] ), .S3(n2652), .Z(n790) );
  HS65_LH_MX41X7 U1155 ( .D0(\registers[20][13] ), .S0(n2613), .D1(
        \registers[21][13] ), .S1(n2610), .D2(\registers[22][13] ), .S2(n2607), 
        .D3(\registers[23][13] ), .S3(n2604), .Z(n781) );
  HS65_LH_MX41X7 U1156 ( .D0(\registers[4][13] ), .S0(n2661), .D1(
        \registers[5][13] ), .S1(n2658), .D2(\registers[6][13] ), .S2(n2655), 
        .D3(\registers[7][13] ), .S3(n2652), .Z(n775) );
  HS65_LH_MX41X7 U1157 ( .D0(\registers[20][14] ), .S0(n2613), .D1(
        \registers[21][14] ), .S1(n2610), .D2(\registers[22][14] ), .S2(n2607), 
        .D3(\registers[23][14] ), .S3(n2604), .Z(n766) );
  HS65_LH_MX41X7 U1158 ( .D0(\registers[4][14] ), .S0(n2661), .D1(
        \registers[5][14] ), .S1(n2658), .D2(\registers[6][14] ), .S2(n2655), 
        .D3(\registers[7][14] ), .S3(n2652), .Z(n760) );
  HS65_LH_MX41X7 U1159 ( .D0(\registers[20][15] ), .S0(n2613), .D1(
        \registers[21][15] ), .S1(n2610), .D2(\registers[22][15] ), .S2(n2607), 
        .D3(\registers[23][15] ), .S3(n2604), .Z(n751) );
  HS65_LH_MX41X7 U1160 ( .D0(\registers[4][15] ), .S0(n2661), .D1(
        \registers[5][15] ), .S1(n2658), .D2(\registers[6][15] ), .S2(n2655), 
        .D3(\registers[7][15] ), .S3(n2652), .Z(n745) );
  HS65_LH_MX41X7 U1161 ( .D0(\registers[20][16] ), .S0(n2613), .D1(
        \registers[21][16] ), .S1(n2610), .D2(\registers[22][16] ), .S2(n2607), 
        .D3(\registers[23][16] ), .S3(n2604), .Z(n736) );
  HS65_LH_MX41X7 U1162 ( .D0(\registers[4][16] ), .S0(n2661), .D1(
        \registers[5][16] ), .S1(n2658), .D2(\registers[6][16] ), .S2(n2655), 
        .D3(\registers[7][16] ), .S3(n2652), .Z(n730) );
  HS65_LH_MX41X7 U1163 ( .D0(\registers[20][17] ), .S0(n2613), .D1(
        \registers[21][17] ), .S1(n2610), .D2(\registers[22][17] ), .S2(n2607), 
        .D3(\registers[23][17] ), .S3(n2604), .Z(n721) );
  HS65_LH_MX41X7 U1164 ( .D0(\registers[4][17] ), .S0(n2661), .D1(
        \registers[5][17] ), .S1(n2658), .D2(\registers[6][17] ), .S2(n2655), 
        .D3(\registers[7][17] ), .S3(n2652), .Z(n715) );
  HS65_LH_MX41X7 U1165 ( .D0(\registers[20][18] ), .S0(n2613), .D1(
        \registers[21][18] ), .S1(n2610), .D2(\registers[22][18] ), .S2(n2607), 
        .D3(\registers[23][18] ), .S3(n2604), .Z(n706) );
  HS65_LH_MX41X7 U1166 ( .D0(\registers[4][18] ), .S0(n2661), .D1(
        \registers[5][18] ), .S1(n2658), .D2(\registers[6][18] ), .S2(n2655), 
        .D3(\registers[7][18] ), .S3(n2652), .Z(n700) );
  HS65_LH_MX41X7 U1167 ( .D0(\registers[20][19] ), .S0(n2613), .D1(
        \registers[21][19] ), .S1(n2610), .D2(\registers[22][19] ), .S2(n2607), 
        .D3(\registers[23][19] ), .S3(n2604), .Z(n691) );
  HS65_LH_MX41X7 U1168 ( .D0(\registers[4][19] ), .S0(n2661), .D1(
        \registers[5][19] ), .S1(n2658), .D2(\registers[6][19] ), .S2(n2655), 
        .D3(\registers[7][19] ), .S3(n2652), .Z(n685) );
  HS65_LH_MX41X7 U1169 ( .D0(\registers[20][20] ), .S0(n2614), .D1(
        \registers[21][20] ), .S1(n2611), .D2(\registers[22][20] ), .S2(n2608), 
        .D3(\registers[23][20] ), .S3(n2605), .Z(n661) );
  HS65_LH_MX41X7 U1170 ( .D0(\registers[4][20] ), .S0(n2662), .D1(
        \registers[5][20] ), .S1(n2659), .D2(\registers[6][20] ), .S2(n2656), 
        .D3(\registers[7][20] ), .S3(n2653), .Z(n655) );
  HS65_LH_MX41X7 U1171 ( .D0(\registers[20][21] ), .S0(n2614), .D1(
        \registers[21][21] ), .S1(n2611), .D2(\registers[22][21] ), .S2(n2608), 
        .D3(\registers[23][21] ), .S3(n2605), .Z(n646) );
  HS65_LH_MX41X7 U1172 ( .D0(\registers[4][21] ), .S0(n2662), .D1(
        \registers[5][21] ), .S1(n2659), .D2(\registers[6][21] ), .S2(n2656), 
        .D3(\registers[7][21] ), .S3(n2653), .Z(n640) );
  HS65_LH_MX41X7 U1173 ( .D0(\registers[20][22] ), .S0(n2614), .D1(
        \registers[21][22] ), .S1(n2611), .D2(\registers[22][22] ), .S2(n2608), 
        .D3(\registers[23][22] ), .S3(n2605), .Z(n631) );
  HS65_LH_MX41X7 U1174 ( .D0(\registers[4][22] ), .S0(n2662), .D1(
        \registers[5][22] ), .S1(n2659), .D2(\registers[6][22] ), .S2(n2656), 
        .D3(\registers[7][22] ), .S3(n2653), .Z(n625) );
  HS65_LH_MX41X7 U1175 ( .D0(\registers[20][23] ), .S0(n2614), .D1(
        \registers[21][23] ), .S1(n2611), .D2(\registers[22][23] ), .S2(n2608), 
        .D3(\registers[23][23] ), .S3(n2605), .Z(n616) );
  HS65_LH_MX41X7 U1176 ( .D0(\registers[4][23] ), .S0(n2662), .D1(
        \registers[5][23] ), .S1(n2659), .D2(\registers[6][23] ), .S2(n2656), 
        .D3(\registers[7][23] ), .S3(n2653), .Z(n610) );
  HS65_LH_MX41X7 U1177 ( .D0(\registers[20][24] ), .S0(n2614), .D1(
        \registers[21][24] ), .S1(n2611), .D2(\registers[22][24] ), .S2(n2608), 
        .D3(\registers[23][24] ), .S3(n2605), .Z(n601) );
  HS65_LH_MX41X7 U1178 ( .D0(\registers[4][24] ), .S0(n2662), .D1(
        \registers[5][24] ), .S1(n2659), .D2(\registers[6][24] ), .S2(n2656), 
        .D3(\registers[7][24] ), .S3(n2653), .Z(n595) );
  HS65_LH_MX41X7 U1179 ( .D0(\registers[20][25] ), .S0(n2614), .D1(
        \registers[21][25] ), .S1(n2611), .D2(\registers[22][25] ), .S2(n2608), 
        .D3(\registers[23][25] ), .S3(n2605), .Z(n586) );
  HS65_LH_MX41X7 U1180 ( .D0(\registers[4][25] ), .S0(n2662), .D1(
        \registers[5][25] ), .S1(n2659), .D2(\registers[6][25] ), .S2(n2656), 
        .D3(\registers[7][25] ), .S3(n2653), .Z(n580) );
  HS65_LH_MX41X7 U1181 ( .D0(\registers[20][26] ), .S0(n2614), .D1(
        \registers[21][26] ), .S1(n2611), .D2(\registers[22][26] ), .S2(n2608), 
        .D3(\registers[23][26] ), .S3(n2605), .Z(n571) );
  HS65_LH_MX41X7 U1182 ( .D0(\registers[4][26] ), .S0(n2662), .D1(
        \registers[5][26] ), .S1(n2659), .D2(\registers[6][26] ), .S2(n2656), 
        .D3(\registers[7][26] ), .S3(n2653), .Z(n565) );
  HS65_LH_MX41X7 U1183 ( .D0(\registers[20][27] ), .S0(n2614), .D1(
        \registers[21][27] ), .S1(n2611), .D2(\registers[22][27] ), .S2(n2608), 
        .D3(\registers[23][27] ), .S3(n2605), .Z(n556) );
  HS65_LH_MX41X7 U1184 ( .D0(\registers[4][27] ), .S0(n2662), .D1(
        \registers[5][27] ), .S1(n2659), .D2(\registers[6][27] ), .S2(n2656), 
        .D3(\registers[7][27] ), .S3(n2653), .Z(n550) );
  HS65_LH_MX41X7 U1185 ( .D0(\registers[20][28] ), .S0(n2614), .D1(
        \registers[21][28] ), .S1(n2611), .D2(\registers[22][28] ), .S2(n2608), 
        .D3(\registers[23][28] ), .S3(n2605), .Z(n541) );
  HS65_LH_MX41X7 U1186 ( .D0(\registers[4][28] ), .S0(n2662), .D1(
        \registers[5][28] ), .S1(n2659), .D2(\registers[6][28] ), .S2(n2656), 
        .D3(\registers[7][28] ), .S3(n2653), .Z(n535) );
  HS65_LH_MX41X7 U1187 ( .D0(\registers[20][29] ), .S0(n2614), .D1(
        \registers[21][29] ), .S1(n2611), .D2(\registers[22][29] ), .S2(n2608), 
        .D3(\registers[23][29] ), .S3(n2605), .Z(n526) );
  HS65_LH_MX41X7 U1188 ( .D0(\registers[4][29] ), .S0(n2662), .D1(
        \registers[5][29] ), .S1(n2659), .D2(\registers[6][29] ), .S2(n2656), 
        .D3(\registers[7][29] ), .S3(n2653), .Z(n520) );
  HS65_LH_MX41X7 U1189 ( .D0(\registers[20][30] ), .S0(n2614), .D1(
        \registers[21][30] ), .S1(n2611), .D2(\registers[22][30] ), .S2(n2608), 
        .D3(\registers[23][30] ), .S3(n2605), .Z(n496) );
  HS65_LH_MX41X7 U1190 ( .D0(\registers[4][30] ), .S0(n2662), .D1(
        \registers[5][30] ), .S1(n2659), .D2(\registers[6][30] ), .S2(n2656), 
        .D3(\registers[7][30] ), .S3(n2653), .Z(n490) );
  HS65_LH_MX41X7 U1191 ( .D0(\registers[20][31] ), .S0(n2615), .D1(
        \registers[21][31] ), .S1(n2612), .D2(\registers[22][31] ), .S2(n2609), 
        .D3(\registers[23][31] ), .S3(n2606), .Z(n481) );
  HS65_LH_MX41X7 U1192 ( .D0(\registers[4][31] ), .S0(n2663), .D1(
        \registers[5][31] ), .S1(n2660), .D2(\registers[6][31] ), .S2(n2657), 
        .D3(\registers[7][31] ), .S3(n2654), .Z(n475) );
  HS65_LH_IVX9 U1193 ( .A(\regfile_i[ADRREAD1][0] ), .Z(n2898) );
  HS65_LH_IVX9 U1194 ( .A(\regfile_i[ADRREAD0][0] ), .Z(n2903) );
  HS65_LH_MX41X7 U1195 ( .D0(n2520), .S0(\registers[20][0] ), .D1(n2517), .S1(
        \registers[21][0] ), .D2(n2514), .S2(\registers[22][0] ), .D3(n2511), 
        .S3(\registers[23][0] ), .Z(n1379) );
  HS65_LH_MX41X7 U1196 ( .D0(n2568), .S0(\registers[4][0] ), .D1(n2565), .S1(
        \registers[5][0] ), .D2(n2562), .S2(\registers[6][0] ), .D3(n2559), 
        .S3(\registers[7][0] ), .Z(n1363) );
  HS65_LH_MX41X7 U1197 ( .D0(n2520), .S0(\registers[20][1] ), .D1(n2517), .S1(
        \registers[21][1] ), .D2(n2514), .S2(\registers[22][1] ), .D3(n2511), 
        .S3(\registers[23][1] ), .Z(n1204) );
  HS65_LH_MX41X7 U1198 ( .D0(n2568), .S0(\registers[4][1] ), .D1(n2565), .S1(
        \registers[5][1] ), .D2(n2562), .S2(\registers[6][1] ), .D3(n2559), 
        .S3(\registers[7][1] ), .Z(n1198) );
  HS65_LH_MX41X7 U1199 ( .D0(n2521), .S0(\registers[20][2] ), .D1(n2518), .S1(
        \registers[21][2] ), .D2(n2515), .S2(\registers[22][2] ), .D3(n2512), 
        .S3(\registers[23][2] ), .Z(n1039) );
  HS65_LH_MX41X7 U1200 ( .D0(n2569), .S0(\registers[4][2] ), .D1(n2566), .S1(
        \registers[5][2] ), .D2(n2563), .S2(\registers[6][2] ), .D3(n2560), 
        .S3(\registers[7][2] ), .Z(n1033) );
  HS65_LH_MX41X7 U1201 ( .D0(n2521), .S0(\registers[20][3] ), .D1(n2519), .S1(
        \registers[21][3] ), .D2(n2515), .S2(\registers[22][3] ), .D3(n2513), 
        .S3(\registers[23][3] ), .Z(n994) );
  HS65_LH_MX41X7 U1202 ( .D0(n2569), .S0(\registers[4][3] ), .D1(n2567), .S1(
        \registers[5][3] ), .D2(n2563), .S2(\registers[6][3] ), .D3(n2561), 
        .S3(\registers[7][3] ), .Z(n988) );
  HS65_LH_MX41X7 U1203 ( .D0(n2522), .S0(\registers[20][4] ), .D1(n2519), .S1(
        \registers[21][4] ), .D2(n2516), .S2(\registers[22][4] ), .D3(n2513), 
        .S3(\registers[23][4] ), .Z(n979) );
  HS65_LH_MX41X7 U1204 ( .D0(n2570), .S0(\registers[4][4] ), .D1(n2567), .S1(
        \registers[5][4] ), .D2(n2564), .S2(\registers[6][4] ), .D3(n2561), 
        .S3(\registers[7][4] ), .Z(n973) );
  HS65_LH_MX41X7 U1205 ( .D0(n2522), .S0(\registers[20][5] ), .D1(n2519), .S1(
        \registers[21][5] ), .D2(n2516), .S2(\registers[22][5] ), .D3(n2513), 
        .S3(\registers[23][5] ), .Z(n964) );
  HS65_LH_MX41X7 U1206 ( .D0(n2570), .S0(\registers[4][5] ), .D1(n2567), .S1(
        \registers[5][5] ), .D2(n2564), .S2(\registers[6][5] ), .D3(n2561), 
        .S3(\registers[7][5] ), .Z(n958) );
  HS65_LH_MX41X7 U1207 ( .D0(n2522), .S0(\registers[20][6] ), .D1(n2519), .S1(
        \registers[21][6] ), .D2(n2516), .S2(\registers[22][6] ), .D3(n2513), 
        .S3(\registers[23][6] ), .Z(n949) );
  HS65_LH_MX41X7 U1208 ( .D0(n2570), .S0(\registers[4][6] ), .D1(n2567), .S1(
        \registers[5][6] ), .D2(n2564), .S2(\registers[6][6] ), .D3(n2561), 
        .S3(\registers[7][6] ), .Z(n943) );
  HS65_LH_MX41X7 U1209 ( .D0(n2522), .S0(\registers[20][7] ), .D1(n2519), .S1(
        \registers[21][7] ), .D2(n2516), .S2(\registers[22][7] ), .D3(n2513), 
        .S3(\registers[23][7] ), .Z(n934) );
  HS65_LH_MX41X7 U1210 ( .D0(n2570), .S0(\registers[4][7] ), .D1(n2567), .S1(
        \registers[5][7] ), .D2(n2564), .S2(\registers[6][7] ), .D3(n2561), 
        .S3(\registers[7][7] ), .Z(n928) );
  HS65_LH_MX41X7 U1211 ( .D0(n2522), .S0(\registers[20][8] ), .D1(n2519), .S1(
        \registers[21][8] ), .D2(n2516), .S2(\registers[22][8] ), .D3(n2513), 
        .S3(\registers[23][8] ), .Z(n919) );
  HS65_LH_MX41X7 U1212 ( .D0(n2570), .S0(\registers[4][8] ), .D1(n2567), .S1(
        \registers[5][8] ), .D2(n2564), .S2(\registers[6][8] ), .D3(n2561), 
        .S3(\registers[7][8] ), .Z(n913) );
  HS65_LH_MX41X7 U1213 ( .D0(n2522), .S0(\registers[20][9] ), .D1(n2519), .S1(
        \registers[21][9] ), .D2(n2516), .S2(\registers[22][9] ), .D3(n2513), 
        .S3(\registers[23][9] ), .Z(n888) );
  HS65_LH_MX41X7 U1214 ( .D0(n2570), .S0(\registers[4][9] ), .D1(n2567), .S1(
        \registers[5][9] ), .D2(n2564), .S2(\registers[6][9] ), .D3(n2561), 
        .S3(\registers[7][9] ), .Z(n866) );
  HS65_LH_MX41X7 U1215 ( .D0(n2520), .S0(\registers[20][10] ), .D1(n2517), 
        .S1(\registers[21][10] ), .D2(n2514), .S2(\registers[22][10] ), .D3(
        n2511), .S3(\registers[23][10] ), .Z(n1354) );
  HS65_LH_MX41X7 U1216 ( .D0(n2568), .S0(\registers[4][10] ), .D1(n2565), .S1(
        \registers[5][10] ), .D2(n2562), .S2(\registers[6][10] ), .D3(n2559), 
        .S3(\registers[7][10] ), .Z(n1348) );
  HS65_LH_MX41X7 U1217 ( .D0(n2520), .S0(\registers[20][11] ), .D1(n2517), 
        .S1(\registers[21][11] ), .D2(n2514), .S2(\registers[22][11] ), .D3(
        n2511), .S3(\registers[23][11] ), .Z(n1339) );
  HS65_LH_MX41X7 U1218 ( .D0(n2568), .S0(\registers[4][11] ), .D1(n2565), .S1(
        \registers[5][11] ), .D2(n2562), .S2(\registers[6][11] ), .D3(n2559), 
        .S3(\registers[7][11] ), .Z(n1333) );
  HS65_LH_MX41X7 U1219 ( .D0(n2520), .S0(\registers[20][12] ), .D1(n2517), 
        .S1(\registers[21][12] ), .D2(n2514), .S2(\registers[22][12] ), .D3(
        n2511), .S3(\registers[23][12] ), .Z(n1324) );
  HS65_LH_MX41X7 U1220 ( .D0(n2568), .S0(\registers[4][12] ), .D1(n2565), .S1(
        \registers[5][12] ), .D2(n2562), .S2(\registers[6][12] ), .D3(n2559), 
        .S3(\registers[7][12] ), .Z(n1318) );
  HS65_LH_MX41X7 U1221 ( .D0(n2520), .S0(\registers[20][13] ), .D1(n2517), 
        .S1(\registers[21][13] ), .D2(n2514), .S2(\registers[22][13] ), .D3(
        n2511), .S3(\registers[23][13] ), .Z(n1309) );
  HS65_LH_MX41X7 U1222 ( .D0(n2568), .S0(\registers[4][13] ), .D1(n2565), .S1(
        \registers[5][13] ), .D2(n2562), .S2(\registers[6][13] ), .D3(n2559), 
        .S3(\registers[7][13] ), .Z(n1303) );
  HS65_LH_MX41X7 U1223 ( .D0(n2520), .S0(\registers[20][14] ), .D1(n2517), 
        .S1(\registers[21][14] ), .D2(n2514), .S2(\registers[22][14] ), .D3(
        n2511), .S3(\registers[23][14] ), .Z(n1294) );
  HS65_LH_MX41X7 U1224 ( .D0(n2568), .S0(\registers[4][14] ), .D1(n2565), .S1(
        \registers[5][14] ), .D2(n2562), .S2(\registers[6][14] ), .D3(n2559), 
        .S3(\registers[7][14] ), .Z(n1288) );
  HS65_LH_MX41X7 U1225 ( .D0(n2520), .S0(\registers[20][15] ), .D1(n2517), 
        .S1(\registers[21][15] ), .D2(n2514), .S2(\registers[22][15] ), .D3(
        n2511), .S3(\registers[23][15] ), .Z(n1279) );
  HS65_LH_MX41X7 U1226 ( .D0(n2568), .S0(\registers[4][15] ), .D1(n2565), .S1(
        \registers[5][15] ), .D2(n2562), .S2(\registers[6][15] ), .D3(n2559), 
        .S3(\registers[7][15] ), .Z(n1273) );
  HS65_LH_MX41X7 U1227 ( .D0(n2520), .S0(\registers[20][16] ), .D1(n2517), 
        .S1(\registers[21][16] ), .D2(n2514), .S2(\registers[22][16] ), .D3(
        n2511), .S3(\registers[23][16] ), .Z(n1264) );
  HS65_LH_MX41X7 U1228 ( .D0(n2568), .S0(\registers[4][16] ), .D1(n2565), .S1(
        \registers[5][16] ), .D2(n2562), .S2(\registers[6][16] ), .D3(n2559), 
        .S3(\registers[7][16] ), .Z(n1258) );
  HS65_LH_MX41X7 U1229 ( .D0(n2520), .S0(\registers[20][17] ), .D1(n2517), 
        .S1(\registers[21][17] ), .D2(n2514), .S2(\registers[22][17] ), .D3(
        n2511), .S3(\registers[23][17] ), .Z(n1249) );
  HS65_LH_MX41X7 U1230 ( .D0(n2568), .S0(\registers[4][17] ), .D1(n2565), .S1(
        \registers[5][17] ), .D2(n2562), .S2(\registers[6][17] ), .D3(n2559), 
        .S3(\registers[7][17] ), .Z(n1243) );
  HS65_LH_MX41X7 U1231 ( .D0(n2520), .S0(\registers[20][18] ), .D1(n2517), 
        .S1(\registers[21][18] ), .D2(n2514), .S2(\registers[22][18] ), .D3(
        n2511), .S3(\registers[23][18] ), .Z(n1234) );
  HS65_LH_MX41X7 U1232 ( .D0(n2568), .S0(\registers[4][18] ), .D1(n2565), .S1(
        \registers[5][18] ), .D2(n2562), .S2(\registers[6][18] ), .D3(n2559), 
        .S3(\registers[7][18] ), .Z(n1228) );
  HS65_LH_MX41X7 U1233 ( .D0(n2520), .S0(\registers[20][19] ), .D1(n2517), 
        .S1(\registers[21][19] ), .D2(n2514), .S2(\registers[22][19] ), .D3(
        n2511), .S3(\registers[23][19] ), .Z(n1219) );
  HS65_LH_MX41X7 U1234 ( .D0(n2568), .S0(\registers[4][19] ), .D1(n2565), .S1(
        \registers[5][19] ), .D2(n2562), .S2(\registers[6][19] ), .D3(n2559), 
        .S3(\registers[7][19] ), .Z(n1213) );
  HS65_LH_MX41X7 U1235 ( .D0(n2520), .S0(\registers[20][20] ), .D1(n2518), 
        .S1(\registers[21][20] ), .D2(n2514), .S2(\registers[22][20] ), .D3(
        n2512), .S3(\registers[23][20] ), .Z(n1189) );
  HS65_LH_MX41X7 U1236 ( .D0(n2568), .S0(\registers[4][20] ), .D1(n2566), .S1(
        \registers[5][20] ), .D2(n2562), .S2(\registers[6][20] ), .D3(n2560), 
        .S3(\registers[7][20] ), .Z(n1183) );
  HS65_LH_MX41X7 U1237 ( .D0(n2521), .S0(\registers[20][21] ), .D1(n2518), 
        .S1(\registers[21][21] ), .D2(n2515), .S2(\registers[22][21] ), .D3(
        n2512), .S3(\registers[23][21] ), .Z(n1174) );
  HS65_LH_MX41X7 U1238 ( .D0(n2569), .S0(\registers[4][21] ), .D1(n2566), .S1(
        \registers[5][21] ), .D2(n2563), .S2(\registers[6][21] ), .D3(n2560), 
        .S3(\registers[7][21] ), .Z(n1168) );
  HS65_LH_MX41X7 U1239 ( .D0(n2521), .S0(\registers[20][22] ), .D1(n2518), 
        .S1(\registers[21][22] ), .D2(n2515), .S2(\registers[22][22] ), .D3(
        n2512), .S3(\registers[23][22] ), .Z(n1159) );
  HS65_LH_MX41X7 U1240 ( .D0(n2569), .S0(\registers[4][22] ), .D1(n2566), .S1(
        \registers[5][22] ), .D2(n2563), .S2(\registers[6][22] ), .D3(n2560), 
        .S3(\registers[7][22] ), .Z(n1153) );
  HS65_LH_MX41X7 U1241 ( .D0(n2521), .S0(\registers[20][23] ), .D1(n2518), 
        .S1(\registers[21][23] ), .D2(n2515), .S2(\registers[22][23] ), .D3(
        n2512), .S3(\registers[23][23] ), .Z(n1144) );
  HS65_LH_MX41X7 U1242 ( .D0(n2569), .S0(\registers[4][23] ), .D1(n2566), .S1(
        \registers[5][23] ), .D2(n2563), .S2(\registers[6][23] ), .D3(n2560), 
        .S3(\registers[7][23] ), .Z(n1138) );
  HS65_LH_MX41X7 U1243 ( .D0(n2521), .S0(\registers[20][24] ), .D1(n2518), 
        .S1(\registers[21][24] ), .D2(n2515), .S2(\registers[22][24] ), .D3(
        n2512), .S3(\registers[23][24] ), .Z(n1129) );
  HS65_LH_MX41X7 U1244 ( .D0(n2569), .S0(\registers[4][24] ), .D1(n2566), .S1(
        \registers[5][24] ), .D2(n2563), .S2(\registers[6][24] ), .D3(n2560), 
        .S3(\registers[7][24] ), .Z(n1123) );
  HS65_LH_MX41X7 U1245 ( .D0(n2521), .S0(\registers[20][25] ), .D1(n2518), 
        .S1(\registers[21][25] ), .D2(n2515), .S2(\registers[22][25] ), .D3(
        n2512), .S3(\registers[23][25] ), .Z(n1114) );
  HS65_LH_MX41X7 U1246 ( .D0(n2569), .S0(\registers[4][25] ), .D1(n2566), .S1(
        \registers[5][25] ), .D2(n2563), .S2(\registers[6][25] ), .D3(n2560), 
        .S3(\registers[7][25] ), .Z(n1108) );
  HS65_LH_MX41X7 U1247 ( .D0(n2521), .S0(\registers[20][26] ), .D1(n2518), 
        .S1(\registers[21][26] ), .D2(n2515), .S2(\registers[22][26] ), .D3(
        n2512), .S3(\registers[23][26] ), .Z(n1099) );
  HS65_LH_MX41X7 U1248 ( .D0(n2569), .S0(\registers[4][26] ), .D1(n2566), .S1(
        \registers[5][26] ), .D2(n2563), .S2(\registers[6][26] ), .D3(n2560), 
        .S3(\registers[7][26] ), .Z(n1093) );
  HS65_LH_MX41X7 U1249 ( .D0(n2521), .S0(\registers[20][27] ), .D1(n2518), 
        .S1(\registers[21][27] ), .D2(n2515), .S2(\registers[22][27] ), .D3(
        n2512), .S3(\registers[23][27] ), .Z(n1084) );
  HS65_LH_MX41X7 U1250 ( .D0(n2569), .S0(\registers[4][27] ), .D1(n2566), .S1(
        \registers[5][27] ), .D2(n2563), .S2(\registers[6][27] ), .D3(n2560), 
        .S3(\registers[7][27] ), .Z(n1078) );
  HS65_LH_MX41X7 U1251 ( .D0(n2521), .S0(\registers[20][28] ), .D1(n2518), 
        .S1(\registers[21][28] ), .D2(n2515), .S2(\registers[22][28] ), .D3(
        n2512), .S3(\registers[23][28] ), .Z(n1069) );
  HS65_LH_MX41X7 U1252 ( .D0(n2569), .S0(\registers[4][28] ), .D1(n2566), .S1(
        \registers[5][28] ), .D2(n2563), .S2(\registers[6][28] ), .D3(n2560), 
        .S3(\registers[7][28] ), .Z(n1063) );
  HS65_LH_MX41X7 U1253 ( .D0(n2521), .S0(\registers[20][29] ), .D1(n2518), 
        .S1(\registers[21][29] ), .D2(n2515), .S2(\registers[22][29] ), .D3(
        n2512), .S3(\registers[23][29] ), .Z(n1054) );
  HS65_LH_MX41X7 U1254 ( .D0(n2569), .S0(\registers[4][29] ), .D1(n2566), .S1(
        \registers[5][29] ), .D2(n2563), .S2(\registers[6][29] ), .D3(n2560), 
        .S3(\registers[7][29] ), .Z(n1048) );
  HS65_LH_MX41X7 U1255 ( .D0(n2521), .S0(\registers[20][30] ), .D1(n2518), 
        .S1(\registers[21][30] ), .D2(n2515), .S2(\registers[22][30] ), .D3(
        n2512), .S3(\registers[23][30] ), .Z(n1024) );
  HS65_LH_MX41X7 U1256 ( .D0(n2569), .S0(\registers[4][30] ), .D1(n2566), .S1(
        \registers[5][30] ), .D2(n2563), .S2(\registers[6][30] ), .D3(n2560), 
        .S3(\registers[7][30] ), .Z(n1018) );
  HS65_LH_MX41X7 U1257 ( .D0(n2521), .S0(\registers[20][31] ), .D1(n2519), 
        .S1(\registers[21][31] ), .D2(n2515), .S2(\registers[22][31] ), .D3(
        n2513), .S3(\registers[23][31] ), .Z(n1009) );
  HS65_LH_MX41X7 U1258 ( .D0(n2569), .S0(\registers[4][31] ), .D1(n2567), .S1(
        \registers[5][31] ), .D2(n2563), .S2(\registers[6][31] ), .D3(n2561), 
        .S3(\registers[7][31] ), .Z(n1003) );
  HS65_LH_IVX9 U1259 ( .A(\regfile_i[ADRREAD1][4] ), .Z(n2902) );
  HS65_LH_IVX9 U1260 ( .A(\regfile_i[ADRREAD0][4] ), .Z(n2907) );
  HS65_LH_IVX9 U1261 ( .A(\regfile_i[ADRREAD1][2] ), .Z(n2900) );
  HS65_LH_IVX9 U1262 ( .A(\regfile_i[ADRREAD0][2] ), .Z(n2905) );
  HS65_LH_IVX9 U1263 ( .A(\regfile_i[ADRREAD1][3] ), .Z(n2901) );
  HS65_LH_IVX9 U1264 ( .A(\regfile_i[ADRREAD0][3] ), .Z(n2906) );
  HS65_LH_IVX9 U1265 ( .A(\regfile_i[ADRREAD1][1] ), .Z(n2899) );
  HS65_LH_IVX9 U1266 ( .A(\regfile_i[ADRREAD0][1] ), .Z(n2904) );
  HS65_LH_OAI21X3 U1267 ( .A(n2698), .B(n280), .C(n1360), .Z(
        \regfile_o[READ_DATA0][0] ) );
  HS65_LH_OAI21X3 U1268 ( .A(n1361), .B(n1362), .C(n278), .Z(n1360) );
  HS65_LH_NAND4ABX3 U1269 ( .A(n1363), .B(n1364), .C(n1365), .D(n1366), .Z(
        n1362) );
  HS65_LH_OAI21X3 U1270 ( .A(n2700), .B(n282), .C(n1195), .Z(
        \regfile_o[READ_DATA0][1] ) );
  HS65_LH_OAI21X3 U1271 ( .A(n1196), .B(n1197), .C(n279), .Z(n1195) );
  HS65_LH_NAND4ABX3 U1272 ( .A(n1198), .B(n1199), .C(n1200), .D(n1201), .Z(
        n1197) );
  HS65_LH_OAI21X3 U1273 ( .A(n2702), .B(n281), .C(n1030), .Z(
        \regfile_o[READ_DATA0][2] ) );
  HS65_LH_OAI21X3 U1274 ( .A(n1031), .B(n1032), .C(n280), .Z(n1030) );
  HS65_LH_NAND4ABX3 U1275 ( .A(n1033), .B(n1034), .C(n1035), .D(n1036), .Z(
        n1032) );
  HS65_LH_OAI21X3 U1276 ( .A(n2704), .B(n280), .C(n985), .Z(
        \regfile_o[READ_DATA0][3] ) );
  HS65_LH_OAI21X3 U1277 ( .A(n986), .B(n987), .C(n279), .Z(n985) );
  HS65_LH_NAND4ABX3 U1278 ( .A(n988), .B(n989), .C(n990), .D(n991), .Z(n987)
         );
  HS65_LH_OAI21X3 U1279 ( .A(n2706), .B(n281), .C(n970), .Z(
        \regfile_o[READ_DATA0][4] ) );
  HS65_LH_OAI21X3 U1280 ( .A(n971), .B(n972), .C(n279), .Z(n970) );
  HS65_LH_NAND4ABX3 U1281 ( .A(n973), .B(n974), .C(n975), .D(n976), .Z(n972)
         );
  HS65_LH_OAI21X3 U1282 ( .A(n2708), .B(n280), .C(n955), .Z(
        \regfile_o[READ_DATA0][5] ) );
  HS65_LH_OAI21X3 U1283 ( .A(n956), .B(n957), .C(n279), .Z(n955) );
  HS65_LH_NAND4ABX3 U1284 ( .A(n958), .B(n959), .C(n960), .D(n961), .Z(n957)
         );
  HS65_LH_OAI21X3 U1285 ( .A(n2710), .B(n280), .C(n940), .Z(
        \regfile_o[READ_DATA0][6] ) );
  HS65_LH_OAI21X3 U1286 ( .A(n941), .B(n942), .C(n278), .Z(n940) );
  HS65_LH_NAND4ABX3 U1287 ( .A(n943), .B(n944), .C(n945), .D(n946), .Z(n942)
         );
  HS65_LH_OAI21X3 U1288 ( .A(n2712), .B(n281), .C(n925), .Z(
        \regfile_o[READ_DATA0][7] ) );
  HS65_LH_OAI21X3 U1289 ( .A(n926), .B(n927), .C(n278), .Z(n925) );
  HS65_LH_NAND4ABX3 U1290 ( .A(n928), .B(n929), .C(n930), .D(n931), .Z(n927)
         );
  HS65_LH_OAI21X3 U1291 ( .A(n2714), .B(n280), .C(n910), .Z(
        \regfile_o[READ_DATA0][8] ) );
  HS65_LH_OAI21X3 U1292 ( .A(n911), .B(n912), .C(n278), .Z(n910) );
  HS65_LH_NAND4ABX3 U1293 ( .A(n913), .B(n914), .C(n915), .D(n916), .Z(n912)
         );
  HS65_LH_OAI21X3 U1294 ( .A(n2716), .B(n281), .C(n863), .Z(
        \regfile_o[READ_DATA0][9] ) );
  HS65_LH_OAI21X3 U1295 ( .A(n864), .B(n865), .C(n278), .Z(n863) );
  HS65_LH_NAND4ABX3 U1296 ( .A(n866), .B(n867), .C(n868), .D(n869), .Z(n865)
         );
  HS65_LH_OAI21X3 U1297 ( .A(n2718), .B(n282), .C(n1345), .Z(
        \regfile_o[READ_DATA0][10] ) );
  HS65_LH_OAI21X3 U1298 ( .A(n1346), .B(n1347), .C(n278), .Z(n1345) );
  HS65_LH_NAND4ABX3 U1299 ( .A(n1348), .B(n1349), .C(n1350), .D(n1351), .Z(
        n1347) );
  HS65_LH_OAI21X3 U1300 ( .A(n2720), .B(n282), .C(n1330), .Z(
        \regfile_o[READ_DATA0][11] ) );
  HS65_LH_OAI21X3 U1301 ( .A(n1331), .B(n1332), .C(n278), .Z(n1330) );
  HS65_LH_NAND4ABX3 U1302 ( .A(n1333), .B(n1334), .C(n1335), .D(n1336), .Z(
        n1332) );
  HS65_LH_OAI21X3 U1303 ( .A(n2722), .B(n282), .C(n1315), .Z(
        \regfile_o[READ_DATA0][12] ) );
  HS65_LH_OAI21X3 U1304 ( .A(n1316), .B(n1317), .C(n278), .Z(n1315) );
  HS65_LH_NAND4ABX3 U1305 ( .A(n1318), .B(n1319), .C(n1320), .D(n1321), .Z(
        n1317) );
  HS65_LH_OAI21X3 U1306 ( .A(n2724), .B(n282), .C(n1300), .Z(
        \regfile_o[READ_DATA0][13] ) );
  HS65_LH_OAI21X3 U1307 ( .A(n1301), .B(n1302), .C(n278), .Z(n1300) );
  HS65_LH_NAND4ABX3 U1308 ( .A(n1303), .B(n1304), .C(n1305), .D(n1306), .Z(
        n1302) );
  HS65_LH_OAI21X3 U1309 ( .A(n2726), .B(n282), .C(n1285), .Z(
        \regfile_o[READ_DATA0][14] ) );
  HS65_LH_OAI21X3 U1310 ( .A(n1286), .B(n1287), .C(n278), .Z(n1285) );
  HS65_LH_NAND4ABX3 U1311 ( .A(n1288), .B(n1289), .C(n1290), .D(n1291), .Z(
        n1287) );
  HS65_LH_OAI21X3 U1312 ( .A(n2728), .B(n282), .C(n1270), .Z(
        \regfile_o[READ_DATA0][15] ) );
  HS65_LH_OAI21X3 U1313 ( .A(n1271), .B(n1272), .C(n278), .Z(n1270) );
  HS65_LH_NAND4ABX3 U1314 ( .A(n1273), .B(n1274), .C(n1275), .D(n1276), .Z(
        n1272) );
  HS65_LH_OAI21X3 U1315 ( .A(n2730), .B(n282), .C(n1255), .Z(
        \regfile_o[READ_DATA0][16] ) );
  HS65_LH_OAI21X3 U1316 ( .A(n1256), .B(n1257), .C(n278), .Z(n1255) );
  HS65_LH_NAND4ABX3 U1317 ( .A(n1258), .B(n1259), .C(n1260), .D(n1261), .Z(
        n1257) );
  HS65_LH_OAI21X3 U1318 ( .A(n2732), .B(n282), .C(n1240), .Z(
        \regfile_o[READ_DATA0][17] ) );
  HS65_LH_OAI21X3 U1319 ( .A(n1241), .B(n1242), .C(n279), .Z(n1240) );
  HS65_LH_NAND4ABX3 U1320 ( .A(n1243), .B(n1244), .C(n1245), .D(n1246), .Z(
        n1242) );
  HS65_LH_OAI21X3 U1321 ( .A(n2734), .B(n282), .C(n1225), .Z(
        \regfile_o[READ_DATA0][18] ) );
  HS65_LH_OAI21X3 U1322 ( .A(n1226), .B(n1227), .C(n279), .Z(n1225) );
  HS65_LH_NAND4ABX3 U1323 ( .A(n1228), .B(n1229), .C(n1230), .D(n1231), .Z(
        n1227) );
  HS65_LH_OAI21X3 U1324 ( .A(n2736), .B(n282), .C(n1210), .Z(
        \regfile_o[READ_DATA0][19] ) );
  HS65_LH_OAI21X3 U1325 ( .A(n1211), .B(n1212), .C(n279), .Z(n1210) );
  HS65_LH_NAND4ABX3 U1326 ( .A(n1213), .B(n1214), .C(n1215), .D(n1216), .Z(
        n1212) );
  HS65_LH_OAI21X3 U1327 ( .A(n2738), .B(n282), .C(n1180), .Z(
        \regfile_o[READ_DATA0][20] ) );
  HS65_LH_OAI21X3 U1328 ( .A(n1181), .B(n1182), .C(n279), .Z(n1180) );
  HS65_LH_NAND4ABX3 U1329 ( .A(n1183), .B(n1184), .C(n1185), .D(n1186), .Z(
        n1182) );
  HS65_LH_OAI21X3 U1330 ( .A(n2740), .B(n282), .C(n1165), .Z(
        \regfile_o[READ_DATA0][21] ) );
  HS65_LH_OAI21X3 U1331 ( .A(n1166), .B(n1167), .C(n279), .Z(n1165) );
  HS65_LH_NAND4ABX3 U1332 ( .A(n1168), .B(n1169), .C(n1170), .D(n1171), .Z(
        n1167) );
  HS65_LH_OAI21X3 U1333 ( .A(n2742), .B(n281), .C(n1150), .Z(
        \regfile_o[READ_DATA0][22] ) );
  HS65_LH_OAI21X3 U1334 ( .A(n1151), .B(n1152), .C(n279), .Z(n1150) );
  HS65_LH_NAND4ABX3 U1335 ( .A(n1153), .B(n1154), .C(n1155), .D(n1156), .Z(
        n1152) );
  HS65_LH_OAI21X3 U1336 ( .A(n2744), .B(n281), .C(n1135), .Z(
        \regfile_o[READ_DATA0][23] ) );
  HS65_LH_OAI21X3 U1337 ( .A(n1136), .B(n1137), .C(n279), .Z(n1135) );
  HS65_LH_NAND4ABX3 U1338 ( .A(n1138), .B(n1139), .C(n1140), .D(n1141), .Z(
        n1137) );
  HS65_LH_OAI21X3 U1339 ( .A(n2746), .B(n281), .C(n1120), .Z(
        \regfile_o[READ_DATA0][24] ) );
  HS65_LH_OAI21X3 U1340 ( .A(n1121), .B(n1122), .C(n280), .Z(n1120) );
  HS65_LH_NAND4ABX3 U1341 ( .A(n1123), .B(n1124), .C(n1125), .D(n1126), .Z(
        n1122) );
  HS65_LH_OAI21X3 U1342 ( .A(n2748), .B(n281), .C(n1105), .Z(
        \regfile_o[READ_DATA0][25] ) );
  HS65_LH_OAI21X3 U1343 ( .A(n1106), .B(n1107), .C(n280), .Z(n1105) );
  HS65_LH_NAND4ABX3 U1344 ( .A(n1108), .B(n1109), .C(n1110), .D(n1111), .Z(
        n1107) );
  HS65_LH_OAI21X3 U1345 ( .A(n2750), .B(n281), .C(n1090), .Z(
        \regfile_o[READ_DATA0][26] ) );
  HS65_LH_OAI21X3 U1346 ( .A(n1091), .B(n1092), .C(n279), .Z(n1090) );
  HS65_LH_NAND4ABX3 U1347 ( .A(n1093), .B(n1094), .C(n1095), .D(n1096), .Z(
        n1092) );
  HS65_LH_OAI21X3 U1348 ( .A(n2752), .B(n281), .C(n1075), .Z(
        \regfile_o[READ_DATA0][27] ) );
  HS65_LH_OAI21X3 U1349 ( .A(n1076), .B(n1077), .C(n280), .Z(n1075) );
  HS65_LH_NAND4ABX3 U1350 ( .A(n1078), .B(n1079), .C(n1080), .D(n1081), .Z(
        n1077) );
  HS65_LH_OAI21X3 U1351 ( .A(n2754), .B(n281), .C(n1060), .Z(
        \regfile_o[READ_DATA0][28] ) );
  HS65_LH_OAI21X3 U1352 ( .A(n1061), .B(n1062), .C(n280), .Z(n1060) );
  HS65_LH_NAND4ABX3 U1353 ( .A(n1063), .B(n1064), .C(n1065), .D(n1066), .Z(
        n1062) );
  HS65_LH_OAI21X3 U1354 ( .A(n2756), .B(n281), .C(n1045), .Z(
        \regfile_o[READ_DATA0][29] ) );
  HS65_LH_OAI21X3 U1355 ( .A(n1046), .B(n1047), .C(n280), .Z(n1045) );
  HS65_LH_NAND4ABX3 U1356 ( .A(n1048), .B(n1049), .C(n1050), .D(n1051), .Z(
        n1047) );
  HS65_LH_OAI21X3 U1357 ( .A(n2758), .B(n281), .C(n1015), .Z(
        \regfile_o[READ_DATA0][30] ) );
  HS65_LH_OAI21X3 U1358 ( .A(n1016), .B(n1017), .C(n280), .Z(n1015) );
  HS65_LH_NAND4ABX3 U1359 ( .A(n1018), .B(n1019), .C(n1020), .D(n1021), .Z(
        n1017) );
  HS65_LH_OAI21X3 U1360 ( .A(n2760), .B(n281), .C(n1000), .Z(
        \regfile_o[READ_DATA0][31] ) );
  HS65_LH_OAI21X3 U1361 ( .A(n1001), .B(n1002), .C(n280), .Z(n1000) );
  HS65_LH_NAND4ABX3 U1362 ( .A(n1003), .B(n1004), .C(n1005), .D(n1006), .Z(
        n1002) );
  HS65_LH_OAI21X3 U1363 ( .A(n285), .B(n2698), .C(n832), .Z(
        \regfile_o[READ_DATA1][0] ) );
  HS65_LH_OAI21X3 U1364 ( .A(n833), .B(n834), .C(n283), .Z(n832) );
  HS65_LH_NAND4ABX3 U1365 ( .A(n835), .B(n836), .C(n837), .D(n838), .Z(n834)
         );
  HS65_LH_OAI21X3 U1366 ( .A(n287), .B(n2700), .C(n667), .Z(
        \regfile_o[READ_DATA1][1] ) );
  HS65_LH_OAI21X3 U1367 ( .A(n668), .B(n669), .C(n284), .Z(n667) );
  HS65_LH_NAND4ABX3 U1368 ( .A(n670), .B(n671), .C(n672), .D(n673), .Z(n669)
         );
  HS65_LH_OAI21X3 U1369 ( .A(n286), .B(n2702), .C(n502), .Z(
        \regfile_o[READ_DATA1][2] ) );
  HS65_LH_OAI21X3 U1370 ( .A(n503), .B(n504), .C(n285), .Z(n502) );
  HS65_LH_NAND4ABX3 U1371 ( .A(n505), .B(n506), .C(n507), .D(n508), .Z(n504)
         );
  HS65_LH_OAI21X3 U1372 ( .A(n285), .B(n2704), .C(n457), .Z(
        \regfile_o[READ_DATA1][3] ) );
  HS65_LH_OAI21X3 U1373 ( .A(n458), .B(n459), .C(n284), .Z(n457) );
  HS65_LH_NAND4ABX3 U1374 ( .A(n460), .B(n461), .C(n462), .D(n463), .Z(n459)
         );
  HS65_LH_OAI21X3 U1375 ( .A(n286), .B(n2706), .C(n442), .Z(
        \regfile_o[READ_DATA1][4] ) );
  HS65_LH_OAI21X3 U1376 ( .A(n443), .B(n444), .C(n284), .Z(n442) );
  HS65_LH_NAND4ABX3 U1377 ( .A(n445), .B(n446), .C(n447), .D(n448), .Z(n444)
         );
  HS65_LH_OAI21X3 U1378 ( .A(n285), .B(n2708), .C(n427), .Z(
        \regfile_o[READ_DATA1][5] ) );
  HS65_LH_OAI21X3 U1379 ( .A(n428), .B(n429), .C(n284), .Z(n427) );
  HS65_LH_NAND4ABX3 U1380 ( .A(n430), .B(n431), .C(n432), .D(n433), .Z(n429)
         );
  HS65_LH_OAI21X3 U1381 ( .A(n285), .B(n2710), .C(n412), .Z(
        \regfile_o[READ_DATA1][6] ) );
  HS65_LH_OAI21X3 U1382 ( .A(n413), .B(n414), .C(n283), .Z(n412) );
  HS65_LH_NAND4ABX3 U1383 ( .A(n415), .B(n416), .C(n417), .D(n418), .Z(n414)
         );
  HS65_LH_OAI21X3 U1384 ( .A(n286), .B(n2712), .C(n397), .Z(
        \regfile_o[READ_DATA1][7] ) );
  HS65_LH_OAI21X3 U1385 ( .A(n398), .B(n399), .C(n283), .Z(n397) );
  HS65_LH_NAND4ABX3 U1386 ( .A(n400), .B(n401), .C(n402), .D(n403), .Z(n399)
         );
  HS65_LH_OAI21X3 U1387 ( .A(n285), .B(n2714), .C(n382), .Z(
        \regfile_o[READ_DATA1][8] ) );
  HS65_LH_OAI21X3 U1388 ( .A(n383), .B(n384), .C(n283), .Z(n382) );
  HS65_LH_NAND4ABX3 U1389 ( .A(n385), .B(n386), .C(n387), .D(n388), .Z(n384)
         );
  HS65_LH_OAI21X3 U1390 ( .A(n286), .B(n2716), .C(n335), .Z(
        \regfile_o[READ_DATA1][9] ) );
  HS65_LH_OAI21X3 U1391 ( .A(n336), .B(n337), .C(n283), .Z(n335) );
  HS65_LH_NAND4ABX3 U1392 ( .A(n338), .B(n339), .C(n340), .D(n341), .Z(n337)
         );
  HS65_LH_OAI21X3 U1393 ( .A(n287), .B(n2720), .C(n802), .Z(
        \regfile_o[READ_DATA1][11] ) );
  HS65_LH_OAI21X3 U1394 ( .A(n803), .B(n804), .C(n283), .Z(n802) );
  HS65_LH_NAND4ABX3 U1395 ( .A(n805), .B(n806), .C(n807), .D(n808), .Z(n804)
         );
  HS65_LH_OAI21X3 U1396 ( .A(n287), .B(n2722), .C(n787), .Z(
        \regfile_o[READ_DATA1][12] ) );
  HS65_LH_OAI21X3 U1397 ( .A(n788), .B(n789), .C(n283), .Z(n787) );
  HS65_LH_NAND4ABX3 U1398 ( .A(n790), .B(n791), .C(n792), .D(n793), .Z(n789)
         );
  HS65_LH_OAI21X3 U1399 ( .A(n287), .B(n2724), .C(n772), .Z(
        \regfile_o[READ_DATA1][13] ) );
  HS65_LH_OAI21X3 U1400 ( .A(n773), .B(n774), .C(n283), .Z(n772) );
  HS65_LH_NAND4ABX3 U1401 ( .A(n775), .B(n776), .C(n777), .D(n778), .Z(n774)
         );
  HS65_LH_OAI21X3 U1402 ( .A(n287), .B(n2726), .C(n757), .Z(
        \regfile_o[READ_DATA1][14] ) );
  HS65_LH_OAI21X3 U1403 ( .A(n758), .B(n759), .C(n283), .Z(n757) );
  HS65_LH_NAND4ABX3 U1404 ( .A(n760), .B(n761), .C(n762), .D(n763), .Z(n759)
         );
  HS65_LH_OAI21X3 U1405 ( .A(n287), .B(n2728), .C(n742), .Z(
        \regfile_o[READ_DATA1][15] ) );
  HS65_LH_OAI21X3 U1406 ( .A(n743), .B(n744), .C(n283), .Z(n742) );
  HS65_LH_NAND4ABX3 U1407 ( .A(n745), .B(n746), .C(n747), .D(n748), .Z(n744)
         );
  HS65_LH_OAI21X3 U1408 ( .A(n287), .B(n2730), .C(n727), .Z(
        \regfile_o[READ_DATA1][16] ) );
  HS65_LH_OAI21X3 U1409 ( .A(n728), .B(n729), .C(n283), .Z(n727) );
  HS65_LH_NAND4ABX3 U1410 ( .A(n730), .B(n731), .C(n732), .D(n733), .Z(n729)
         );
  HS65_LH_OAI21X3 U1411 ( .A(n287), .B(n2732), .C(n712), .Z(
        \regfile_o[READ_DATA1][17] ) );
  HS65_LH_OAI21X3 U1412 ( .A(n713), .B(n714), .C(n284), .Z(n712) );
  HS65_LH_NAND4ABX3 U1413 ( .A(n715), .B(n716), .C(n717), .D(n718), .Z(n714)
         );
  HS65_LH_OAI21X3 U1414 ( .A(n287), .B(n2734), .C(n697), .Z(
        \regfile_o[READ_DATA1][18] ) );
  HS65_LH_OAI21X3 U1415 ( .A(n698), .B(n699), .C(n284), .Z(n697) );
  HS65_LH_NAND4ABX3 U1416 ( .A(n700), .B(n701), .C(n702), .D(n703), .Z(n699)
         );
  HS65_LH_OAI21X3 U1417 ( .A(n287), .B(n2736), .C(n682), .Z(
        \regfile_o[READ_DATA1][19] ) );
  HS65_LH_OAI21X3 U1418 ( .A(n683), .B(n684), .C(n284), .Z(n682) );
  HS65_LH_NAND4ABX3 U1419 ( .A(n685), .B(n686), .C(n687), .D(n688), .Z(n684)
         );
  HS65_LH_OAI21X3 U1420 ( .A(n287), .B(n2738), .C(n652), .Z(
        \regfile_o[READ_DATA1][20] ) );
  HS65_LH_OAI21X3 U1421 ( .A(n653), .B(n654), .C(n284), .Z(n652) );
  HS65_LH_NAND4ABX3 U1422 ( .A(n655), .B(n656), .C(n657), .D(n658), .Z(n654)
         );
  HS65_LH_OAI21X3 U1423 ( .A(n287), .B(n2740), .C(n637), .Z(
        \regfile_o[READ_DATA1][21] ) );
  HS65_LH_OAI21X3 U1424 ( .A(n638), .B(n639), .C(n284), .Z(n637) );
  HS65_LH_NAND4ABX3 U1425 ( .A(n640), .B(n641), .C(n642), .D(n643), .Z(n639)
         );
  HS65_LH_OAI21X3 U1426 ( .A(n287), .B(n2742), .C(n622), .Z(
        \regfile_o[READ_DATA1][22] ) );
  HS65_LH_OAI21X3 U1427 ( .A(n623), .B(n624), .C(n284), .Z(n622) );
  HS65_LH_NAND4ABX3 U1428 ( .A(n625), .B(n626), .C(n627), .D(n628), .Z(n624)
         );
  HS65_LH_OAI21X3 U1429 ( .A(n286), .B(n2744), .C(n607), .Z(
        \regfile_o[READ_DATA1][23] ) );
  HS65_LH_OAI21X3 U1430 ( .A(n608), .B(n609), .C(n284), .Z(n607) );
  HS65_LH_NAND4ABX3 U1431 ( .A(n610), .B(n611), .C(n612), .D(n613), .Z(n609)
         );
  HS65_LH_OAI21X3 U1432 ( .A(n286), .B(n2746), .C(n592), .Z(
        \regfile_o[READ_DATA1][24] ) );
  HS65_LH_OAI21X3 U1433 ( .A(n593), .B(n594), .C(n285), .Z(n592) );
  HS65_LH_NAND4ABX3 U1434 ( .A(n595), .B(n596), .C(n597), .D(n598), .Z(n594)
         );
  HS65_LH_OAI21X3 U1435 ( .A(n286), .B(n2748), .C(n577), .Z(
        \regfile_o[READ_DATA1][25] ) );
  HS65_LH_OAI21X3 U1436 ( .A(n578), .B(n579), .C(n285), .Z(n577) );
  HS65_LH_NAND4ABX3 U1437 ( .A(n580), .B(n581), .C(n582), .D(n583), .Z(n579)
         );
  HS65_LH_OAI21X3 U1438 ( .A(n286), .B(n2750), .C(n562), .Z(
        \regfile_o[READ_DATA1][26] ) );
  HS65_LH_OAI21X3 U1439 ( .A(n563), .B(n564), .C(n284), .Z(n562) );
  HS65_LH_NAND4ABX3 U1440 ( .A(n565), .B(n566), .C(n567), .D(n568), .Z(n564)
         );
  HS65_LH_OAI21X3 U1441 ( .A(n286), .B(n2752), .C(n547), .Z(
        \regfile_o[READ_DATA1][27] ) );
  HS65_LH_OAI21X3 U1442 ( .A(n548), .B(n549), .C(n285), .Z(n547) );
  HS65_LH_NAND4ABX3 U1443 ( .A(n550), .B(n551), .C(n552), .D(n553), .Z(n549)
         );
  HS65_LH_OAI21X3 U1444 ( .A(n286), .B(n2754), .C(n532), .Z(
        \regfile_o[READ_DATA1][28] ) );
  HS65_LH_OAI21X3 U1445 ( .A(n533), .B(n534), .C(n285), .Z(n532) );
  HS65_LH_NAND4ABX3 U1446 ( .A(n535), .B(n536), .C(n537), .D(n538), .Z(n534)
         );
  HS65_LH_OAI21X3 U1447 ( .A(n286), .B(n2756), .C(n517), .Z(
        \regfile_o[READ_DATA1][29] ) );
  HS65_LH_OAI21X3 U1448 ( .A(n518), .B(n519), .C(n285), .Z(n517) );
  HS65_LH_NAND4ABX3 U1449 ( .A(n520), .B(n521), .C(n522), .D(n523), .Z(n519)
         );
  HS65_LH_OAI21X3 U1450 ( .A(n286), .B(n2758), .C(n487), .Z(
        \regfile_o[READ_DATA1][30] ) );
  HS65_LH_OAI21X3 U1451 ( .A(n488), .B(n489), .C(n285), .Z(n487) );
  HS65_LH_NAND4ABX3 U1452 ( .A(n490), .B(n491), .C(n492), .D(n493), .Z(n489)
         );
  HS65_LH_OAI21X3 U1453 ( .A(n286), .B(n2760), .C(n472), .Z(
        \regfile_o[READ_DATA1][31] ) );
  HS65_LH_OAI21X3 U1454 ( .A(n473), .B(n474), .C(n285), .Z(n472) );
  HS65_LH_NAND4ABX3 U1455 ( .A(n475), .B(n476), .C(n477), .D(n478), .Z(n474)
         );
  HS65_LH_OAI21X3 U1456 ( .A(n287), .B(n2718), .C(n817), .Z(
        \regfile_o[READ_DATA1][10] ) );
  HS65_LH_OAI21X3 U1457 ( .A(n818), .B(n819), .C(n283), .Z(n817) );
  HS65_LH_AOI212X4 U1458 ( .A(\registers[11][3] ), .B(n2684), .C(
        \registers[10][3] ), .D(n2680), .E(n465), .Z(n462) );
  HS65_LH_OAI22X6 U1459 ( .A(n2678), .B(n253), .C(n2674), .D(n221), .Z(n465)
         );
  HS65_LH_AOI212X4 U1460 ( .A(\registers[11][4] ), .B(n2684), .C(
        \registers[10][4] ), .D(n2681), .E(n450), .Z(n447) );
  HS65_LH_OAI22X6 U1461 ( .A(n2678), .B(n252), .C(n2675), .D(n220), .Z(n450)
         );
  HS65_LH_AOI212X4 U1462 ( .A(\registers[11][5] ), .B(n2684), .C(
        \registers[10][5] ), .D(n2681), .E(n435), .Z(n432) );
  HS65_LH_OAI22X6 U1463 ( .A(n2678), .B(n251), .C(n2675), .D(n219), .Z(n435)
         );
  HS65_LH_AOI212X4 U1464 ( .A(\registers[11][6] ), .B(n2684), .C(
        \registers[10][6] ), .D(n2681), .E(n420), .Z(n417) );
  HS65_LH_OAI22X6 U1465 ( .A(n2678), .B(n250), .C(n2675), .D(n218), .Z(n420)
         );
  HS65_LH_AOI212X4 U1466 ( .A(\registers[11][7] ), .B(n2684), .C(
        \registers[10][7] ), .D(n2681), .E(n405), .Z(n402) );
  HS65_LH_OAI22X6 U1467 ( .A(n2678), .B(n249), .C(n2675), .D(n217), .Z(n405)
         );
  HS65_LH_AOI212X4 U1468 ( .A(\registers[11][8] ), .B(n2684), .C(
        \registers[10][8] ), .D(n2681), .E(n390), .Z(n387) );
  HS65_LH_OAI22X6 U1469 ( .A(n2678), .B(n248), .C(n2675), .D(n216), .Z(n390)
         );
  HS65_LH_AOI212X4 U1470 ( .A(\registers[11][9] ), .B(n2684), .C(
        \registers[10][9] ), .D(n2681), .E(n349), .Z(n340) );
  HS65_LH_OAI22X6 U1471 ( .A(n2678), .B(n247), .C(n2675), .D(n215), .Z(n349)
         );
  HS65_LH_AOI212X4 U1472 ( .A(\registers[11][31] ), .B(n2684), .C(
        \registers[10][31] ), .D(n2680), .E(n480), .Z(n477) );
  HS65_LH_OAI22X6 U1473 ( .A(n2678), .B(n225), .C(n2674), .D(n193), .Z(n480)
         );
  HS65_LH_AOI212X4 U1474 ( .A(\registers[13][0] ), .B(n2694), .C(
        \registers[12][0] ), .D(n2691), .E(n839), .Z(n838) );
  HS65_LH_OAI22X6 U1475 ( .A(n2688), .B(n192), .C(n2685), .D(n160), .Z(n839)
         );
  HS65_LH_AOI212X4 U1476 ( .A(\registers[13][1] ), .B(n2694), .C(
        \registers[12][1] ), .D(n2691), .E(n674), .Z(n673) );
  HS65_LH_OAI22X6 U1477 ( .A(n2688), .B(n191), .C(n2685), .D(n159), .Z(n674)
         );
  HS65_LH_AOI212X4 U1478 ( .A(\registers[13][2] ), .B(n2695), .C(
        \registers[12][2] ), .D(n2692), .E(n509), .Z(n508) );
  HS65_LH_OAI22X6 U1479 ( .A(n2689), .B(n190), .C(n2686), .D(n158), .Z(n509)
         );
  HS65_LH_AOI212X4 U1480 ( .A(\registers[13][3] ), .B(n2696), .C(
        \registers[12][3] ), .D(n2692), .E(n464), .Z(n463) );
  HS65_LH_OAI22X6 U1481 ( .A(n2690), .B(n189), .C(n2686), .D(n157), .Z(n464)
         );
  HS65_LH_AOI212X4 U1482 ( .A(\registers[13][4] ), .B(n2696), .C(
        \registers[12][4] ), .D(n2693), .E(n449), .Z(n448) );
  HS65_LH_OAI22X6 U1483 ( .A(n2690), .B(n188), .C(n2687), .D(n156), .Z(n449)
         );
  HS65_LH_AOI212X4 U1484 ( .A(\registers[13][5] ), .B(n2696), .C(
        \registers[12][5] ), .D(n2693), .E(n434), .Z(n433) );
  HS65_LH_OAI22X6 U1485 ( .A(n2690), .B(n187), .C(n2687), .D(n155), .Z(n434)
         );
  HS65_LH_AOI212X4 U1486 ( .A(\registers[13][6] ), .B(n2696), .C(
        \registers[12][6] ), .D(n2693), .E(n419), .Z(n418) );
  HS65_LH_OAI22X6 U1487 ( .A(n2690), .B(n186), .C(n2687), .D(n154), .Z(n419)
         );
  HS65_LH_AOI212X4 U1488 ( .A(\registers[13][7] ), .B(n2696), .C(
        \registers[12][7] ), .D(n2693), .E(n404), .Z(n403) );
  HS65_LH_OAI22X6 U1489 ( .A(n2690), .B(n185), .C(n2687), .D(n153), .Z(n404)
         );
  HS65_LH_AOI212X4 U1490 ( .A(\registers[13][8] ), .B(n2696), .C(
        \registers[12][8] ), .D(n2693), .E(n389), .Z(n388) );
  HS65_LH_OAI22X6 U1491 ( .A(n2690), .B(n184), .C(n2687), .D(n152), .Z(n389)
         );
  HS65_LH_AOI212X4 U1492 ( .A(\registers[13][9] ), .B(n2696), .C(
        \registers[12][9] ), .D(n2693), .E(n344), .Z(n341) );
  HS65_LH_OAI22X6 U1493 ( .A(n2690), .B(n183), .C(n2687), .D(n151), .Z(n344)
         );
  HS65_LH_AOI212X4 U1494 ( .A(\registers[13][11] ), .B(n2694), .C(
        \registers[12][11] ), .D(n2691), .E(n809), .Z(n808) );
  HS65_LH_OAI22X6 U1495 ( .A(n2688), .B(n181), .C(n2685), .D(n149), .Z(n809)
         );
  HS65_LH_AOI212X4 U1496 ( .A(\registers[13][12] ), .B(n2694), .C(
        \registers[12][12] ), .D(n2691), .E(n794), .Z(n793) );
  HS65_LH_OAI22X6 U1497 ( .A(n2688), .B(n180), .C(n2685), .D(n148), .Z(n794)
         );
  HS65_LH_AOI212X4 U1498 ( .A(\registers[13][13] ), .B(n2694), .C(
        \registers[12][13] ), .D(n2691), .E(n779), .Z(n778) );
  HS65_LH_OAI22X6 U1499 ( .A(n2688), .B(n179), .C(n2685), .D(n147), .Z(n779)
         );
  HS65_LH_AOI212X4 U1500 ( .A(\registers[13][14] ), .B(n2694), .C(
        \registers[12][14] ), .D(n2691), .E(n764), .Z(n763) );
  HS65_LH_OAI22X6 U1501 ( .A(n2688), .B(n178), .C(n2685), .D(n146), .Z(n764)
         );
  HS65_LH_AOI212X4 U1502 ( .A(\registers[13][15] ), .B(n2694), .C(
        \registers[12][15] ), .D(n2691), .E(n749), .Z(n748) );
  HS65_LH_OAI22X6 U1503 ( .A(n2688), .B(n177), .C(n2685), .D(n145), .Z(n749)
         );
  HS65_LH_AOI212X4 U1504 ( .A(\registers[13][16] ), .B(n2694), .C(
        \registers[12][16] ), .D(n2691), .E(n734), .Z(n733) );
  HS65_LH_OAI22X6 U1505 ( .A(n2688), .B(n176), .C(n2685), .D(n144), .Z(n734)
         );
  HS65_LH_AOI212X4 U1506 ( .A(\registers[13][17] ), .B(n2694), .C(
        \registers[12][17] ), .D(n2691), .E(n719), .Z(n718) );
  HS65_LH_OAI22X6 U1507 ( .A(n2688), .B(n175), .C(n2685), .D(n143), .Z(n719)
         );
  HS65_LH_AOI212X4 U1508 ( .A(\registers[13][18] ), .B(n2694), .C(
        \registers[12][18] ), .D(n2691), .E(n704), .Z(n703) );
  HS65_LH_OAI22X6 U1509 ( .A(n2688), .B(n174), .C(n2685), .D(n142), .Z(n704)
         );
  HS65_LH_AOI212X4 U1510 ( .A(\registers[13][19] ), .B(n2694), .C(
        \registers[12][19] ), .D(n2691), .E(n689), .Z(n688) );
  HS65_LH_OAI22X6 U1511 ( .A(n2688), .B(n173), .C(n2685), .D(n141), .Z(n689)
         );
  HS65_LH_AOI212X4 U1512 ( .A(\registers[13][20] ), .B(n2695), .C(
        \registers[12][20] ), .D(n2691), .E(n659), .Z(n658) );
  HS65_LH_OAI22X6 U1513 ( .A(n2689), .B(n172), .C(n2685), .D(n140), .Z(n659)
         );
  HS65_LH_AOI212X4 U1514 ( .A(\registers[13][21] ), .B(n2695), .C(
        \registers[12][21] ), .D(n2692), .E(n644), .Z(n643) );
  HS65_LH_OAI22X6 U1515 ( .A(n2689), .B(n171), .C(n2686), .D(n139), .Z(n644)
         );
  HS65_LH_AOI212X4 U1516 ( .A(\registers[13][22] ), .B(n2695), .C(
        \registers[12][22] ), .D(n2692), .E(n629), .Z(n628) );
  HS65_LH_OAI22X6 U1517 ( .A(n2689), .B(n170), .C(n2686), .D(n138), .Z(n629)
         );
  HS65_LH_AOI212X4 U1518 ( .A(\registers[13][23] ), .B(n2695), .C(
        \registers[12][23] ), .D(n2692), .E(n614), .Z(n613) );
  HS65_LH_OAI22X6 U1519 ( .A(n2689), .B(n169), .C(n2686), .D(n137), .Z(n614)
         );
  HS65_LH_AOI212X4 U1520 ( .A(\registers[13][24] ), .B(n2695), .C(
        \registers[12][24] ), .D(n2692), .E(n599), .Z(n598) );
  HS65_LH_OAI22X6 U1521 ( .A(n2689), .B(n168), .C(n2686), .D(n136), .Z(n599)
         );
  HS65_LH_AOI212X4 U1522 ( .A(\registers[13][25] ), .B(n2695), .C(
        \registers[12][25] ), .D(n2692), .E(n584), .Z(n583) );
  HS65_LH_OAI22X6 U1523 ( .A(n2689), .B(n167), .C(n2686), .D(n135), .Z(n584)
         );
  HS65_LH_AOI212X4 U1524 ( .A(\registers[13][26] ), .B(n2695), .C(
        \registers[12][26] ), .D(n2692), .E(n569), .Z(n568) );
  HS65_LH_OAI22X6 U1525 ( .A(n2689), .B(n166), .C(n2686), .D(n134), .Z(n569)
         );
  HS65_LH_AOI212X4 U1526 ( .A(\registers[13][27] ), .B(n2695), .C(
        \registers[12][27] ), .D(n2692), .E(n554), .Z(n553) );
  HS65_LH_OAI22X6 U1527 ( .A(n2689), .B(n165), .C(n2686), .D(n133), .Z(n554)
         );
  HS65_LH_AOI212X4 U1528 ( .A(\registers[13][28] ), .B(n2695), .C(
        \registers[12][28] ), .D(n2692), .E(n539), .Z(n538) );
  HS65_LH_OAI22X6 U1529 ( .A(n2689), .B(n164), .C(n2686), .D(n132), .Z(n539)
         );
  HS65_LH_AOI212X4 U1530 ( .A(\registers[13][29] ), .B(n2695), .C(
        \registers[12][29] ), .D(n2692), .E(n524), .Z(n523) );
  HS65_LH_OAI22X6 U1531 ( .A(n2689), .B(n163), .C(n2686), .D(n131), .Z(n524)
         );
  HS65_LH_AOI212X4 U1532 ( .A(\registers[13][30] ), .B(n2695), .C(
        \registers[12][30] ), .D(n2692), .E(n494), .Z(n493) );
  HS65_LH_OAI22X6 U1533 ( .A(n2689), .B(n162), .C(n2686), .D(n130), .Z(n494)
         );
  HS65_LH_AOI212X4 U1534 ( .A(\registers[13][31] ), .B(n2696), .C(
        \registers[12][31] ), .D(n2692), .E(n479), .Z(n478) );
  HS65_LH_OAI22X6 U1535 ( .A(n2690), .B(n161), .C(n2686), .D(n129), .Z(n479)
         );
  HS65_LH_AOI212X4 U1536 ( .A(n2603), .B(\registers[13][4] ), .C(n2600), .D(
        \registers[12][4] ), .E(n977), .Z(n976) );
  HS65_LH_OAI22X6 U1537 ( .A(n188), .B(n2597), .C(n156), .D(n2594), .Z(n977)
         );
  HS65_LH_AOI212X4 U1538 ( .A(n2603), .B(\registers[13][5] ), .C(n2600), .D(
        \registers[12][5] ), .E(n962), .Z(n961) );
  HS65_LH_OAI22X6 U1539 ( .A(n187), .B(n2597), .C(n155), .D(n2594), .Z(n962)
         );
  HS65_LH_AOI212X4 U1540 ( .A(n2603), .B(\registers[13][6] ), .C(n2600), .D(
        \registers[12][6] ), .E(n947), .Z(n946) );
  HS65_LH_OAI22X6 U1541 ( .A(n186), .B(n2597), .C(n154), .D(n2594), .Z(n947)
         );
  HS65_LH_AOI212X4 U1542 ( .A(n2603), .B(\registers[13][7] ), .C(n2600), .D(
        \registers[12][7] ), .E(n932), .Z(n931) );
  HS65_LH_OAI22X6 U1543 ( .A(n185), .B(n2597), .C(n153), .D(n2594), .Z(n932)
         );
  HS65_LH_AOI212X4 U1544 ( .A(n2603), .B(\registers[13][8] ), .C(n2600), .D(
        \registers[12][8] ), .E(n917), .Z(n916) );
  HS65_LH_OAI22X6 U1545 ( .A(n184), .B(n2597), .C(n152), .D(n2594), .Z(n917)
         );
  HS65_LH_AOI212X4 U1546 ( .A(n2603), .B(\registers[13][9] ), .C(n2600), .D(
        \registers[12][9] ), .E(n872), .Z(n869) );
  HS65_LH_OAI22X6 U1547 ( .A(n183), .B(n2597), .C(n151), .D(n2594), .Z(n872)
         );
  HS65_LH_OAI22X6 U1548 ( .A(n2643), .B(n64), .C(n2640), .D(n32), .Z(n855) );
  HS65_LH_OAI22X6 U1549 ( .A(n2643), .B(n63), .C(n2640), .D(n31), .Z(n680) );
  HS65_LH_OAI22X6 U1550 ( .A(n2644), .B(n62), .C(n2641), .D(n30), .Z(n515) );
  HS65_LH_OAI22X6 U1551 ( .A(n2633), .B(n125), .C(n2629), .D(n93), .Z(n471) );
  HS65_LH_OAI22X6 U1552 ( .A(n2645), .B(n61), .C(n2641), .D(n29), .Z(n470) );
  HS65_LH_OAI22X6 U1553 ( .A(n2633), .B(n124), .C(n2630), .D(n92), .Z(n456) );
  HS65_LH_OAI22X6 U1554 ( .A(n2645), .B(n60), .C(n2642), .D(n28), .Z(n455) );
  HS65_LH_OAI22X6 U1555 ( .A(n2633), .B(n123), .C(n2630), .D(n91), .Z(n441) );
  HS65_LH_OAI22X6 U1556 ( .A(n2645), .B(n59), .C(n2642), .D(n27), .Z(n440) );
  HS65_LH_OAI22X6 U1557 ( .A(n2633), .B(n122), .C(n2630), .D(n90), .Z(n426) );
  HS65_LH_OAI22X6 U1558 ( .A(n2645), .B(n58), .C(n2642), .D(n26), .Z(n425) );
  HS65_LH_OAI22X6 U1559 ( .A(n2633), .B(n121), .C(n2630), .D(n89), .Z(n411) );
  HS65_LH_OAI22X6 U1560 ( .A(n2645), .B(n57), .C(n2642), .D(n25), .Z(n410) );
  HS65_LH_OAI22X6 U1561 ( .A(n2633), .B(n120), .C(n2630), .D(n88), .Z(n396) );
  HS65_LH_OAI22X6 U1562 ( .A(n2645), .B(n56), .C(n2642), .D(n24), .Z(n395) );
  HS65_LH_OAI22X6 U1563 ( .A(n2633), .B(n119), .C(n2630), .D(n87), .Z(n371) );
  HS65_LH_OAI22X6 U1564 ( .A(n2645), .B(n55), .C(n2642), .D(n23), .Z(n366) );
  HS65_LH_OAI22X6 U1565 ( .A(n2643), .B(n54), .C(n2640), .D(n22), .Z(n830) );
  HS65_LH_OAI22X6 U1566 ( .A(n2676), .B(n246), .C(n2673), .D(n214), .Z(n825)
         );
  HS65_LH_OAI22X6 U1567 ( .A(n2688), .B(n182), .C(n2685), .D(n150), .Z(n824)
         );
  HS65_LH_OAI22X6 U1568 ( .A(n2643), .B(n53), .C(n2640), .D(n21), .Z(n815) );
  HS65_LH_OAI22X6 U1569 ( .A(n2643), .B(n52), .C(n2640), .D(n20), .Z(n800) );
  HS65_LH_OAI22X6 U1570 ( .A(n2643), .B(n51), .C(n2640), .D(n19), .Z(n785) );
  HS65_LH_OAI22X6 U1571 ( .A(n2643), .B(n50), .C(n2640), .D(n18), .Z(n770) );
  HS65_LH_OAI22X6 U1572 ( .A(n2643), .B(n49), .C(n2640), .D(n17), .Z(n755) );
  HS65_LH_OAI22X6 U1573 ( .A(n2643), .B(n48), .C(n2640), .D(n16), .Z(n740) );
  HS65_LH_OAI22X6 U1574 ( .A(n2643), .B(n47), .C(n2640), .D(n15), .Z(n725) );
  HS65_LH_OAI22X6 U1575 ( .A(n2643), .B(n46), .C(n2640), .D(n14), .Z(n710) );
  HS65_LH_OAI22X6 U1576 ( .A(n2643), .B(n45), .C(n2640), .D(n13), .Z(n695) );
  HS65_LH_OAI22X6 U1577 ( .A(n2644), .B(n44), .C(n2640), .D(n12), .Z(n665) );
  HS65_LH_OAI22X6 U1578 ( .A(n2644), .B(n43), .C(n2641), .D(n11), .Z(n650) );
  HS65_LH_OAI22X6 U1579 ( .A(n2644), .B(n42), .C(n2641), .D(n10), .Z(n635) );
  HS65_LH_OAI22X6 U1580 ( .A(n2644), .B(n41), .C(n2641), .D(n9), .Z(n620) );
  HS65_LH_OAI22X6 U1581 ( .A(n2644), .B(n40), .C(n2641), .D(n8), .Z(n605) );
  HS65_LH_OAI22X6 U1582 ( .A(n2644), .B(n39), .C(n2641), .D(n7), .Z(n590) );
  HS65_LH_OAI22X6 U1583 ( .A(n2644), .B(n38), .C(n2641), .D(n6), .Z(n575) );
  HS65_LH_OAI22X6 U1584 ( .A(n2644), .B(n37), .C(n2641), .D(n5), .Z(n560) );
  HS65_LH_OAI22X6 U1585 ( .A(n2644), .B(n36), .C(n2641), .D(n4), .Z(n545) );
  HS65_LH_OAI22X6 U1586 ( .A(n2644), .B(n35), .C(n2641), .D(n3), .Z(n530) );
  HS65_LH_OAI22X6 U1587 ( .A(n2644), .B(n34), .C(n2641), .D(n2), .Z(n500) );
  HS65_LH_OAI22X6 U1588 ( .A(n2633), .B(n97), .C(n2629), .D(n65), .Z(n486) );
  HS65_LH_OAI22X6 U1589 ( .A(n2645), .B(n33), .C(n2641), .D(n1), .Z(n485) );
  HS65_LH_OAI22X6 U1590 ( .A(n128), .B(n2538), .C(n96), .D(n2535), .Z(n1386)
         );
  HS65_LH_OAI22X6 U1591 ( .A(n64), .B(n2550), .C(n32), .D(n2547), .Z(n1383) );
  HS65_LH_OAI22X6 U1592 ( .A(n127), .B(n2538), .C(n95), .D(n2535), .Z(n1209)
         );
  HS65_LH_OAI22X6 U1593 ( .A(n63), .B(n2550), .C(n31), .D(n2547), .Z(n1208) );
  HS65_LH_OAI22X6 U1594 ( .A(n126), .B(n2539), .C(n94), .D(n2536), .Z(n1044)
         );
  HS65_LH_OAI22X6 U1595 ( .A(n62), .B(n2551), .C(n30), .D(n2548), .Z(n1043) );
  HS65_LH_OAI22X6 U1596 ( .A(n118), .B(n2538), .C(n86), .D(n2535), .Z(n1359)
         );
  HS65_LH_OAI22X6 U1597 ( .A(n54), .B(n2550), .C(n22), .D(n2547), .Z(n1358) );
  HS65_LH_OAI22X6 U1598 ( .A(n117), .B(n2538), .C(n85), .D(n2535), .Z(n1344)
         );
  HS65_LH_OAI22X6 U1599 ( .A(n53), .B(n2550), .C(n21), .D(n2547), .Z(n1343) );
  HS65_LH_OAI22X6 U1600 ( .A(n116), .B(n2538), .C(n84), .D(n2535), .Z(n1329)
         );
  HS65_LH_OAI22X6 U1601 ( .A(n52), .B(n2550), .C(n20), .D(n2547), .Z(n1328) );
  HS65_LH_OAI22X6 U1602 ( .A(n115), .B(n2538), .C(n83), .D(n2535), .Z(n1314)
         );
  HS65_LH_OAI22X6 U1603 ( .A(n51), .B(n2550), .C(n19), .D(n2547), .Z(n1313) );
  HS65_LH_OAI22X6 U1604 ( .A(n114), .B(n2538), .C(n82), .D(n2535), .Z(n1299)
         );
  HS65_LH_OAI22X6 U1605 ( .A(n50), .B(n2550), .C(n18), .D(n2547), .Z(n1298) );
  HS65_LH_OAI22X6 U1606 ( .A(n113), .B(n2538), .C(n81), .D(n2535), .Z(n1284)
         );
  HS65_LH_OAI22X6 U1607 ( .A(n49), .B(n2550), .C(n17), .D(n2547), .Z(n1283) );
  HS65_LH_OAI22X6 U1608 ( .A(n112), .B(n2538), .C(n80), .D(n2535), .Z(n1269)
         );
  HS65_LH_OAI22X6 U1609 ( .A(n48), .B(n2550), .C(n16), .D(n2547), .Z(n1268) );
  HS65_LH_OAI22X6 U1610 ( .A(n111), .B(n2538), .C(n79), .D(n2535), .Z(n1254)
         );
  HS65_LH_OAI22X6 U1611 ( .A(n47), .B(n2550), .C(n15), .D(n2547), .Z(n1253) );
  HS65_LH_OAI22X6 U1612 ( .A(n110), .B(n2538), .C(n78), .D(n2535), .Z(n1239)
         );
  HS65_LH_OAI22X6 U1613 ( .A(n46), .B(n2550), .C(n14), .D(n2547), .Z(n1238) );
  HS65_LH_OAI22X6 U1614 ( .A(n109), .B(n2538), .C(n77), .D(n2535), .Z(n1224)
         );
  HS65_LH_OAI22X6 U1615 ( .A(n45), .B(n2550), .C(n13), .D(n2547), .Z(n1223) );
  HS65_LH_OAI22X6 U1616 ( .A(n108), .B(n2539), .C(n76), .D(n2535), .Z(n1194)
         );
  HS65_LH_OAI22X6 U1617 ( .A(n44), .B(n2551), .C(n12), .D(n2547), .Z(n1193) );
  HS65_LH_OAI22X6 U1618 ( .A(n107), .B(n2539), .C(n75), .D(n2536), .Z(n1179)
         );
  HS65_LH_OAI22X6 U1619 ( .A(n43), .B(n2551), .C(n11), .D(n2548), .Z(n1178) );
  HS65_LH_OAI22X6 U1620 ( .A(n106), .B(n2539), .C(n74), .D(n2536), .Z(n1164)
         );
  HS65_LH_OAI22X6 U1621 ( .A(n42), .B(n2551), .C(n10), .D(n2548), .Z(n1163) );
  HS65_LH_OAI22X6 U1622 ( .A(n105), .B(n2539), .C(n73), .D(n2536), .Z(n1149)
         );
  HS65_LH_OAI22X6 U1623 ( .A(n41), .B(n2551), .C(n9), .D(n2548), .Z(n1148) );
  HS65_LH_OAI22X6 U1624 ( .A(n104), .B(n2539), .C(n72), .D(n2536), .Z(n1134)
         );
  HS65_LH_OAI22X6 U1625 ( .A(n40), .B(n2551), .C(n8), .D(n2548), .Z(n1133) );
  HS65_LH_OAI22X6 U1626 ( .A(n103), .B(n2539), .C(n71), .D(n2536), .Z(n1119)
         );
  HS65_LH_OAI22X6 U1627 ( .A(n39), .B(n2551), .C(n7), .D(n2548), .Z(n1118) );
  HS65_LH_OAI22X6 U1628 ( .A(n102), .B(n2539), .C(n70), .D(n2536), .Z(n1104)
         );
  HS65_LH_OAI22X6 U1629 ( .A(n38), .B(n2551), .C(n6), .D(n2548), .Z(n1103) );
  HS65_LH_OAI22X6 U1630 ( .A(n101), .B(n2539), .C(n69), .D(n2536), .Z(n1089)
         );
  HS65_LH_OAI22X6 U1631 ( .A(n37), .B(n2551), .C(n5), .D(n2548), .Z(n1088) );
  HS65_LH_OAI22X6 U1632 ( .A(n100), .B(n2539), .C(n68), .D(n2536), .Z(n1074)
         );
  HS65_LH_OAI22X6 U1633 ( .A(n36), .B(n2551), .C(n4), .D(n2548), .Z(n1073) );
  HS65_LH_OAI22X6 U1634 ( .A(n99), .B(n2539), .C(n67), .D(n2536), .Z(n1059) );
  HS65_LH_OAI22X6 U1635 ( .A(n35), .B(n2551), .C(n3), .D(n2548), .Z(n1058) );
  HS65_LH_OAI22X6 U1636 ( .A(n98), .B(n2539), .C(n66), .D(n2536), .Z(n1029) );
  HS65_LH_OAI22X6 U1637 ( .A(n34), .B(n2551), .C(n2), .D(n2548), .Z(n1028) );
  HS65_LH_OAI22X6 U1638 ( .A(n125), .B(n2540), .C(n93), .D(n2536), .Z(n999) );
  HS65_LH_OAI22X6 U1639 ( .A(n61), .B(n2552), .C(n29), .D(n2548), .Z(n998) );
  HS65_LH_OAI22X6 U1640 ( .A(n124), .B(n2540), .C(n92), .D(n2537), .Z(n984) );
  HS65_LH_OAI22X6 U1641 ( .A(n60), .B(n2552), .C(n28), .D(n2549), .Z(n983) );
  HS65_LH_OAI22X6 U1642 ( .A(n123), .B(n2540), .C(n91), .D(n2537), .Z(n969) );
  HS65_LH_OAI22X6 U1643 ( .A(n59), .B(n2552), .C(n27), .D(n2549), .Z(n968) );
  HS65_LH_OAI22X6 U1644 ( .A(n122), .B(n2540), .C(n90), .D(n2537), .Z(n954) );
  HS65_LH_OAI22X6 U1645 ( .A(n58), .B(n2552), .C(n26), .D(n2549), .Z(n953) );
  HS65_LH_OAI22X6 U1646 ( .A(n121), .B(n2540), .C(n89), .D(n2537), .Z(n939) );
  HS65_LH_OAI22X6 U1647 ( .A(n57), .B(n2552), .C(n25), .D(n2549), .Z(n938) );
  HS65_LH_OAI22X6 U1648 ( .A(n120), .B(n2540), .C(n88), .D(n2537), .Z(n924) );
  HS65_LH_OAI22X6 U1649 ( .A(n56), .B(n2552), .C(n24), .D(n2549), .Z(n923) );
  HS65_LH_OAI22X6 U1650 ( .A(n119), .B(n2540), .C(n87), .D(n2537), .Z(n899) );
  HS65_LH_OAI22X6 U1651 ( .A(n55), .B(n2552), .C(n23), .D(n2549), .Z(n894) );
  HS65_LH_OAI22X6 U1652 ( .A(n97), .B(n2540), .C(n65), .D(n2536), .Z(n1014) );
  HS65_LH_OAI22X6 U1653 ( .A(n33), .B(n2552), .C(n1), .D(n2548), .Z(n1013) );
  HS65_LH_OAI22X6 U1654 ( .A(n2760), .B(n2473), .C(n2471), .D(n225), .Z(n1689)
         );
  HS65_LH_OAI22X6 U1655 ( .A(n2760), .B(n2468), .C(n2466), .D(n193), .Z(n1721)
         );
  HS65_LH_OAI22X6 U1656 ( .A(n2760), .B(n2443), .C(n2441), .D(n161), .Z(n1881)
         );
  HS65_LH_OAI22X6 U1657 ( .A(n2760), .B(n2438), .C(n2436), .D(n129), .Z(n1913)
         );
  HS65_LH_OAI22X6 U1658 ( .A(n2760), .B(n305), .C(n303), .D(n33), .Z(n2329) );
  HS65_LH_OAI22X6 U1659 ( .A(n2760), .B(n300), .C(n298), .D(n1), .Z(n2361) );
  HS65_LH_OAI22X6 U1660 ( .A(n2760), .B(n315), .C(n313), .D(n97), .Z(n2265) );
  HS65_LH_OAI22X6 U1661 ( .A(n2760), .B(n310), .C(n308), .D(n65), .Z(n2297) );
  HS65_LH_OAI22X6 U1662 ( .A(n2724), .B(n2474), .C(n2472), .D(n243), .Z(n1671)
         );
  HS65_LH_OAI22X6 U1663 ( .A(n2726), .B(n2474), .C(n2472), .D(n242), .Z(n1672)
         );
  HS65_LH_OAI22X6 U1664 ( .A(n2728), .B(n2474), .C(n2472), .D(n241), .Z(n1673)
         );
  HS65_LH_OAI22X6 U1665 ( .A(n2730), .B(n2474), .C(n2472), .D(n240), .Z(n1674)
         );
  HS65_LH_OAI22X6 U1666 ( .A(n2732), .B(n2474), .C(n2472), .D(n239), .Z(n1675)
         );
  HS65_LH_OAI22X6 U1667 ( .A(n2734), .B(n2474), .C(n2472), .D(n238), .Z(n1676)
         );
  HS65_LH_OAI22X6 U1668 ( .A(n2736), .B(n2474), .C(n2471), .D(n237), .Z(n1677)
         );
  HS65_LH_OAI22X6 U1669 ( .A(n2738), .B(n2474), .C(n2471), .D(n236), .Z(n1678)
         );
  HS65_LH_OAI22X6 U1670 ( .A(n2740), .B(n2474), .C(n2471), .D(n235), .Z(n1679)
         );
  HS65_LH_OAI22X6 U1671 ( .A(n2742), .B(n2474), .C(n2471), .D(n234), .Z(n1680)
         );
  HS65_LH_OAI22X6 U1672 ( .A(n2744), .B(n2474), .C(n2471), .D(n233), .Z(n1681)
         );
  HS65_LH_OAI22X6 U1673 ( .A(n2746), .B(n2474), .C(n2471), .D(n232), .Z(n1682)
         );
  HS65_LH_OAI22X6 U1674 ( .A(n2748), .B(n2474), .C(n2471), .D(n231), .Z(n1683)
         );
  HS65_LH_OAI22X6 U1675 ( .A(n2750), .B(n2474), .C(n2471), .D(n230), .Z(n1684)
         );
  HS65_LH_OAI22X6 U1676 ( .A(n2752), .B(n2474), .C(n2471), .D(n229), .Z(n1685)
         );
  HS65_LH_OAI22X6 U1677 ( .A(n2754), .B(n2474), .C(n2471), .D(n228), .Z(n1686)
         );
  HS65_LH_OAI22X6 U1678 ( .A(n2756), .B(n2474), .C(n2471), .D(n227), .Z(n1687)
         );
  HS65_LH_OAI22X6 U1679 ( .A(n2758), .B(n2474), .C(n2471), .D(n226), .Z(n1688)
         );
  HS65_LH_OAI22X6 U1680 ( .A(n2724), .B(n2469), .C(n2467), .D(n211), .Z(n1703)
         );
  HS65_LH_OAI22X6 U1681 ( .A(n2726), .B(n2469), .C(n2467), .D(n210), .Z(n1704)
         );
  HS65_LH_OAI22X6 U1682 ( .A(n2728), .B(n2469), .C(n2467), .D(n209), .Z(n1705)
         );
  HS65_LH_OAI22X6 U1683 ( .A(n2730), .B(n2469), .C(n2467), .D(n208), .Z(n1706)
         );
  HS65_LH_OAI22X6 U1684 ( .A(n2732), .B(n2469), .C(n2467), .D(n207), .Z(n1707)
         );
  HS65_LH_OAI22X6 U1685 ( .A(n2734), .B(n2469), .C(n2467), .D(n206), .Z(n1708)
         );
  HS65_LH_OAI22X6 U1686 ( .A(n2736), .B(n2469), .C(n2466), .D(n205), .Z(n1709)
         );
  HS65_LH_OAI22X6 U1687 ( .A(n2738), .B(n2469), .C(n2466), .D(n204), .Z(n1710)
         );
  HS65_LH_OAI22X6 U1688 ( .A(n2740), .B(n2469), .C(n2466), .D(n203), .Z(n1711)
         );
  HS65_LH_OAI22X6 U1689 ( .A(n2742), .B(n2469), .C(n2466), .D(n202), .Z(n1712)
         );
  HS65_LH_OAI22X6 U1690 ( .A(n2744), .B(n2469), .C(n2466), .D(n201), .Z(n1713)
         );
  HS65_LH_OAI22X6 U1691 ( .A(n2746), .B(n2469), .C(n2466), .D(n200), .Z(n1714)
         );
  HS65_LH_OAI22X6 U1692 ( .A(n2748), .B(n2469), .C(n2466), .D(n199), .Z(n1715)
         );
  HS65_LH_OAI22X6 U1693 ( .A(n2750), .B(n2469), .C(n2466), .D(n198), .Z(n1716)
         );
  HS65_LH_OAI22X6 U1694 ( .A(n2752), .B(n2469), .C(n2466), .D(n197), .Z(n1717)
         );
  HS65_LH_OAI22X6 U1695 ( .A(n2754), .B(n2469), .C(n2466), .D(n196), .Z(n1718)
         );
  HS65_LH_OAI22X6 U1696 ( .A(n2756), .B(n2469), .C(n2466), .D(n195), .Z(n1719)
         );
  HS65_LH_OAI22X6 U1697 ( .A(n2758), .B(n2469), .C(n2466), .D(n194), .Z(n1720)
         );
  HS65_LH_OAI22X6 U1698 ( .A(n2724), .B(n2444), .C(n2442), .D(n179), .Z(n1863)
         );
  HS65_LH_OAI22X6 U1699 ( .A(n2726), .B(n2444), .C(n2442), .D(n178), .Z(n1864)
         );
  HS65_LH_OAI22X6 U1700 ( .A(n2728), .B(n2444), .C(n2442), .D(n177), .Z(n1865)
         );
  HS65_LH_OAI22X6 U1701 ( .A(n2730), .B(n2444), .C(n2442), .D(n176), .Z(n1866)
         );
  HS65_LH_OAI22X6 U1702 ( .A(n2732), .B(n2444), .C(n2442), .D(n175), .Z(n1867)
         );
  HS65_LH_OAI22X6 U1703 ( .A(n2734), .B(n2444), .C(n2442), .D(n174), .Z(n1868)
         );
  HS65_LH_OAI22X6 U1704 ( .A(n2736), .B(n2444), .C(n2441), .D(n173), .Z(n1869)
         );
  HS65_LH_OAI22X6 U1705 ( .A(n2738), .B(n2444), .C(n2441), .D(n172), .Z(n1870)
         );
  HS65_LH_OAI22X6 U1706 ( .A(n2740), .B(n2444), .C(n2441), .D(n171), .Z(n1871)
         );
  HS65_LH_OAI22X6 U1707 ( .A(n2742), .B(n2444), .C(n2441), .D(n170), .Z(n1872)
         );
  HS65_LH_OAI22X6 U1708 ( .A(n2744), .B(n2444), .C(n2441), .D(n169), .Z(n1873)
         );
  HS65_LH_OAI22X6 U1709 ( .A(n2746), .B(n2444), .C(n2441), .D(n168), .Z(n1874)
         );
  HS65_LH_OAI22X6 U1710 ( .A(n2748), .B(n2444), .C(n2441), .D(n167), .Z(n1875)
         );
  HS65_LH_OAI22X6 U1711 ( .A(n2750), .B(n2444), .C(n2441), .D(n166), .Z(n1876)
         );
  HS65_LH_OAI22X6 U1712 ( .A(n2752), .B(n2444), .C(n2441), .D(n165), .Z(n1877)
         );
  HS65_LH_OAI22X6 U1713 ( .A(n2754), .B(n2444), .C(n2441), .D(n164), .Z(n1878)
         );
  HS65_LH_OAI22X6 U1714 ( .A(n2756), .B(n2444), .C(n2441), .D(n163), .Z(n1879)
         );
  HS65_LH_OAI22X6 U1715 ( .A(n2758), .B(n2444), .C(n2441), .D(n162), .Z(n1880)
         );
  HS65_LH_OAI22X6 U1716 ( .A(n2724), .B(n2439), .C(n2437), .D(n147), .Z(n1895)
         );
  HS65_LH_OAI22X6 U1717 ( .A(n2726), .B(n2439), .C(n2437), .D(n146), .Z(n1896)
         );
  HS65_LH_OAI22X6 U1718 ( .A(n2728), .B(n2439), .C(n2437), .D(n145), .Z(n1897)
         );
  HS65_LH_OAI22X6 U1719 ( .A(n2730), .B(n2439), .C(n2437), .D(n144), .Z(n1898)
         );
  HS65_LH_OAI22X6 U1720 ( .A(n2732), .B(n2439), .C(n2437), .D(n143), .Z(n1899)
         );
  HS65_LH_OAI22X6 U1721 ( .A(n2734), .B(n2439), .C(n2437), .D(n142), .Z(n1900)
         );
  HS65_LH_OAI22X6 U1722 ( .A(n2736), .B(n2439), .C(n2436), .D(n141), .Z(n1901)
         );
  HS65_LH_OAI22X6 U1723 ( .A(n2738), .B(n2439), .C(n2436), .D(n140), .Z(n1902)
         );
  HS65_LH_OAI22X6 U1724 ( .A(n2740), .B(n2439), .C(n2436), .D(n139), .Z(n1903)
         );
  HS65_LH_OAI22X6 U1725 ( .A(n2742), .B(n2439), .C(n2436), .D(n138), .Z(n1904)
         );
  HS65_LH_OAI22X6 U1726 ( .A(n2744), .B(n2439), .C(n2436), .D(n137), .Z(n1905)
         );
  HS65_LH_OAI22X6 U1727 ( .A(n2746), .B(n2439), .C(n2436), .D(n136), .Z(n1906)
         );
  HS65_LH_OAI22X6 U1728 ( .A(n2748), .B(n2439), .C(n2436), .D(n135), .Z(n1907)
         );
  HS65_LH_OAI22X6 U1729 ( .A(n2750), .B(n2439), .C(n2436), .D(n134), .Z(n1908)
         );
  HS65_LH_OAI22X6 U1730 ( .A(n2752), .B(n2439), .C(n2436), .D(n133), .Z(n1909)
         );
  HS65_LH_OAI22X6 U1731 ( .A(n2754), .B(n2439), .C(n2436), .D(n132), .Z(n1910)
         );
  HS65_LH_OAI22X6 U1732 ( .A(n2756), .B(n2439), .C(n2436), .D(n131), .Z(n1911)
         );
  HS65_LH_OAI22X6 U1733 ( .A(n2758), .B(n2439), .C(n2436), .D(n130), .Z(n1912)
         );
  HS65_LH_OAI22X6 U1734 ( .A(n2724), .B(n306), .C(n304), .D(n51), .Z(n2311) );
  HS65_LH_OAI22X6 U1735 ( .A(n2726), .B(n306), .C(n304), .D(n50), .Z(n2312) );
  HS65_LH_OAI22X6 U1736 ( .A(n2728), .B(n306), .C(n304), .D(n49), .Z(n2313) );
  HS65_LH_OAI22X6 U1737 ( .A(n2730), .B(n306), .C(n304), .D(n48), .Z(n2314) );
  HS65_LH_OAI22X6 U1738 ( .A(n2732), .B(n306), .C(n304), .D(n47), .Z(n2315) );
  HS65_LH_OAI22X6 U1739 ( .A(n2734), .B(n306), .C(n304), .D(n46), .Z(n2316) );
  HS65_LH_OAI22X6 U1740 ( .A(n2736), .B(n306), .C(n303), .D(n45), .Z(n2317) );
  HS65_LH_OAI22X6 U1741 ( .A(n2738), .B(n306), .C(n303), .D(n44), .Z(n2318) );
  HS65_LH_OAI22X6 U1742 ( .A(n2740), .B(n306), .C(n303), .D(n43), .Z(n2319) );
  HS65_LH_OAI22X6 U1743 ( .A(n2742), .B(n306), .C(n303), .D(n42), .Z(n2320) );
  HS65_LH_OAI22X6 U1744 ( .A(n2744), .B(n306), .C(n303), .D(n41), .Z(n2321) );
  HS65_LH_OAI22X6 U1745 ( .A(n2746), .B(n306), .C(n303), .D(n40), .Z(n2322) );
  HS65_LH_OAI22X6 U1746 ( .A(n2748), .B(n306), .C(n303), .D(n39), .Z(n2323) );
  HS65_LH_OAI22X6 U1747 ( .A(n2750), .B(n306), .C(n303), .D(n38), .Z(n2324) );
  HS65_LH_OAI22X6 U1748 ( .A(n2752), .B(n306), .C(n303), .D(n37), .Z(n2325) );
  HS65_LH_OAI22X6 U1749 ( .A(n2754), .B(n306), .C(n303), .D(n36), .Z(n2326) );
  HS65_LH_OAI22X6 U1750 ( .A(n2756), .B(n306), .C(n303), .D(n35), .Z(n2327) );
  HS65_LH_OAI22X6 U1751 ( .A(n2758), .B(n306), .C(n303), .D(n34), .Z(n2328) );
  HS65_LH_OAI22X6 U1752 ( .A(n2724), .B(n301), .C(n299), .D(n19), .Z(n2343) );
  HS65_LH_OAI22X6 U1753 ( .A(n2726), .B(n301), .C(n299), .D(n18), .Z(n2344) );
  HS65_LH_OAI22X6 U1754 ( .A(n2728), .B(n301), .C(n299), .D(n17), .Z(n2345) );
  HS65_LH_OAI22X6 U1755 ( .A(n2730), .B(n301), .C(n299), .D(n16), .Z(n2346) );
  HS65_LH_OAI22X6 U1756 ( .A(n2732), .B(n301), .C(n299), .D(n15), .Z(n2347) );
  HS65_LH_OAI22X6 U1757 ( .A(n2734), .B(n301), .C(n299), .D(n14), .Z(n2348) );
  HS65_LH_OAI22X6 U1758 ( .A(n2736), .B(n301), .C(n298), .D(n13), .Z(n2349) );
  HS65_LH_OAI22X6 U1759 ( .A(n2738), .B(n301), .C(n298), .D(n12), .Z(n2350) );
  HS65_LH_OAI22X6 U1760 ( .A(n2740), .B(n301), .C(n298), .D(n11), .Z(n2351) );
  HS65_LH_OAI22X6 U1761 ( .A(n2742), .B(n301), .C(n298), .D(n10), .Z(n2352) );
  HS65_LH_OAI22X6 U1762 ( .A(n2744), .B(n301), .C(n298), .D(n9), .Z(n2353) );
  HS65_LH_OAI22X6 U1763 ( .A(n2746), .B(n301), .C(n298), .D(n8), .Z(n2354) );
  HS65_LH_OAI22X6 U1764 ( .A(n2748), .B(n301), .C(n298), .D(n7), .Z(n2355) );
  HS65_LH_OAI22X6 U1765 ( .A(n2750), .B(n301), .C(n298), .D(n6), .Z(n2356) );
  HS65_LH_OAI22X6 U1766 ( .A(n2752), .B(n301), .C(n298), .D(n5), .Z(n2357) );
  HS65_LH_OAI22X6 U1767 ( .A(n2754), .B(n301), .C(n298), .D(n4), .Z(n2358) );
  HS65_LH_OAI22X6 U1768 ( .A(n2756), .B(n301), .C(n298), .D(n3), .Z(n2359) );
  HS65_LH_OAI22X6 U1769 ( .A(n2758), .B(n301), .C(n298), .D(n2), .Z(n2360) );
  HS65_LH_OAI22X6 U1770 ( .A(n2724), .B(n316), .C(n314), .D(n115), .Z(n2247)
         );
  HS65_LH_OAI22X6 U1771 ( .A(n2726), .B(n316), .C(n314), .D(n114), .Z(n2248)
         );
  HS65_LH_OAI22X6 U1772 ( .A(n2728), .B(n316), .C(n314), .D(n113), .Z(n2249)
         );
  HS65_LH_OAI22X6 U1773 ( .A(n2730), .B(n316), .C(n314), .D(n112), .Z(n2250)
         );
  HS65_LH_OAI22X6 U1774 ( .A(n2732), .B(n316), .C(n314), .D(n111), .Z(n2251)
         );
  HS65_LH_OAI22X6 U1775 ( .A(n2734), .B(n316), .C(n314), .D(n110), .Z(n2252)
         );
  HS65_LH_OAI22X6 U1776 ( .A(n2736), .B(n316), .C(n313), .D(n109), .Z(n2253)
         );
  HS65_LH_OAI22X6 U1777 ( .A(n2738), .B(n316), .C(n313), .D(n108), .Z(n2254)
         );
  HS65_LH_OAI22X6 U1778 ( .A(n2740), .B(n316), .C(n313), .D(n107), .Z(n2255)
         );
  HS65_LH_OAI22X6 U1779 ( .A(n2742), .B(n316), .C(n313), .D(n106), .Z(n2256)
         );
  HS65_LH_OAI22X6 U1780 ( .A(n2744), .B(n316), .C(n313), .D(n105), .Z(n2257)
         );
  HS65_LH_OAI22X6 U1781 ( .A(n2746), .B(n316), .C(n313), .D(n104), .Z(n2258)
         );
  HS65_LH_OAI22X6 U1782 ( .A(n2748), .B(n316), .C(n313), .D(n103), .Z(n2259)
         );
  HS65_LH_OAI22X6 U1783 ( .A(n2750), .B(n316), .C(n313), .D(n102), .Z(n2260)
         );
  HS65_LH_OAI22X6 U1784 ( .A(n2752), .B(n316), .C(n313), .D(n101), .Z(n2261)
         );
  HS65_LH_OAI22X6 U1785 ( .A(n2754), .B(n316), .C(n313), .D(n100), .Z(n2262)
         );
  HS65_LH_OAI22X6 U1786 ( .A(n2756), .B(n316), .C(n313), .D(n99), .Z(n2263) );
  HS65_LH_OAI22X6 U1787 ( .A(n2758), .B(n316), .C(n313), .D(n98), .Z(n2264) );
  HS65_LH_OAI22X6 U1788 ( .A(n2724), .B(n311), .C(n309), .D(n83), .Z(n2279) );
  HS65_LH_OAI22X6 U1789 ( .A(n2726), .B(n311), .C(n309), .D(n82), .Z(n2280) );
  HS65_LH_OAI22X6 U1790 ( .A(n2728), .B(n311), .C(n309), .D(n81), .Z(n2281) );
  HS65_LH_OAI22X6 U1791 ( .A(n2730), .B(n311), .C(n309), .D(n80), .Z(n2282) );
  HS65_LH_OAI22X6 U1792 ( .A(n2732), .B(n311), .C(n309), .D(n79), .Z(n2283) );
  HS65_LH_OAI22X6 U1793 ( .A(n2734), .B(n311), .C(n309), .D(n78), .Z(n2284) );
  HS65_LH_OAI22X6 U1794 ( .A(n2736), .B(n311), .C(n308), .D(n77), .Z(n2285) );
  HS65_LH_OAI22X6 U1795 ( .A(n2738), .B(n311), .C(n308), .D(n76), .Z(n2286) );
  HS65_LH_OAI22X6 U1796 ( .A(n2740), .B(n311), .C(n308), .D(n75), .Z(n2287) );
  HS65_LH_OAI22X6 U1797 ( .A(n2742), .B(n311), .C(n308), .D(n74), .Z(n2288) );
  HS65_LH_OAI22X6 U1798 ( .A(n2744), .B(n311), .C(n308), .D(n73), .Z(n2289) );
  HS65_LH_OAI22X6 U1799 ( .A(n2746), .B(n311), .C(n308), .D(n72), .Z(n2290) );
  HS65_LH_OAI22X6 U1800 ( .A(n2748), .B(n311), .C(n308), .D(n71), .Z(n2291) );
  HS65_LH_OAI22X6 U1801 ( .A(n2750), .B(n311), .C(n308), .D(n70), .Z(n2292) );
  HS65_LH_OAI22X6 U1802 ( .A(n2752), .B(n311), .C(n308), .D(n69), .Z(n2293) );
  HS65_LH_OAI22X6 U1803 ( .A(n2754), .B(n311), .C(n308), .D(n68), .Z(n2294) );
  HS65_LH_OAI22X6 U1804 ( .A(n2756), .B(n311), .C(n308), .D(n67), .Z(n2295) );
  HS65_LH_OAI22X6 U1805 ( .A(n2758), .B(n311), .C(n308), .D(n66), .Z(n2296) );
  HS65_LH_OAI22X6 U1806 ( .A(n2698), .B(n2475), .C(n2472), .D(n256), .Z(n1658)
         );
  HS65_LH_OAI22X6 U1807 ( .A(n2700), .B(n2475), .C(n2471), .D(n255), .Z(n1659)
         );
  HS65_LH_OAI22X6 U1808 ( .A(n2702), .B(n2475), .C(n2472), .D(n254), .Z(n1660)
         );
  HS65_LH_OAI22X6 U1809 ( .A(n2704), .B(n2475), .C(n2471), .D(n253), .Z(n1661)
         );
  HS65_LH_OAI22X6 U1810 ( .A(n2706), .B(n2475), .C(n2472), .D(n252), .Z(n1662)
         );
  HS65_LH_OAI22X6 U1811 ( .A(n2708), .B(n2475), .C(n2471), .D(n251), .Z(n1663)
         );
  HS65_LH_OAI22X6 U1812 ( .A(n2710), .B(n2475), .C(n2472), .D(n250), .Z(n1664)
         );
  HS65_LH_OAI22X6 U1813 ( .A(n2712), .B(n2475), .C(n2472), .D(n249), .Z(n1665)
         );
  HS65_LH_OAI22X6 U1814 ( .A(n2714), .B(n2475), .C(n2472), .D(n248), .Z(n1666)
         );
  HS65_LH_OAI22X6 U1815 ( .A(n2716), .B(n2475), .C(n2472), .D(n247), .Z(n1667)
         );
  HS65_LH_OAI22X6 U1816 ( .A(n2718), .B(n2475), .C(n2472), .D(n246), .Z(n1668)
         );
  HS65_LH_OAI22X6 U1817 ( .A(n2720), .B(n2475), .C(n2472), .D(n245), .Z(n1669)
         );
  HS65_LH_OAI22X6 U1818 ( .A(n2722), .B(n2475), .C(n2472), .D(n244), .Z(n1670)
         );
  HS65_LH_OAI22X6 U1819 ( .A(n2698), .B(n2470), .C(n2467), .D(n224), .Z(n1690)
         );
  HS65_LH_OAI22X6 U1820 ( .A(n2700), .B(n2470), .C(n2466), .D(n223), .Z(n1691)
         );
  HS65_LH_OAI22X6 U1821 ( .A(n2702), .B(n2470), .C(n2467), .D(n222), .Z(n1692)
         );
  HS65_LH_OAI22X6 U1822 ( .A(n2704), .B(n2470), .C(n2466), .D(n221), .Z(n1693)
         );
  HS65_LH_OAI22X6 U1823 ( .A(n2706), .B(n2470), .C(n2467), .D(n220), .Z(n1694)
         );
  HS65_LH_OAI22X6 U1824 ( .A(n2708), .B(n2470), .C(n2466), .D(n219), .Z(n1695)
         );
  HS65_LH_OAI22X6 U1825 ( .A(n2710), .B(n2470), .C(n2467), .D(n218), .Z(n1696)
         );
  HS65_LH_OAI22X6 U1826 ( .A(n2712), .B(n2470), .C(n2467), .D(n217), .Z(n1697)
         );
  HS65_LH_OAI22X6 U1827 ( .A(n2714), .B(n2470), .C(n2467), .D(n216), .Z(n1698)
         );
  HS65_LH_OAI22X6 U1828 ( .A(n2716), .B(n2470), .C(n2467), .D(n215), .Z(n1699)
         );
  HS65_LH_OAI22X6 U1829 ( .A(n2718), .B(n2470), .C(n2467), .D(n214), .Z(n1700)
         );
  HS65_LH_OAI22X6 U1830 ( .A(n2720), .B(n2470), .C(n2467), .D(n213), .Z(n1701)
         );
  HS65_LH_OAI22X6 U1831 ( .A(n2722), .B(n2470), .C(n2467), .D(n212), .Z(n1702)
         );
  HS65_LH_OAI22X6 U1832 ( .A(n2698), .B(n2445), .C(n2442), .D(n192), .Z(n1850)
         );
  HS65_LH_OAI22X6 U1833 ( .A(n2700), .B(n2445), .C(n2441), .D(n191), .Z(n1851)
         );
  HS65_LH_OAI22X6 U1834 ( .A(n2702), .B(n2445), .C(n2442), .D(n190), .Z(n1852)
         );
  HS65_LH_OAI22X6 U1835 ( .A(n2704), .B(n2445), .C(n2441), .D(n189), .Z(n1853)
         );
  HS65_LH_OAI22X6 U1836 ( .A(n2706), .B(n2445), .C(n2442), .D(n188), .Z(n1854)
         );
  HS65_LH_OAI22X6 U1837 ( .A(n2708), .B(n2445), .C(n2441), .D(n187), .Z(n1855)
         );
  HS65_LH_OAI22X6 U1838 ( .A(n2710), .B(n2445), .C(n2442), .D(n186), .Z(n1856)
         );
  HS65_LH_OAI22X6 U1839 ( .A(n2712), .B(n2445), .C(n2442), .D(n185), .Z(n1857)
         );
  HS65_LH_OAI22X6 U1840 ( .A(n2714), .B(n2445), .C(n2442), .D(n184), .Z(n1858)
         );
  HS65_LH_OAI22X6 U1841 ( .A(n2716), .B(n2445), .C(n2442), .D(n183), .Z(n1859)
         );
  HS65_LH_OAI22X6 U1842 ( .A(n2718), .B(n2445), .C(n2442), .D(n182), .Z(n1860)
         );
  HS65_LH_OAI22X6 U1843 ( .A(n2720), .B(n2445), .C(n2442), .D(n181), .Z(n1861)
         );
  HS65_LH_OAI22X6 U1844 ( .A(n2722), .B(n2445), .C(n2442), .D(n180), .Z(n1862)
         );
  HS65_LH_OAI22X6 U1845 ( .A(n2698), .B(n2440), .C(n2437), .D(n160), .Z(n1882)
         );
  HS65_LH_OAI22X6 U1846 ( .A(n2700), .B(n2440), .C(n2436), .D(n159), .Z(n1883)
         );
  HS65_LH_OAI22X6 U1847 ( .A(n2702), .B(n2440), .C(n2437), .D(n158), .Z(n1884)
         );
  HS65_LH_OAI22X6 U1848 ( .A(n2704), .B(n2440), .C(n2436), .D(n157), .Z(n1885)
         );
  HS65_LH_OAI22X6 U1849 ( .A(n2706), .B(n2440), .C(n2437), .D(n156), .Z(n1886)
         );
  HS65_LH_OAI22X6 U1850 ( .A(n2708), .B(n2440), .C(n2436), .D(n155), .Z(n1887)
         );
  HS65_LH_OAI22X6 U1851 ( .A(n2710), .B(n2440), .C(n2437), .D(n154), .Z(n1888)
         );
  HS65_LH_OAI22X6 U1852 ( .A(n2712), .B(n2440), .C(n2437), .D(n153), .Z(n1889)
         );
  HS65_LH_OAI22X6 U1853 ( .A(n2714), .B(n2440), .C(n2437), .D(n152), .Z(n1890)
         );
  HS65_LH_OAI22X6 U1854 ( .A(n2716), .B(n2440), .C(n2437), .D(n151), .Z(n1891)
         );
  HS65_LH_OAI22X6 U1855 ( .A(n2718), .B(n2440), .C(n2437), .D(n150), .Z(n1892)
         );
  HS65_LH_OAI22X6 U1856 ( .A(n2720), .B(n2440), .C(n2437), .D(n149), .Z(n1893)
         );
  HS65_LH_OAI22X6 U1857 ( .A(n2722), .B(n2440), .C(n2437), .D(n148), .Z(n1894)
         );
  HS65_LH_OAI22X6 U1858 ( .A(n2698), .B(n307), .C(n304), .D(n64), .Z(n2298) );
  HS65_LH_OAI22X6 U1859 ( .A(n2700), .B(n307), .C(n303), .D(n63), .Z(n2299) );
  HS65_LH_OAI22X6 U1860 ( .A(n2702), .B(n307), .C(n304), .D(n62), .Z(n2300) );
  HS65_LH_OAI22X6 U1861 ( .A(n2704), .B(n307), .C(n303), .D(n61), .Z(n2301) );
  HS65_LH_OAI22X6 U1862 ( .A(n2706), .B(n307), .C(n304), .D(n60), .Z(n2302) );
  HS65_LH_OAI22X6 U1863 ( .A(n2708), .B(n307), .C(n303), .D(n59), .Z(n2303) );
  HS65_LH_OAI22X6 U1864 ( .A(n2710), .B(n307), .C(n304), .D(n58), .Z(n2304) );
  HS65_LH_OAI22X6 U1865 ( .A(n2712), .B(n307), .C(n304), .D(n57), .Z(n2305) );
  HS65_LH_OAI22X6 U1866 ( .A(n2714), .B(n307), .C(n304), .D(n56), .Z(n2306) );
  HS65_LH_OAI22X6 U1867 ( .A(n2716), .B(n307), .C(n304), .D(n55), .Z(n2307) );
  HS65_LH_OAI22X6 U1868 ( .A(n2718), .B(n307), .C(n304), .D(n54), .Z(n2308) );
  HS65_LH_OAI22X6 U1869 ( .A(n2720), .B(n307), .C(n304), .D(n53), .Z(n2309) );
  HS65_LH_OAI22X6 U1870 ( .A(n2722), .B(n307), .C(n304), .D(n52), .Z(n2310) );
  HS65_LH_OAI22X6 U1871 ( .A(n2698), .B(n302), .C(n299), .D(n32), .Z(n2330) );
  HS65_LH_OAI22X6 U1872 ( .A(n2700), .B(n302), .C(n298), .D(n31), .Z(n2331) );
  HS65_LH_OAI22X6 U1873 ( .A(n2702), .B(n302), .C(n299), .D(n30), .Z(n2332) );
  HS65_LH_OAI22X6 U1874 ( .A(n2704), .B(n302), .C(n298), .D(n29), .Z(n2333) );
  HS65_LH_OAI22X6 U1875 ( .A(n2706), .B(n302), .C(n299), .D(n28), .Z(n2334) );
  HS65_LH_OAI22X6 U1876 ( .A(n2708), .B(n302), .C(n298), .D(n27), .Z(n2335) );
  HS65_LH_OAI22X6 U1877 ( .A(n2710), .B(n302), .C(n299), .D(n26), .Z(n2336) );
  HS65_LH_OAI22X6 U1878 ( .A(n2712), .B(n302), .C(n299), .D(n25), .Z(n2337) );
  HS65_LH_OAI22X6 U1879 ( .A(n2714), .B(n302), .C(n299), .D(n24), .Z(n2338) );
  HS65_LH_OAI22X6 U1880 ( .A(n2716), .B(n302), .C(n299), .D(n23), .Z(n2339) );
  HS65_LH_OAI22X6 U1881 ( .A(n2718), .B(n302), .C(n299), .D(n22), .Z(n2340) );
  HS65_LH_OAI22X6 U1882 ( .A(n2720), .B(n302), .C(n299), .D(n21), .Z(n2341) );
  HS65_LH_OAI22X6 U1883 ( .A(n2722), .B(n302), .C(n299), .D(n20), .Z(n2342) );
  HS65_LH_OAI22X6 U1884 ( .A(n2698), .B(n317), .C(n314), .D(n128), .Z(n2234)
         );
  HS65_LH_OAI22X6 U1885 ( .A(n2700), .B(n317), .C(n313), .D(n127), .Z(n2235)
         );
  HS65_LH_OAI22X6 U1886 ( .A(n2702), .B(n317), .C(n314), .D(n126), .Z(n2236)
         );
  HS65_LH_OAI22X6 U1887 ( .A(n2704), .B(n317), .C(n313), .D(n125), .Z(n2237)
         );
  HS65_LH_OAI22X6 U1888 ( .A(n2706), .B(n317), .C(n314), .D(n124), .Z(n2238)
         );
  HS65_LH_OAI22X6 U1889 ( .A(n2708), .B(n317), .C(n313), .D(n123), .Z(n2239)
         );
  HS65_LH_OAI22X6 U1890 ( .A(n2710), .B(n317), .C(n314), .D(n122), .Z(n2240)
         );
  HS65_LH_OAI22X6 U1891 ( .A(n2712), .B(n317), .C(n314), .D(n121), .Z(n2241)
         );
  HS65_LH_OAI22X6 U1892 ( .A(n2714), .B(n317), .C(n314), .D(n120), .Z(n2242)
         );
  HS65_LH_OAI22X6 U1893 ( .A(n2716), .B(n317), .C(n314), .D(n119), .Z(n2243)
         );
  HS65_LH_OAI22X6 U1894 ( .A(n2718), .B(n317), .C(n314), .D(n118), .Z(n2244)
         );
  HS65_LH_OAI22X6 U1895 ( .A(n2720), .B(n317), .C(n314), .D(n117), .Z(n2245)
         );
  HS65_LH_OAI22X6 U1896 ( .A(n2722), .B(n317), .C(n314), .D(n116), .Z(n2246)
         );
  HS65_LH_OAI22X6 U1897 ( .A(n2698), .B(n312), .C(n309), .D(n96), .Z(n2266) );
  HS65_LH_OAI22X6 U1898 ( .A(n2700), .B(n312), .C(n308), .D(n95), .Z(n2267) );
  HS65_LH_OAI22X6 U1899 ( .A(n2702), .B(n312), .C(n309), .D(n94), .Z(n2268) );
  HS65_LH_OAI22X6 U1900 ( .A(n2704), .B(n312), .C(n308), .D(n93), .Z(n2269) );
  HS65_LH_OAI22X6 U1901 ( .A(n2706), .B(n312), .C(n309), .D(n92), .Z(n2270) );
  HS65_LH_OAI22X6 U1902 ( .A(n2708), .B(n312), .C(n308), .D(n91), .Z(n2271) );
  HS65_LH_OAI22X6 U1903 ( .A(n2710), .B(n312), .C(n309), .D(n90), .Z(n2272) );
  HS65_LH_OAI22X6 U1904 ( .A(n2712), .B(n312), .C(n309), .D(n89), .Z(n2273) );
  HS65_LH_OAI22X6 U1905 ( .A(n2714), .B(n312), .C(n309), .D(n88), .Z(n2274) );
  HS65_LH_OAI22X6 U1906 ( .A(n2716), .B(n312), .C(n309), .D(n87), .Z(n2275) );
  HS65_LH_OAI22X6 U1907 ( .A(n2718), .B(n312), .C(n309), .D(n86), .Z(n2276) );
  HS65_LH_OAI22X6 U1908 ( .A(n2720), .B(n312), .C(n309), .D(n85), .Z(n2277) );
  HS65_LH_OAI22X6 U1909 ( .A(n2722), .B(n312), .C(n309), .D(n84), .Z(n2278) );
  HS65_LH_NAND3X5 U1910 ( .A(n2908), .B(n2909), .C(n2910), .Z(n836) );
  HS65_LH_NAND2X7 U1911 ( .A(\registers[1][0] ), .B(n2670), .Z(n2910) );
  HS65_LH_NAND2X7 U1912 ( .A(\registers[3][0] ), .B(n2664), .Z(n2909) );
  HS65_LH_NAND2X7 U1913 ( .A(\registers[2][0] ), .B(n2667), .Z(n2908) );
  HS65_LH_NAND3X5 U1914 ( .A(n2914), .B(n2915), .C(n2916), .Z(n671) );
  HS65_LH_NAND2X7 U1915 ( .A(\registers[1][1] ), .B(n2670), .Z(n2916) );
  HS65_LH_NAND2X7 U1916 ( .A(\registers[3][1] ), .B(n2664), .Z(n2915) );
  HS65_LH_NAND2X7 U1917 ( .A(\registers[2][1] ), .B(n2667), .Z(n2914) );
  HS65_LH_NAND3X5 U1918 ( .A(n2920), .B(n2921), .C(n2922), .Z(n506) );
  HS65_LH_NAND2X7 U1919 ( .A(\registers[1][2] ), .B(n2670), .Z(n2922) );
  HS65_LH_NAND2X7 U1920 ( .A(\registers[3][2] ), .B(n2664), .Z(n2921) );
  HS65_LH_NAND2X7 U1921 ( .A(\registers[2][2] ), .B(n2667), .Z(n2920) );
  HS65_LH_NAND3X5 U1922 ( .A(n2926), .B(n2927), .C(n2928), .Z(n461) );
  HS65_LH_NAND2X7 U1923 ( .A(\registers[1][3] ), .B(n2670), .Z(n2928) );
  HS65_LH_NAND2X7 U1924 ( .A(\registers[3][3] ), .B(n2664), .Z(n2927) );
  HS65_LH_NAND2X7 U1925 ( .A(\registers[2][3] ), .B(n2667), .Z(n2926) );
  HS65_LH_NAND3X5 U1926 ( .A(n2932), .B(n2933), .C(n2934), .Z(n446) );
  HS65_LH_NAND2X7 U1927 ( .A(\registers[1][4] ), .B(n2670), .Z(n2934) );
  HS65_LH_NAND2X7 U1928 ( .A(\registers[3][4] ), .B(n2664), .Z(n2933) );
  HS65_LH_NAND2X7 U1929 ( .A(\registers[2][4] ), .B(n2667), .Z(n2932) );
  HS65_LH_NAND3X5 U1930 ( .A(n2938), .B(n2939), .C(n2940), .Z(n431) );
  HS65_LH_NAND2X7 U1931 ( .A(\registers[1][5] ), .B(n2670), .Z(n2940) );
  HS65_LH_NAND2X7 U1932 ( .A(\registers[3][5] ), .B(n2664), .Z(n2939) );
  HS65_LH_NAND2X7 U1933 ( .A(\registers[2][5] ), .B(n2667), .Z(n2938) );
  HS65_LH_NAND3X5 U1934 ( .A(n2944), .B(n2945), .C(n2946), .Z(n416) );
  HS65_LH_NAND2X7 U1935 ( .A(\registers[1][6] ), .B(n2670), .Z(n2946) );
  HS65_LH_NAND2X7 U1936 ( .A(\registers[3][6] ), .B(n2664), .Z(n2945) );
  HS65_LH_NAND2X7 U1937 ( .A(\registers[2][6] ), .B(n2667), .Z(n2944) );
  HS65_LH_NAND3X5 U1938 ( .A(n2950), .B(n2951), .C(n2952), .Z(n401) );
  HS65_LH_NAND2X7 U1939 ( .A(\registers[1][7] ), .B(n2670), .Z(n2952) );
  HS65_LH_NAND2X7 U1940 ( .A(\registers[3][7] ), .B(n2664), .Z(n2951) );
  HS65_LH_NAND2X7 U1941 ( .A(\registers[2][7] ), .B(n2667), .Z(n2950) );
  HS65_LH_NAND3X5 U1942 ( .A(n2956), .B(n2957), .C(n2958), .Z(n386) );
  HS65_LH_NAND2X7 U1943 ( .A(\registers[1][8] ), .B(n2670), .Z(n2958) );
  HS65_LH_NAND2X7 U1944 ( .A(\registers[3][8] ), .B(n2664), .Z(n2957) );
  HS65_LH_NAND2X7 U1945 ( .A(\registers[2][8] ), .B(n2667), .Z(n2956) );
  HS65_LH_NAND3X5 U1946 ( .A(n2962), .B(n2963), .C(n2964), .Z(n339) );
  HS65_LH_NAND2X7 U1947 ( .A(\registers[1][9] ), .B(n2670), .Z(n2964) );
  HS65_LH_NAND2X7 U1948 ( .A(\registers[3][9] ), .B(n2664), .Z(n2963) );
  HS65_LH_NAND2X7 U1949 ( .A(\registers[2][9] ), .B(n2667), .Z(n2962) );
  HS65_LH_NAND3X5 U1950 ( .A(n2974), .B(n2975), .C(n2976), .Z(n806) );
  HS65_LH_NAND2X7 U1951 ( .A(\registers[1][11] ), .B(n2670), .Z(n2976) );
  HS65_LH_NAND2X7 U1952 ( .A(\registers[3][11] ), .B(n2664), .Z(n2975) );
  HS65_LH_NAND2X7 U1953 ( .A(\registers[2][11] ), .B(n2667), .Z(n2974) );
  HS65_LH_NAND3X5 U1954 ( .A(n2980), .B(n2981), .C(n2982), .Z(n791) );
  HS65_LH_NAND2X7 U1955 ( .A(\registers[1][12] ), .B(n2671), .Z(n2982) );
  HS65_LH_NAND2X7 U1956 ( .A(\registers[3][12] ), .B(n2665), .Z(n2981) );
  HS65_LH_NAND2X7 U1957 ( .A(\registers[2][12] ), .B(n2668), .Z(n2980) );
  HS65_LH_NAND3X5 U1958 ( .A(n2986), .B(n2987), .C(n2988), .Z(n776) );
  HS65_LH_NAND2X7 U1959 ( .A(\registers[1][13] ), .B(n2671), .Z(n2988) );
  HS65_LH_NAND2X7 U1960 ( .A(\registers[3][13] ), .B(n2665), .Z(n2987) );
  HS65_LH_NAND2X7 U1961 ( .A(\registers[2][13] ), .B(n2668), .Z(n2986) );
  HS65_LH_NAND3X5 U1962 ( .A(n2992), .B(n2993), .C(n2994), .Z(n761) );
  HS65_LH_NAND2X7 U1963 ( .A(\registers[1][14] ), .B(n2671), .Z(n2994) );
  HS65_LH_NAND2X7 U1964 ( .A(\registers[3][14] ), .B(n2665), .Z(n2993) );
  HS65_LH_NAND2X7 U1965 ( .A(\registers[2][14] ), .B(n2668), .Z(n2992) );
  HS65_LH_NAND3X5 U1966 ( .A(n2998), .B(n2999), .C(n3000), .Z(n746) );
  HS65_LH_NAND2X7 U1967 ( .A(\registers[1][15] ), .B(n2671), .Z(n3000) );
  HS65_LH_NAND2X7 U1968 ( .A(\registers[3][15] ), .B(n2665), .Z(n2999) );
  HS65_LH_NAND2X7 U1969 ( .A(\registers[2][15] ), .B(n2668), .Z(n2998) );
  HS65_LH_NAND3X5 U1970 ( .A(n3004), .B(n3005), .C(n3006), .Z(n731) );
  HS65_LH_NAND2X7 U1971 ( .A(\registers[1][16] ), .B(n2671), .Z(n3006) );
  HS65_LH_NAND2X7 U1972 ( .A(\registers[3][16] ), .B(n2665), .Z(n3005) );
  HS65_LH_NAND2X7 U1973 ( .A(\registers[2][16] ), .B(n2668), .Z(n3004) );
  HS65_LH_NAND3X5 U1974 ( .A(n3010), .B(n3011), .C(n3012), .Z(n716) );
  HS65_LH_NAND2X7 U1975 ( .A(\registers[1][17] ), .B(n2671), .Z(n3012) );
  HS65_LH_NAND2X7 U1976 ( .A(\registers[3][17] ), .B(n2665), .Z(n3011) );
  HS65_LH_NAND2X7 U1977 ( .A(\registers[2][17] ), .B(n2668), .Z(n3010) );
  HS65_LH_NAND3X5 U1978 ( .A(n3016), .B(n3017), .C(n3018), .Z(n701) );
  HS65_LH_NAND2X7 U1979 ( .A(\registers[1][18] ), .B(n2671), .Z(n3018) );
  HS65_LH_NAND2X7 U1980 ( .A(\registers[3][18] ), .B(n2665), .Z(n3017) );
  HS65_LH_NAND2X7 U1981 ( .A(\registers[2][18] ), .B(n2668), .Z(n3016) );
  HS65_LH_NAND3X5 U1982 ( .A(n3022), .B(n3023), .C(n3024), .Z(n686) );
  HS65_LH_NAND2X7 U1983 ( .A(\registers[1][19] ), .B(n2671), .Z(n3024) );
  HS65_LH_NAND2X7 U1984 ( .A(\registers[3][19] ), .B(n2665), .Z(n3023) );
  HS65_LH_NAND2X7 U1985 ( .A(\registers[2][19] ), .B(n2668), .Z(n3022) );
  HS65_LH_NAND3X5 U1986 ( .A(n3028), .B(n3029), .C(n3030), .Z(n656) );
  HS65_LH_NAND2X7 U1987 ( .A(\registers[1][20] ), .B(n2671), .Z(n3030) );
  HS65_LH_NAND2X7 U1988 ( .A(\registers[3][20] ), .B(n2665), .Z(n3029) );
  HS65_LH_NAND2X7 U1989 ( .A(\registers[2][20] ), .B(n2668), .Z(n3028) );
  HS65_LH_NAND3X5 U1990 ( .A(n3034), .B(n3035), .C(n3036), .Z(n641) );
  HS65_LH_NAND2X7 U1991 ( .A(\registers[1][21] ), .B(n2671), .Z(n3036) );
  HS65_LH_NAND2X7 U1992 ( .A(\registers[3][21] ), .B(n2665), .Z(n3035) );
  HS65_LH_NAND2X7 U1993 ( .A(\registers[2][21] ), .B(n2668), .Z(n3034) );
  HS65_LH_NAND3X5 U1994 ( .A(n3040), .B(n3041), .C(n3042), .Z(n626) );
  HS65_LH_NAND2X7 U1995 ( .A(\registers[1][22] ), .B(n2671), .Z(n3042) );
  HS65_LH_NAND2X7 U1996 ( .A(\registers[3][22] ), .B(n2665), .Z(n3041) );
  HS65_LH_NAND2X7 U1997 ( .A(\registers[2][22] ), .B(n2668), .Z(n3040) );
  HS65_LH_NAND3X5 U1998 ( .A(n3046), .B(n3047), .C(n3048), .Z(n611) );
  HS65_LH_NAND2X7 U1999 ( .A(\registers[1][23] ), .B(n2671), .Z(n3048) );
  HS65_LH_NAND2X7 U2000 ( .A(\registers[3][23] ), .B(n2665), .Z(n3047) );
  HS65_LH_NAND2X7 U2001 ( .A(\registers[2][23] ), .B(n2668), .Z(n3046) );
  HS65_LH_NAND3X5 U2002 ( .A(n3052), .B(n3053), .C(n3054), .Z(n596) );
  HS65_LH_NAND2X7 U2003 ( .A(\registers[1][24] ), .B(n2672), .Z(n3054) );
  HS65_LH_NAND2X7 U2004 ( .A(\registers[3][24] ), .B(n2666), .Z(n3053) );
  HS65_LH_NAND2X7 U2005 ( .A(\registers[2][24] ), .B(n2669), .Z(n3052) );
  HS65_LH_NAND3X5 U2006 ( .A(n3058), .B(n3059), .C(n3060), .Z(n581) );
  HS65_LH_NAND2X7 U2007 ( .A(\registers[1][25] ), .B(n2672), .Z(n3060) );
  HS65_LH_NAND2X7 U2008 ( .A(\registers[3][25] ), .B(n2666), .Z(n3059) );
  HS65_LH_NAND2X7 U2009 ( .A(\registers[2][25] ), .B(n2669), .Z(n3058) );
  HS65_LH_NAND3X5 U2010 ( .A(n3064), .B(n3065), .C(n3066), .Z(n566) );
  HS65_LH_NAND2X7 U2011 ( .A(\registers[1][26] ), .B(n2672), .Z(n3066) );
  HS65_LH_NAND2X7 U2012 ( .A(\registers[3][26] ), .B(n2666), .Z(n3065) );
  HS65_LH_NAND2X7 U2013 ( .A(\registers[2][26] ), .B(n2669), .Z(n3064) );
  HS65_LH_NAND3X5 U2014 ( .A(n3070), .B(n3071), .C(n3072), .Z(n551) );
  HS65_LH_NAND2X7 U2015 ( .A(\registers[1][27] ), .B(n2672), .Z(n3072) );
  HS65_LH_NAND2X7 U2016 ( .A(\registers[3][27] ), .B(n2666), .Z(n3071) );
  HS65_LH_NAND2X7 U2017 ( .A(\registers[2][27] ), .B(n2669), .Z(n3070) );
  HS65_LH_NAND3X5 U2018 ( .A(n3076), .B(n3077), .C(n3078), .Z(n536) );
  HS65_LH_NAND2X7 U2019 ( .A(\registers[1][28] ), .B(n2672), .Z(n3078) );
  HS65_LH_NAND2X7 U2020 ( .A(\registers[3][28] ), .B(n2666), .Z(n3077) );
  HS65_LH_NAND2X7 U2021 ( .A(\registers[2][28] ), .B(n2669), .Z(n3076) );
  HS65_LH_NAND3X5 U2022 ( .A(n3082), .B(n3083), .C(n3084), .Z(n521) );
  HS65_LH_NAND2X7 U2023 ( .A(\registers[1][29] ), .B(n2672), .Z(n3084) );
  HS65_LH_NAND2X7 U2024 ( .A(\registers[3][29] ), .B(n2666), .Z(n3083) );
  HS65_LH_NAND2X7 U2025 ( .A(\registers[2][29] ), .B(n2669), .Z(n3082) );
  HS65_LH_NAND3X5 U2026 ( .A(n3088), .B(n3089), .C(n3090), .Z(n491) );
  HS65_LH_NAND2X7 U2027 ( .A(\registers[1][30] ), .B(n2672), .Z(n3090) );
  HS65_LH_NAND2X7 U2028 ( .A(\registers[3][30] ), .B(n2666), .Z(n3089) );
  HS65_LH_NAND2X7 U2029 ( .A(\registers[2][30] ), .B(n2669), .Z(n3088) );
  HS65_LH_NAND3X5 U2030 ( .A(n3094), .B(n3095), .C(n3096), .Z(n476) );
  HS65_LH_NAND2X7 U2031 ( .A(\registers[1][31] ), .B(n2672), .Z(n3096) );
  HS65_LH_NAND2X7 U2032 ( .A(\registers[3][31] ), .B(n2666), .Z(n3095) );
  HS65_LH_NAND2X7 U2033 ( .A(\registers[2][31] ), .B(n2669), .Z(n3094) );
  HS65_LH_NAND3X5 U2034 ( .A(n2911), .B(n2912), .C(n2913), .Z(n1364) );
  HS65_LH_NAND2X7 U2035 ( .A(n2577), .B(\registers[1][0] ), .Z(n2913) );
  HS65_LH_NAND2X7 U2036 ( .A(n2571), .B(\registers[3][0] ), .Z(n2912) );
  HS65_LH_NAND2X7 U2037 ( .A(n2574), .B(\registers[2][0] ), .Z(n2911) );
  HS65_LH_NAND3X5 U2038 ( .A(n2917), .B(n2918), .C(n2919), .Z(n1199) );
  HS65_LH_NAND2X7 U2039 ( .A(n2577), .B(\registers[1][1] ), .Z(n2919) );
  HS65_LH_NAND2X7 U2040 ( .A(n2571), .B(\registers[3][1] ), .Z(n2918) );
  HS65_LH_NAND2X7 U2041 ( .A(n2574), .B(\registers[2][1] ), .Z(n2917) );
  HS65_LH_NAND3X5 U2042 ( .A(n2923), .B(n2924), .C(n2925), .Z(n1034) );
  HS65_LH_NAND2X7 U2043 ( .A(n2577), .B(\registers[1][2] ), .Z(n2925) );
  HS65_LH_NAND2X7 U2044 ( .A(n2571), .B(\registers[3][2] ), .Z(n2924) );
  HS65_LH_NAND2X7 U2045 ( .A(n2574), .B(\registers[2][2] ), .Z(n2923) );
  HS65_LH_NAND3X5 U2046 ( .A(n2929), .B(n2930), .C(n2931), .Z(n989) );
  HS65_LH_NAND2X7 U2047 ( .A(n2577), .B(\registers[1][3] ), .Z(n2931) );
  HS65_LH_NAND2X7 U2048 ( .A(n2571), .B(\registers[3][3] ), .Z(n2930) );
  HS65_LH_NAND2X7 U2049 ( .A(n2574), .B(\registers[2][3] ), .Z(n2929) );
  HS65_LH_NAND3X5 U2050 ( .A(n2935), .B(n2936), .C(n2937), .Z(n974) );
  HS65_LH_NAND2X7 U2051 ( .A(n2577), .B(\registers[1][4] ), .Z(n2937) );
  HS65_LH_NAND2X7 U2052 ( .A(n2571), .B(\registers[3][4] ), .Z(n2936) );
  HS65_LH_NAND2X7 U2053 ( .A(n2574), .B(\registers[2][4] ), .Z(n2935) );
  HS65_LH_NAND3X5 U2054 ( .A(n2941), .B(n2942), .C(n2943), .Z(n959) );
  HS65_LH_NAND2X7 U2055 ( .A(n2577), .B(\registers[1][5] ), .Z(n2943) );
  HS65_LH_NAND2X7 U2056 ( .A(n2571), .B(\registers[3][5] ), .Z(n2942) );
  HS65_LH_NAND2X7 U2057 ( .A(n2574), .B(\registers[2][5] ), .Z(n2941) );
  HS65_LH_NAND3X5 U2058 ( .A(n2947), .B(n2948), .C(n2949), .Z(n944) );
  HS65_LH_NAND2X7 U2059 ( .A(n2577), .B(\registers[1][6] ), .Z(n2949) );
  HS65_LH_NAND2X7 U2060 ( .A(n2571), .B(\registers[3][6] ), .Z(n2948) );
  HS65_LH_NAND2X7 U2061 ( .A(n2574), .B(\registers[2][6] ), .Z(n2947) );
  HS65_LH_NAND3X5 U2062 ( .A(n2953), .B(n2954), .C(n2955), .Z(n929) );
  HS65_LH_NAND2X7 U2063 ( .A(n2577), .B(\registers[1][7] ), .Z(n2955) );
  HS65_LH_NAND2X7 U2064 ( .A(n2571), .B(\registers[3][7] ), .Z(n2954) );
  HS65_LH_NAND2X7 U2065 ( .A(n2574), .B(\registers[2][7] ), .Z(n2953) );
  HS65_LH_NAND3X5 U2066 ( .A(n2959), .B(n2960), .C(n2961), .Z(n914) );
  HS65_LH_NAND2X7 U2067 ( .A(n2577), .B(\registers[1][8] ), .Z(n2961) );
  HS65_LH_NAND2X7 U2068 ( .A(n2571), .B(\registers[3][8] ), .Z(n2960) );
  HS65_LH_NAND2X7 U2069 ( .A(n2574), .B(\registers[2][8] ), .Z(n2959) );
  HS65_LH_NAND3X5 U2070 ( .A(n2965), .B(n2966), .C(n2967), .Z(n867) );
  HS65_LH_NAND2X7 U2071 ( .A(n2577), .B(\registers[1][9] ), .Z(n2967) );
  HS65_LH_NAND2X7 U2072 ( .A(n2571), .B(\registers[3][9] ), .Z(n2966) );
  HS65_LH_NAND2X7 U2073 ( .A(n2574), .B(\registers[2][9] ), .Z(n2965) );
  HS65_LH_NAND3X5 U2074 ( .A(n2971), .B(n2972), .C(n2973), .Z(n1349) );
  HS65_LH_NAND2X7 U2075 ( .A(n2577), .B(\registers[1][10] ), .Z(n2973) );
  HS65_LH_NAND2X7 U2076 ( .A(n2571), .B(\registers[3][10] ), .Z(n2972) );
  HS65_LH_NAND2X7 U2077 ( .A(n2574), .B(\registers[2][10] ), .Z(n2971) );
  HS65_LH_NAND3X5 U2078 ( .A(n2977), .B(n2978), .C(n2979), .Z(n1334) );
  HS65_LH_NAND2X7 U2079 ( .A(n2577), .B(\registers[1][11] ), .Z(n2979) );
  HS65_LH_NAND2X7 U2080 ( .A(n2571), .B(\registers[3][11] ), .Z(n2978) );
  HS65_LH_NAND2X7 U2081 ( .A(n2574), .B(\registers[2][11] ), .Z(n2977) );
  HS65_LH_NAND3X5 U2082 ( .A(n2983), .B(n2984), .C(n2985), .Z(n1319) );
  HS65_LH_NAND2X7 U2083 ( .A(n2577), .B(\registers[1][12] ), .Z(n2985) );
  HS65_LH_NAND2X7 U2084 ( .A(n2571), .B(\registers[3][12] ), .Z(n2984) );
  HS65_LH_NAND2X7 U2085 ( .A(n2574), .B(\registers[2][12] ), .Z(n2983) );
  HS65_LH_NAND3X5 U2086 ( .A(n2989), .B(n2990), .C(n2991), .Z(n1304) );
  HS65_LH_NAND2X7 U2087 ( .A(n2578), .B(\registers[1][13] ), .Z(n2991) );
  HS65_LH_NAND2X7 U2088 ( .A(n2572), .B(\registers[3][13] ), .Z(n2990) );
  HS65_LH_NAND2X7 U2089 ( .A(n2575), .B(\registers[2][13] ), .Z(n2989) );
  HS65_LH_NAND3X5 U2090 ( .A(n2995), .B(n2996), .C(n2997), .Z(n1289) );
  HS65_LH_NAND2X7 U2091 ( .A(n2578), .B(\registers[1][14] ), .Z(n2997) );
  HS65_LH_NAND2X7 U2092 ( .A(n2572), .B(\registers[3][14] ), .Z(n2996) );
  HS65_LH_NAND2X7 U2093 ( .A(n2575), .B(\registers[2][14] ), .Z(n2995) );
  HS65_LH_NAND3X5 U2094 ( .A(n3001), .B(n3002), .C(n3003), .Z(n1274) );
  HS65_LH_NAND2X7 U2095 ( .A(n2578), .B(\registers[1][15] ), .Z(n3003) );
  HS65_LH_NAND2X7 U2096 ( .A(n2572), .B(\registers[3][15] ), .Z(n3002) );
  HS65_LH_NAND2X7 U2097 ( .A(n2575), .B(\registers[2][15] ), .Z(n3001) );
  HS65_LH_NAND3X5 U2098 ( .A(n3007), .B(n3008), .C(n3009), .Z(n1259) );
  HS65_LH_NAND2X7 U2099 ( .A(n2578), .B(\registers[1][16] ), .Z(n3009) );
  HS65_LH_NAND2X7 U2100 ( .A(n2572), .B(\registers[3][16] ), .Z(n3008) );
  HS65_LH_NAND2X7 U2101 ( .A(n2575), .B(\registers[2][16] ), .Z(n3007) );
  HS65_LH_NAND3X5 U2102 ( .A(n3013), .B(n3014), .C(n3015), .Z(n1244) );
  HS65_LH_NAND2X7 U2103 ( .A(n2578), .B(\registers[1][17] ), .Z(n3015) );
  HS65_LH_NAND2X7 U2104 ( .A(n2572), .B(\registers[3][17] ), .Z(n3014) );
  HS65_LH_NAND2X7 U2105 ( .A(n2575), .B(\registers[2][17] ), .Z(n3013) );
  HS65_LH_NAND3X5 U2106 ( .A(n3019), .B(n3020), .C(n3021), .Z(n1229) );
  HS65_LH_NAND2X7 U2107 ( .A(n2578), .B(\registers[1][18] ), .Z(n3021) );
  HS65_LH_NAND2X7 U2108 ( .A(n2572), .B(\registers[3][18] ), .Z(n3020) );
  HS65_LH_NAND2X7 U2109 ( .A(n2575), .B(\registers[2][18] ), .Z(n3019) );
  HS65_LH_NAND3X5 U2110 ( .A(n3025), .B(n3026), .C(n3027), .Z(n1214) );
  HS65_LH_NAND2X7 U2111 ( .A(n2578), .B(\registers[1][19] ), .Z(n3027) );
  HS65_LH_NAND2X7 U2112 ( .A(n2572), .B(\registers[3][19] ), .Z(n3026) );
  HS65_LH_NAND2X7 U2113 ( .A(n2575), .B(\registers[2][19] ), .Z(n3025) );
  HS65_LH_NAND3X5 U2114 ( .A(n3031), .B(n3032), .C(n3033), .Z(n1184) );
  HS65_LH_NAND2X7 U2115 ( .A(n2578), .B(\registers[1][20] ), .Z(n3033) );
  HS65_LH_NAND2X7 U2116 ( .A(n2572), .B(\registers[3][20] ), .Z(n3032) );
  HS65_LH_NAND2X7 U2117 ( .A(n2575), .B(\registers[2][20] ), .Z(n3031) );
  HS65_LH_NAND3X5 U2118 ( .A(n3037), .B(n3038), .C(n3039), .Z(n1169) );
  HS65_LH_NAND2X7 U2119 ( .A(n2578), .B(\registers[1][21] ), .Z(n3039) );
  HS65_LH_NAND2X7 U2120 ( .A(n2572), .B(\registers[3][21] ), .Z(n3038) );
  HS65_LH_NAND2X7 U2121 ( .A(n2575), .B(\registers[2][21] ), .Z(n3037) );
  HS65_LH_NAND3X5 U2122 ( .A(n3043), .B(n3044), .C(n3045), .Z(n1154) );
  HS65_LH_NAND2X7 U2123 ( .A(n2578), .B(\registers[1][22] ), .Z(n3045) );
  HS65_LH_NAND2X7 U2124 ( .A(n2572), .B(\registers[3][22] ), .Z(n3044) );
  HS65_LH_NAND2X7 U2125 ( .A(n2575), .B(\registers[2][22] ), .Z(n3043) );
  HS65_LH_NAND3X5 U2126 ( .A(n3049), .B(n3050), .C(n3051), .Z(n1139) );
  HS65_LH_NAND2X7 U2127 ( .A(n2578), .B(\registers[1][23] ), .Z(n3051) );
  HS65_LH_NAND2X7 U2128 ( .A(n2572), .B(\registers[3][23] ), .Z(n3050) );
  HS65_LH_NAND2X7 U2129 ( .A(n2575), .B(\registers[2][23] ), .Z(n3049) );
  HS65_LH_NAND3X5 U2130 ( .A(n3055), .B(n3056), .C(n3057), .Z(n1124) );
  HS65_LH_NAND2X7 U2131 ( .A(n2578), .B(\registers[1][24] ), .Z(n3057) );
  HS65_LH_NAND2X7 U2132 ( .A(n2572), .B(\registers[3][24] ), .Z(n3056) );
  HS65_LH_NAND2X7 U2133 ( .A(n2575), .B(\registers[2][24] ), .Z(n3055) );
  HS65_LH_NAND3X5 U2134 ( .A(n3061), .B(n3062), .C(n3063), .Z(n1109) );
  HS65_LH_NAND2X7 U2135 ( .A(n2578), .B(\registers[1][25] ), .Z(n3063) );
  HS65_LH_NAND2X7 U2136 ( .A(n2572), .B(\registers[3][25] ), .Z(n3062) );
  HS65_LH_NAND2X7 U2137 ( .A(n2575), .B(\registers[2][25] ), .Z(n3061) );
  HS65_LH_NAND3X5 U2138 ( .A(n3067), .B(n3068), .C(n3069), .Z(n1094) );
  HS65_LH_NAND2X7 U2139 ( .A(n2579), .B(\registers[1][26] ), .Z(n3069) );
  HS65_LH_NAND2X7 U2140 ( .A(n2573), .B(\registers[3][26] ), .Z(n3068) );
  HS65_LH_NAND2X7 U2141 ( .A(n2576), .B(\registers[2][26] ), .Z(n3067) );
  HS65_LH_NAND3X5 U2142 ( .A(n3073), .B(n3074), .C(n3075), .Z(n1079) );
  HS65_LH_NAND2X7 U2143 ( .A(n2579), .B(\registers[1][27] ), .Z(n3075) );
  HS65_LH_NAND2X7 U2144 ( .A(n2573), .B(\registers[3][27] ), .Z(n3074) );
  HS65_LH_NAND2X7 U2145 ( .A(n2576), .B(\registers[2][27] ), .Z(n3073) );
  HS65_LH_NAND3X5 U2146 ( .A(n3079), .B(n3080), .C(n3081), .Z(n1064) );
  HS65_LH_NAND2X7 U2147 ( .A(n2579), .B(\registers[1][28] ), .Z(n3081) );
  HS65_LH_NAND2X7 U2148 ( .A(n2573), .B(\registers[3][28] ), .Z(n3080) );
  HS65_LH_NAND2X7 U2149 ( .A(n2576), .B(\registers[2][28] ), .Z(n3079) );
  HS65_LH_NAND3X5 U2150 ( .A(n3085), .B(n3086), .C(n3087), .Z(n1049) );
  HS65_LH_NAND2X7 U2151 ( .A(n2579), .B(\registers[1][29] ), .Z(n3087) );
  HS65_LH_NAND2X7 U2152 ( .A(n2573), .B(\registers[3][29] ), .Z(n3086) );
  HS65_LH_NAND2X7 U2153 ( .A(n2576), .B(\registers[2][29] ), .Z(n3085) );
  HS65_LH_NAND3X5 U2154 ( .A(n3091), .B(n3092), .C(n3093), .Z(n1019) );
  HS65_LH_NAND2X7 U2155 ( .A(n2579), .B(\registers[1][30] ), .Z(n3093) );
  HS65_LH_NAND2X7 U2156 ( .A(n2573), .B(\registers[3][30] ), .Z(n3092) );
  HS65_LH_NAND2X7 U2157 ( .A(n2576), .B(\registers[2][30] ), .Z(n3091) );
  HS65_LH_NAND3X5 U2158 ( .A(n3097), .B(n3098), .C(n3099), .Z(n1004) );
  HS65_LH_NAND2X7 U2159 ( .A(n2579), .B(\registers[1][31] ), .Z(n3099) );
  HS65_LH_NAND2X7 U2160 ( .A(n2573), .B(\registers[3][31] ), .Z(n3098) );
  HS65_LH_NAND2X7 U2161 ( .A(n2576), .B(\registers[2][31] ), .Z(n3097) );
  HS65_LH_NAND2X7 U2162 ( .A(\registers[2][10] ), .B(n2667), .Z(n2968) );
  HS65_LH_NAND2X7 U2163 ( .A(\registers[3][10] ), .B(n2664), .Z(n2969) );
  HS65_LH_NAND2X7 U2164 ( .A(\registers[1][10] ), .B(n2670), .Z(n2970) );
  HS65_LH_AO22X9 U2165 ( .A(n2697), .B(n2510), .C(n2507), .D(\registers[1][0] ), .Z(n1434) );
  HS65_LH_AO22X9 U2166 ( .A(n2699), .B(n2510), .C(n2506), .D(\registers[1][1] ), .Z(n1435) );
  HS65_LH_AO22X9 U2167 ( .A(n2701), .B(n2510), .C(n2507), .D(\registers[1][2] ), .Z(n1436) );
  HS65_LH_AO22X9 U2168 ( .A(n2703), .B(n2510), .C(n2506), .D(\registers[1][3] ), .Z(n1437) );
  HS65_LH_AO22X9 U2169 ( .A(n2705), .B(n2510), .C(n2507), .D(\registers[1][4] ), .Z(n1438) );
  HS65_LH_AO22X9 U2170 ( .A(n2707), .B(n2510), .C(n2506), .D(\registers[1][5] ), .Z(n1439) );
  HS65_LH_AO22X9 U2171 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2510), .C(n2507), 
        .D(\registers[1][6] ), .Z(n1440) );
  HS65_LH_AO22X9 U2172 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2510), .C(n2507), 
        .D(\registers[1][7] ), .Z(n1441) );
  HS65_LH_AO22X9 U2173 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2510), .C(n2507), 
        .D(\registers[1][8] ), .Z(n1442) );
  HS65_LH_AO22X9 U2174 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2510), .C(n2507), 
        .D(\registers[1][9] ), .Z(n1443) );
  HS65_LH_AO22X9 U2175 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2510), .C(n2507), 
        .D(\registers[1][10] ), .Z(n1444) );
  HS65_LH_AO22X9 U2176 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2509), .C(n2507), 
        .D(\registers[1][11] ), .Z(n1445) );
  HS65_LH_AO22X9 U2177 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2509), .C(n2507), 
        .D(\registers[1][12] ), .Z(n1446) );
  HS65_LH_AO22X9 U2178 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2509), .C(n2507), 
        .D(\registers[1][13] ), .Z(n1447) );
  HS65_LH_AO22X9 U2179 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2509), .C(n2507), 
        .D(\registers[1][14] ), .Z(n1448) );
  HS65_LH_AO22X9 U2180 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2509), .C(n2507), 
        .D(\registers[1][15] ), .Z(n1449) );
  HS65_LH_AO22X9 U2181 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2509), .C(n2507), 
        .D(\registers[1][16] ), .Z(n1450) );
  HS65_LH_AO22X9 U2182 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2509), .C(n2507), 
        .D(\registers[1][17] ), .Z(n1451) );
  HS65_LH_AO22X9 U2183 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2509), .C(n2507), 
        .D(\registers[1][18] ), .Z(n1452) );
  HS65_LH_AO22X9 U2184 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2509), .C(n2506), 
        .D(\registers[1][19] ), .Z(n1453) );
  HS65_LH_AO22X9 U2185 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2509), .C(n2506), 
        .D(\registers[1][20] ), .Z(n1454) );
  HS65_LH_AO22X9 U2186 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2509), .C(n2506), 
        .D(\registers[1][21] ), .Z(n1455) );
  HS65_LH_AO22X9 U2187 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2509), .C(n2506), 
        .D(\registers[1][22] ), .Z(n1456) );
  HS65_LH_AO22X9 U2188 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2509), .C(n2506), 
        .D(\registers[1][23] ), .Z(n1457) );
  HS65_LH_AO22X9 U2189 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2509), .C(n2506), 
        .D(\registers[1][24] ), .Z(n1458) );
  HS65_LH_AO22X9 U2190 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2509), .C(n2506), 
        .D(\registers[1][25] ), .Z(n1459) );
  HS65_LH_AO22X9 U2191 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2509), .C(n2506), 
        .D(\registers[1][26] ), .Z(n1460) );
  HS65_LH_AO22X9 U2192 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2509), .C(n2506), 
        .D(\registers[1][27] ), .Z(n1461) );
  HS65_LH_AO22X9 U2193 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2509), .C(n2506), 
        .D(\registers[1][28] ), .Z(n1462) );
  HS65_LH_AO22X9 U2194 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2509), .C(n2506), 
        .D(\registers[1][29] ), .Z(n1463) );
  HS65_LH_AO22X9 U2195 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2509), .C(n2506), 
        .D(\registers[1][30] ), .Z(n1464) );
  HS65_LH_AO22X9 U2196 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2508), .C(n2506), 
        .D(\registers[1][31] ), .Z(n1465) );
  HS65_LH_AO22X9 U2197 ( .A(n2697), .B(n2505), .C(n2502), .D(\registers[2][0] ), .Z(n1466) );
  HS65_LH_AO22X9 U2198 ( .A(n2699), .B(n2505), .C(n2501), .D(\registers[2][1] ), .Z(n1467) );
  HS65_LH_AO22X9 U2199 ( .A(n2701), .B(n2505), .C(n2502), .D(\registers[2][2] ), .Z(n1468) );
  HS65_LH_AO22X9 U2200 ( .A(n2703), .B(n2505), .C(n2501), .D(\registers[2][3] ), .Z(n1469) );
  HS65_LH_AO22X9 U2201 ( .A(n2705), .B(n2505), .C(n2502), .D(\registers[2][4] ), .Z(n1470) );
  HS65_LH_AO22X9 U2202 ( .A(n2707), .B(n2505), .C(n2501), .D(\registers[2][5] ), .Z(n1471) );
  HS65_LH_AO22X9 U2203 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2505), .C(n2502), 
        .D(\registers[2][6] ), .Z(n1472) );
  HS65_LH_AO22X9 U2204 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2505), .C(n2502), 
        .D(\registers[2][7] ), .Z(n1473) );
  HS65_LH_AO22X9 U2205 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2505), .C(n2502), 
        .D(\registers[2][8] ), .Z(n1474) );
  HS65_LH_AO22X9 U2206 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2505), .C(n2502), 
        .D(\registers[2][9] ), .Z(n1475) );
  HS65_LH_AO22X9 U2207 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2505), .C(n2502), 
        .D(\registers[2][10] ), .Z(n1476) );
  HS65_LH_AO22X9 U2208 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2504), .C(n2502), 
        .D(\registers[2][11] ), .Z(n1477) );
  HS65_LH_AO22X9 U2209 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2504), .C(n2502), 
        .D(\registers[2][12] ), .Z(n1478) );
  HS65_LH_AO22X9 U2210 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2504), .C(n2502), 
        .D(\registers[2][13] ), .Z(n1479) );
  HS65_LH_AO22X9 U2211 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2504), .C(n2502), 
        .D(\registers[2][14] ), .Z(n1480) );
  HS65_LH_AO22X9 U2212 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2504), .C(n2502), 
        .D(\registers[2][15] ), .Z(n1481) );
  HS65_LH_AO22X9 U2213 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2504), .C(n2502), 
        .D(\registers[2][16] ), .Z(n1482) );
  HS65_LH_AO22X9 U2214 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2504), .C(n2502), 
        .D(\registers[2][17] ), .Z(n1483) );
  HS65_LH_AO22X9 U2215 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2504), .C(n2502), 
        .D(\registers[2][18] ), .Z(n1484) );
  HS65_LH_AO22X9 U2216 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2504), .C(n2501), 
        .D(\registers[2][19] ), .Z(n1485) );
  HS65_LH_AO22X9 U2217 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2504), .C(n2501), 
        .D(\registers[2][20] ), .Z(n1486) );
  HS65_LH_AO22X9 U2218 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2504), .C(n2501), 
        .D(\registers[2][21] ), .Z(n1487) );
  HS65_LH_AO22X9 U2219 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2504), .C(n2501), 
        .D(\registers[2][22] ), .Z(n1488) );
  HS65_LH_AO22X9 U2220 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2504), .C(n2501), 
        .D(\registers[2][23] ), .Z(n1489) );
  HS65_LH_AO22X9 U2221 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2504), .C(n2501), 
        .D(\registers[2][24] ), .Z(n1490) );
  HS65_LH_AO22X9 U2222 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2504), .C(n2501), 
        .D(\registers[2][25] ), .Z(n1491) );
  HS65_LH_AO22X9 U2223 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2504), .C(n2501), 
        .D(\registers[2][26] ), .Z(n1492) );
  HS65_LH_AO22X9 U2224 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2504), .C(n2501), 
        .D(\registers[2][27] ), .Z(n1493) );
  HS65_LH_AO22X9 U2225 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2504), .C(n2501), 
        .D(\registers[2][28] ), .Z(n1494) );
  HS65_LH_AO22X9 U2226 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2504), .C(n2501), 
        .D(\registers[2][29] ), .Z(n1495) );
  HS65_LH_AO22X9 U2227 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2504), .C(n2501), 
        .D(\registers[2][30] ), .Z(n1496) );
  HS65_LH_AO22X9 U2228 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2503), .C(n2501), 
        .D(\registers[2][31] ), .Z(n1497) );
  HS65_LH_AO22X9 U2229 ( .A(n2697), .B(n2500), .C(n2497), .D(\registers[3][0] ), .Z(n1498) );
  HS65_LH_AO22X9 U2230 ( .A(n2699), .B(n2500), .C(n2496), .D(\registers[3][1] ), .Z(n1499) );
  HS65_LH_AO22X9 U2231 ( .A(n2701), .B(n2500), .C(n2497), .D(\registers[3][2] ), .Z(n1500) );
  HS65_LH_AO22X9 U2232 ( .A(n2703), .B(n2500), .C(n2496), .D(\registers[3][3] ), .Z(n1501) );
  HS65_LH_AO22X9 U2233 ( .A(n2705), .B(n2500), .C(n2497), .D(\registers[3][4] ), .Z(n1502) );
  HS65_LH_AO22X9 U2234 ( .A(n2707), .B(n2500), .C(n2496), .D(\registers[3][5] ), .Z(n1503) );
  HS65_LH_AO22X9 U2235 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2500), .C(n2497), 
        .D(\registers[3][6] ), .Z(n1504) );
  HS65_LH_AO22X9 U2236 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2500), .C(n2497), 
        .D(\registers[3][7] ), .Z(n1505) );
  HS65_LH_AO22X9 U2237 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2500), .C(n2497), 
        .D(\registers[3][8] ), .Z(n1506) );
  HS65_LH_AO22X9 U2238 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2500), .C(n2497), 
        .D(\registers[3][9] ), .Z(n1507) );
  HS65_LH_AO22X9 U2239 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2500), .C(n2497), 
        .D(\registers[3][10] ), .Z(n1508) );
  HS65_LH_AO22X9 U2240 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2499), .C(n2497), 
        .D(\registers[3][11] ), .Z(n1509) );
  HS65_LH_AO22X9 U2241 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2499), .C(n2497), 
        .D(\registers[3][12] ), .Z(n1510) );
  HS65_LH_AO22X9 U2242 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2499), .C(n2497), 
        .D(\registers[3][13] ), .Z(n1511) );
  HS65_LH_AO22X9 U2243 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2499), .C(n2497), 
        .D(\registers[3][14] ), .Z(n1512) );
  HS65_LH_AO22X9 U2244 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2499), .C(n2497), 
        .D(\registers[3][15] ), .Z(n1513) );
  HS65_LH_AO22X9 U2245 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2499), .C(n2497), 
        .D(\registers[3][16] ), .Z(n1514) );
  HS65_LH_AO22X9 U2246 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2499), .C(n2497), 
        .D(\registers[3][17] ), .Z(n1515) );
  HS65_LH_AO22X9 U2247 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2499), .C(n2497), 
        .D(\registers[3][18] ), .Z(n1516) );
  HS65_LH_AO22X9 U2248 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2499), .C(n2496), 
        .D(\registers[3][19] ), .Z(n1517) );
  HS65_LH_AO22X9 U2249 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2499), .C(n2496), 
        .D(\registers[3][20] ), .Z(n1518) );
  HS65_LH_AO22X9 U2250 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2499), .C(n2496), 
        .D(\registers[3][21] ), .Z(n1519) );
  HS65_LH_AO22X9 U2251 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2499), .C(n2496), 
        .D(\registers[3][22] ), .Z(n1520) );
  HS65_LH_AO22X9 U2252 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2499), .C(n2496), 
        .D(\registers[3][23] ), .Z(n1521) );
  HS65_LH_AO22X9 U2253 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2499), .C(n2496), 
        .D(\registers[3][24] ), .Z(n1522) );
  HS65_LH_AO22X9 U2254 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2499), .C(n2496), 
        .D(\registers[3][25] ), .Z(n1523) );
  HS65_LH_AO22X9 U2255 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2499), .C(n2496), 
        .D(\registers[3][26] ), .Z(n1524) );
  HS65_LH_AO22X9 U2256 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2499), .C(n2496), 
        .D(\registers[3][27] ), .Z(n1525) );
  HS65_LH_AO22X9 U2257 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2499), .C(n2496), 
        .D(\registers[3][28] ), .Z(n1526) );
  HS65_LH_AO22X9 U2258 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2499), .C(n2496), 
        .D(\registers[3][29] ), .Z(n1527) );
  HS65_LH_AO22X9 U2259 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2499), .C(n2496), 
        .D(\registers[3][30] ), .Z(n1528) );
  HS65_LH_AO22X9 U2260 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2498), .C(n2496), 
        .D(\registers[3][31] ), .Z(n1529) );
  HS65_LH_AO22X9 U2261 ( .A(n2697), .B(n2460), .C(n2457), .D(
        \registers[11][0] ), .Z(n1754) );
  HS65_LH_AO22X9 U2262 ( .A(n2699), .B(n2460), .C(n2456), .D(
        \registers[11][1] ), .Z(n1755) );
  HS65_LH_AO22X9 U2263 ( .A(n2701), .B(n2460), .C(n2457), .D(
        \registers[11][2] ), .Z(n1756) );
  HS65_LH_AO22X9 U2264 ( .A(n2703), .B(n2460), .C(n2456), .D(
        \registers[11][3] ), .Z(n1757) );
  HS65_LH_AO22X9 U2265 ( .A(n2705), .B(n2460), .C(n2457), .D(
        \registers[11][4] ), .Z(n1758) );
  HS65_LH_AO22X9 U2266 ( .A(n2707), .B(n2460), .C(n2456), .D(
        \registers[11][5] ), .Z(n1759) );
  HS65_LH_AO22X9 U2267 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2460), .C(n2457), 
        .D(\registers[11][6] ), .Z(n1760) );
  HS65_LH_AO22X9 U2268 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2460), .C(n2457), 
        .D(\registers[11][7] ), .Z(n1761) );
  HS65_LH_AO22X9 U2269 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2460), .C(n2457), 
        .D(\registers[11][8] ), .Z(n1762) );
  HS65_LH_AO22X9 U2270 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2460), .C(n2457), 
        .D(\registers[11][9] ), .Z(n1763) );
  HS65_LH_AO22X9 U2271 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2460), .C(n2457), 
        .D(\registers[11][10] ), .Z(n1764) );
  HS65_LH_AO22X9 U2272 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2459), .C(n2457), 
        .D(\registers[11][11] ), .Z(n1765) );
  HS65_LH_AO22X9 U2273 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2459), .C(n2457), 
        .D(\registers[11][12] ), .Z(n1766) );
  HS65_LH_AO22X9 U2274 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2459), .C(n2457), 
        .D(\registers[11][13] ), .Z(n1767) );
  HS65_LH_AO22X9 U2275 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2459), .C(n2457), 
        .D(\registers[11][14] ), .Z(n1768) );
  HS65_LH_AO22X9 U2276 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2459), .C(n2457), 
        .D(\registers[11][15] ), .Z(n1769) );
  HS65_LH_AO22X9 U2277 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2459), .C(n2457), 
        .D(\registers[11][16] ), .Z(n1770) );
  HS65_LH_AO22X9 U2278 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2459), .C(n2457), 
        .D(\registers[11][17] ), .Z(n1771) );
  HS65_LH_AO22X9 U2279 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2459), .C(n2457), 
        .D(\registers[11][18] ), .Z(n1772) );
  HS65_LH_AO22X9 U2280 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2459), .C(n2456), 
        .D(\registers[11][19] ), .Z(n1773) );
  HS65_LH_AO22X9 U2281 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2459), .C(n2456), 
        .D(\registers[11][20] ), .Z(n1774) );
  HS65_LH_AO22X9 U2282 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2459), .C(n2456), 
        .D(\registers[11][21] ), .Z(n1775) );
  HS65_LH_AO22X9 U2283 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2459), .C(n2456), 
        .D(\registers[11][22] ), .Z(n1776) );
  HS65_LH_AO22X9 U2284 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2459), .C(n2456), 
        .D(\registers[11][23] ), .Z(n1777) );
  HS65_LH_AO22X9 U2285 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2459), .C(n2456), 
        .D(\registers[11][24] ), .Z(n1778) );
  HS65_LH_AO22X9 U2286 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2459), .C(n2456), 
        .D(\registers[11][25] ), .Z(n1779) );
  HS65_LH_AO22X9 U2287 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2459), .C(n2456), 
        .D(\registers[11][26] ), .Z(n1780) );
  HS65_LH_AO22X9 U2288 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2459), .C(n2456), 
        .D(\registers[11][27] ), .Z(n1781) );
  HS65_LH_AO22X9 U2289 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2459), .C(n2456), 
        .D(\registers[11][28] ), .Z(n1782) );
  HS65_LH_AO22X9 U2290 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2459), .C(n2456), 
        .D(\registers[11][29] ), .Z(n1783) );
  HS65_LH_AO22X9 U2291 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2459), .C(n2456), 
        .D(\registers[11][30] ), .Z(n1784) );
  HS65_LH_AO22X9 U2292 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2458), .C(n2456), 
        .D(\registers[11][31] ), .Z(n1785) );
  HS65_LH_AO22X9 U2293 ( .A(n2697), .B(n2450), .C(n2447), .D(
        \registers[13][0] ), .Z(n1818) );
  HS65_LH_AO22X9 U2294 ( .A(n2699), .B(n2450), .C(n2446), .D(
        \registers[13][1] ), .Z(n1819) );
  HS65_LH_AO22X9 U2295 ( .A(n2701), .B(n2450), .C(n2447), .D(
        \registers[13][2] ), .Z(n1820) );
  HS65_LH_AO22X9 U2296 ( .A(n2703), .B(n2450), .C(n2446), .D(
        \registers[13][3] ), .Z(n1821) );
  HS65_LH_AO22X9 U2297 ( .A(n2705), .B(n2450), .C(n2447), .D(
        \registers[13][4] ), .Z(n1822) );
  HS65_LH_AO22X9 U2298 ( .A(n2707), .B(n2450), .C(n2446), .D(
        \registers[13][5] ), .Z(n1823) );
  HS65_LH_AO22X9 U2299 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2450), .C(n2447), 
        .D(\registers[13][6] ), .Z(n1824) );
  HS65_LH_AO22X9 U2300 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2450), .C(n2447), 
        .D(\registers[13][7] ), .Z(n1825) );
  HS65_LH_AO22X9 U2301 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2450), .C(n2447), 
        .D(\registers[13][8] ), .Z(n1826) );
  HS65_LH_AO22X9 U2302 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2450), .C(n2447), 
        .D(\registers[13][9] ), .Z(n1827) );
  HS65_LH_AO22X9 U2303 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2450), .C(n2447), 
        .D(\registers[13][10] ), .Z(n1828) );
  HS65_LH_AO22X9 U2304 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2449), .C(n2447), 
        .D(\registers[13][11] ), .Z(n1829) );
  HS65_LH_AO22X9 U2305 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2449), .C(n2447), 
        .D(\registers[13][12] ), .Z(n1830) );
  HS65_LH_AO22X9 U2306 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2449), .C(n2447), 
        .D(\registers[13][13] ), .Z(n1831) );
  HS65_LH_AO22X9 U2307 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2449), .C(n2447), 
        .D(\registers[13][14] ), .Z(n1832) );
  HS65_LH_AO22X9 U2308 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2449), .C(n2447), 
        .D(\registers[13][15] ), .Z(n1833) );
  HS65_LH_AO22X9 U2309 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2449), .C(n2447), 
        .D(\registers[13][16] ), .Z(n1834) );
  HS65_LH_AO22X9 U2310 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2449), .C(n2447), 
        .D(\registers[13][17] ), .Z(n1835) );
  HS65_LH_AO22X9 U2311 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2449), .C(n2447), 
        .D(\registers[13][18] ), .Z(n1836) );
  HS65_LH_AO22X9 U2312 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2449), .C(n2446), 
        .D(\registers[13][19] ), .Z(n1837) );
  HS65_LH_AO22X9 U2313 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2449), .C(n2446), 
        .D(\registers[13][20] ), .Z(n1838) );
  HS65_LH_AO22X9 U2314 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2449), .C(n2446), 
        .D(\registers[13][21] ), .Z(n1839) );
  HS65_LH_AO22X9 U2315 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2449), .C(n2446), 
        .D(\registers[13][22] ), .Z(n1840) );
  HS65_LH_AO22X9 U2316 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2449), .C(n2446), 
        .D(\registers[13][23] ), .Z(n1841) );
  HS65_LH_AO22X9 U2317 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2449), .C(n2446), 
        .D(\registers[13][24] ), .Z(n1842) );
  HS65_LH_AO22X9 U2318 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2449), .C(n2446), 
        .D(\registers[13][25] ), .Z(n1843) );
  HS65_LH_AO22X9 U2319 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2449), .C(n2446), 
        .D(\registers[13][26] ), .Z(n1844) );
  HS65_LH_AO22X9 U2320 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2449), .C(n2446), 
        .D(\registers[13][27] ), .Z(n1845) );
  HS65_LH_AO22X9 U2321 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2449), .C(n2446), 
        .D(\registers[13][28] ), .Z(n1846) );
  HS65_LH_AO22X9 U2322 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2449), .C(n2446), 
        .D(\registers[13][29] ), .Z(n1847) );
  HS65_LH_AO22X9 U2323 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2449), .C(n2446), 
        .D(\registers[13][30] ), .Z(n1848) );
  HS65_LH_AO22X9 U2324 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2448), .C(n2446), 
        .D(\registers[13][31] ), .Z(n1849) );
  HS65_LH_AO22X9 U2325 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n322), .C(n319), 
        .D(\registers[25][0] ), .Z(n2202) );
  HS65_LH_AO22X9 U2326 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n322), .C(n318), 
        .D(\registers[25][1] ), .Z(n2203) );
  HS65_LH_AO22X9 U2327 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n322), .C(n319), 
        .D(\registers[25][2] ), .Z(n2204) );
  HS65_LH_AO22X9 U2328 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n322), .C(n318), 
        .D(\registers[25][3] ), .Z(n2205) );
  HS65_LH_AO22X9 U2329 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n322), .C(n319), 
        .D(\registers[25][4] ), .Z(n2206) );
  HS65_LH_AO22X9 U2330 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n322), .C(n318), 
        .D(\registers[25][5] ), .Z(n2207) );
  HS65_LH_AO22X9 U2331 ( .A(n2709), .B(n322), .C(n319), .D(\registers[25][6] ), 
        .Z(n2208) );
  HS65_LH_AO22X9 U2332 ( .A(n2711), .B(n322), .C(n319), .D(\registers[25][7] ), 
        .Z(n2209) );
  HS65_LH_AO22X9 U2333 ( .A(n2713), .B(n322), .C(n319), .D(\registers[25][8] ), 
        .Z(n2210) );
  HS65_LH_AO22X9 U2334 ( .A(n2715), .B(n322), .C(n319), .D(\registers[25][9] ), 
        .Z(n2211) );
  HS65_LH_AO22X9 U2335 ( .A(n2717), .B(n322), .C(n319), .D(\registers[25][10] ), .Z(n2212) );
  HS65_LH_AO22X9 U2336 ( .A(n2719), .B(n321), .C(n319), .D(\registers[25][11] ), .Z(n2213) );
  HS65_LH_AO22X9 U2337 ( .A(n2721), .B(n321), .C(n319), .D(\registers[25][12] ), .Z(n2214) );
  HS65_LH_AO22X9 U2338 ( .A(n2723), .B(n321), .C(n319), .D(\registers[25][13] ), .Z(n2215) );
  HS65_LH_AO22X9 U2339 ( .A(n2725), .B(n321), .C(n319), .D(\registers[25][14] ), .Z(n2216) );
  HS65_LH_AO22X9 U2340 ( .A(n2727), .B(n321), .C(n319), .D(\registers[25][15] ), .Z(n2217) );
  HS65_LH_AO22X9 U2341 ( .A(n2729), .B(n321), .C(n319), .D(\registers[25][16] ), .Z(n2218) );
  HS65_LH_AO22X9 U2342 ( .A(n2731), .B(n321), .C(n319), .D(\registers[25][17] ), .Z(n2219) );
  HS65_LH_AO22X9 U2343 ( .A(n2733), .B(n321), .C(n319), .D(\registers[25][18] ), .Z(n2220) );
  HS65_LH_AO22X9 U2344 ( .A(n2735), .B(n321), .C(n318), .D(\registers[25][19] ), .Z(n2221) );
  HS65_LH_AO22X9 U2345 ( .A(n2737), .B(n321), .C(n318), .D(\registers[25][20] ), .Z(n2222) );
  HS65_LH_AO22X9 U2346 ( .A(n2739), .B(n321), .C(n318), .D(\registers[25][21] ), .Z(n2223) );
  HS65_LH_AO22X9 U2347 ( .A(n2741), .B(n321), .C(n318), .D(\registers[25][22] ), .Z(n2224) );
  HS65_LH_AO22X9 U2348 ( .A(n2743), .B(n321), .C(n318), .D(\registers[25][23] ), .Z(n2225) );
  HS65_LH_AO22X9 U2349 ( .A(n2745), .B(n321), .C(n318), .D(\registers[25][24] ), .Z(n2226) );
  HS65_LH_AO22X9 U2350 ( .A(n2747), .B(n321), .C(n318), .D(\registers[25][25] ), .Z(n2227) );
  HS65_LH_AO22X9 U2351 ( .A(n2749), .B(n321), .C(n318), .D(\registers[25][26] ), .Z(n2228) );
  HS65_LH_AO22X9 U2352 ( .A(n2751), .B(n321), .C(n318), .D(\registers[25][27] ), .Z(n2229) );
  HS65_LH_AO22X9 U2353 ( .A(n2753), .B(n321), .C(n318), .D(\registers[25][28] ), .Z(n2230) );
  HS65_LH_AO22X9 U2354 ( .A(n2755), .B(n321), .C(n318), .D(\registers[25][29] ), .Z(n2231) );
  HS65_LH_AO22X9 U2355 ( .A(n2757), .B(n321), .C(n318), .D(\registers[25][30] ), .Z(n2232) );
  HS65_LH_AO22X9 U2356 ( .A(n2759), .B(n320), .C(n318), .D(\registers[25][31] ), .Z(n2233) );
  HS65_LH_AO22X9 U2357 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n292), .C(n289), 
        .D(\registers[31][0] ), .Z(n2394) );
  HS65_LH_AO22X9 U2358 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n292), .C(n288), 
        .D(\registers[31][1] ), .Z(n2395) );
  HS65_LH_AO22X9 U2359 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n292), .C(n289), 
        .D(\registers[31][2] ), .Z(n2396) );
  HS65_LH_AO22X9 U2360 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n292), .C(n288), 
        .D(\registers[31][3] ), .Z(n2397) );
  HS65_LH_AO22X9 U2361 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n292), .C(n289), 
        .D(\registers[31][4] ), .Z(n2398) );
  HS65_LH_AO22X9 U2362 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n292), .C(n288), 
        .D(\registers[31][5] ), .Z(n2399) );
  HS65_LH_AO22X9 U2363 ( .A(n2709), .B(n292), .C(n289), .D(\registers[31][6] ), 
        .Z(n2400) );
  HS65_LH_AO22X9 U2364 ( .A(n2711), .B(n292), .C(n289), .D(\registers[31][7] ), 
        .Z(n2401) );
  HS65_LH_AO22X9 U2365 ( .A(n2713), .B(n292), .C(n289), .D(\registers[31][8] ), 
        .Z(n2402) );
  HS65_LH_AO22X9 U2366 ( .A(n2715), .B(n292), .C(n289), .D(\registers[31][9] ), 
        .Z(n2403) );
  HS65_LH_AO22X9 U2367 ( .A(n2717), .B(n292), .C(n289), .D(\registers[31][10] ), .Z(n2404) );
  HS65_LH_AO22X9 U2368 ( .A(n2719), .B(n291), .C(n289), .D(\registers[31][11] ), .Z(n2405) );
  HS65_LH_AO22X9 U2369 ( .A(n2721), .B(n291), .C(n289), .D(\registers[31][12] ), .Z(n2406) );
  HS65_LH_AO22X9 U2370 ( .A(n2723), .B(n291), .C(n289), .D(\registers[31][13] ), .Z(n2407) );
  HS65_LH_AO22X9 U2371 ( .A(n2725), .B(n291), .C(n289), .D(\registers[31][14] ), .Z(n2408) );
  HS65_LH_AO22X9 U2372 ( .A(n2727), .B(n291), .C(n289), .D(\registers[31][15] ), .Z(n2409) );
  HS65_LH_AO22X9 U2373 ( .A(n2729), .B(n291), .C(n289), .D(\registers[31][16] ), .Z(n2410) );
  HS65_LH_AO22X9 U2374 ( .A(n2731), .B(n291), .C(n289), .D(\registers[31][17] ), .Z(n2411) );
  HS65_LH_AO22X9 U2375 ( .A(n2733), .B(n291), .C(n289), .D(\registers[31][18] ), .Z(n2412) );
  HS65_LH_AO22X9 U2376 ( .A(n2735), .B(n291), .C(n288), .D(\registers[31][19] ), .Z(n2413) );
  HS65_LH_AO22X9 U2377 ( .A(n2737), .B(n291), .C(n288), .D(\registers[31][20] ), .Z(n2414) );
  HS65_LH_AO22X9 U2378 ( .A(n2739), .B(n291), .C(n288), .D(\registers[31][21] ), .Z(n2415) );
  HS65_LH_AO22X9 U2379 ( .A(n2741), .B(n291), .C(n288), .D(\registers[31][22] ), .Z(n2416) );
  HS65_LH_AO22X9 U2380 ( .A(n2743), .B(n291), .C(n288), .D(\registers[31][23] ), .Z(n2417) );
  HS65_LH_AO22X9 U2381 ( .A(n2745), .B(n291), .C(n288), .D(\registers[31][24] ), .Z(n2418) );
  HS65_LH_AO22X9 U2382 ( .A(n2747), .B(n291), .C(n288), .D(\registers[31][25] ), .Z(n2419) );
  HS65_LH_AO22X9 U2383 ( .A(n2749), .B(n291), .C(n288), .D(\registers[31][26] ), .Z(n2420) );
  HS65_LH_AO22X9 U2384 ( .A(n2751), .B(n291), .C(n288), .D(\registers[31][27] ), .Z(n2421) );
  HS65_LH_AO22X9 U2385 ( .A(n2753), .B(n291), .C(n288), .D(\registers[31][28] ), .Z(n2422) );
  HS65_LH_AO22X9 U2386 ( .A(n2755), .B(n291), .C(n288), .D(\registers[31][29] ), .Z(n2423) );
  HS65_LH_AO22X9 U2387 ( .A(n2757), .B(n291), .C(n288), .D(\registers[31][30] ), .Z(n2424) );
  HS65_LH_AO22X9 U2388 ( .A(n2759), .B(n290), .C(n288), .D(\registers[31][31] ), .Z(n2425) );
  HS65_LH_AO22X9 U2389 ( .A(n2697), .B(n2465), .C(n2462), .D(
        \registers[10][0] ), .Z(n1722) );
  HS65_LH_AO22X9 U2390 ( .A(n2699), .B(n2465), .C(n2461), .D(
        \registers[10][1] ), .Z(n1723) );
  HS65_LH_AO22X9 U2391 ( .A(n2701), .B(n2465), .C(n2462), .D(
        \registers[10][2] ), .Z(n1724) );
  HS65_LH_AO22X9 U2392 ( .A(n2703), .B(n2465), .C(n2461), .D(
        \registers[10][3] ), .Z(n1725) );
  HS65_LH_AO22X9 U2393 ( .A(n2705), .B(n2465), .C(n2462), .D(
        \registers[10][4] ), .Z(n1726) );
  HS65_LH_AO22X9 U2394 ( .A(n2707), .B(n2465), .C(n2461), .D(
        \registers[10][5] ), .Z(n1727) );
  HS65_LH_AO22X9 U2395 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2465), .C(n2462), 
        .D(\registers[10][6] ), .Z(n1728) );
  HS65_LH_AO22X9 U2396 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2465), .C(n2462), 
        .D(\registers[10][7] ), .Z(n1729) );
  HS65_LH_AO22X9 U2397 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2465), .C(n2462), 
        .D(\registers[10][8] ), .Z(n1730) );
  HS65_LH_AO22X9 U2398 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2465), .C(n2462), 
        .D(\registers[10][9] ), .Z(n1731) );
  HS65_LH_AO22X9 U2399 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2465), .C(n2462), 
        .D(\registers[10][10] ), .Z(n1732) );
  HS65_LH_AO22X9 U2400 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2464), .C(n2462), 
        .D(\registers[10][11] ), .Z(n1733) );
  HS65_LH_AO22X9 U2401 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2464), .C(n2462), 
        .D(\registers[10][12] ), .Z(n1734) );
  HS65_LH_AO22X9 U2402 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2464), .C(n2462), 
        .D(\registers[10][13] ), .Z(n1735) );
  HS65_LH_AO22X9 U2403 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2464), .C(n2462), 
        .D(\registers[10][14] ), .Z(n1736) );
  HS65_LH_AO22X9 U2404 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2464), .C(n2462), 
        .D(\registers[10][15] ), .Z(n1737) );
  HS65_LH_AO22X9 U2405 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2464), .C(n2462), 
        .D(\registers[10][16] ), .Z(n1738) );
  HS65_LH_AO22X9 U2406 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2464), .C(n2462), 
        .D(\registers[10][17] ), .Z(n1739) );
  HS65_LH_AO22X9 U2407 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2464), .C(n2462), 
        .D(\registers[10][18] ), .Z(n1740) );
  HS65_LH_AO22X9 U2408 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2464), .C(n2461), 
        .D(\registers[10][19] ), .Z(n1741) );
  HS65_LH_AO22X9 U2409 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2464), .C(n2461), 
        .D(\registers[10][20] ), .Z(n1742) );
  HS65_LH_AO22X9 U2410 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2464), .C(n2461), 
        .D(\registers[10][21] ), .Z(n1743) );
  HS65_LH_AO22X9 U2411 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2464), .C(n2461), 
        .D(\registers[10][22] ), .Z(n1744) );
  HS65_LH_AO22X9 U2412 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2464), .C(n2461), 
        .D(\registers[10][23] ), .Z(n1745) );
  HS65_LH_AO22X9 U2413 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2464), .C(n2461), 
        .D(\registers[10][24] ), .Z(n1746) );
  HS65_LH_AO22X9 U2414 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2464), .C(n2461), 
        .D(\registers[10][25] ), .Z(n1747) );
  HS65_LH_AO22X9 U2415 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2464), .C(n2461), 
        .D(\registers[10][26] ), .Z(n1748) );
  HS65_LH_AO22X9 U2416 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2464), .C(n2461), 
        .D(\registers[10][27] ), .Z(n1749) );
  HS65_LH_AO22X9 U2417 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2464), .C(n2461), 
        .D(\registers[10][28] ), .Z(n1750) );
  HS65_LH_AO22X9 U2418 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2464), .C(n2461), 
        .D(\registers[10][29] ), .Z(n1751) );
  HS65_LH_AO22X9 U2419 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2464), .C(n2461), 
        .D(\registers[10][30] ), .Z(n1752) );
  HS65_LH_AO22X9 U2420 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2463), .C(n2461), 
        .D(\registers[10][31] ), .Z(n1753) );
  HS65_LH_AO22X9 U2421 ( .A(n2697), .B(n2455), .C(n2452), .D(
        \registers[12][0] ), .Z(n1786) );
  HS65_LH_AO22X9 U2422 ( .A(n2699), .B(n2455), .C(n2451), .D(
        \registers[12][1] ), .Z(n1787) );
  HS65_LH_AO22X9 U2423 ( .A(n2701), .B(n2455), .C(n2452), .D(
        \registers[12][2] ), .Z(n1788) );
  HS65_LH_AO22X9 U2424 ( .A(n2703), .B(n2455), .C(n2451), .D(
        \registers[12][3] ), .Z(n1789) );
  HS65_LH_AO22X9 U2425 ( .A(n2705), .B(n2455), .C(n2452), .D(
        \registers[12][4] ), .Z(n1790) );
  HS65_LH_AO22X9 U2426 ( .A(n2707), .B(n2455), .C(n2451), .D(
        \registers[12][5] ), .Z(n1791) );
  HS65_LH_AO22X9 U2427 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2455), .C(n2452), 
        .D(\registers[12][6] ), .Z(n1792) );
  HS65_LH_AO22X9 U2428 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2455), .C(n2452), 
        .D(\registers[12][7] ), .Z(n1793) );
  HS65_LH_AO22X9 U2429 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2455), .C(n2452), 
        .D(\registers[12][8] ), .Z(n1794) );
  HS65_LH_AO22X9 U2430 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2455), .C(n2452), 
        .D(\registers[12][9] ), .Z(n1795) );
  HS65_LH_AO22X9 U2431 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2455), .C(n2452), 
        .D(\registers[12][10] ), .Z(n1796) );
  HS65_LH_AO22X9 U2432 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2454), .C(n2452), 
        .D(\registers[12][11] ), .Z(n1797) );
  HS65_LH_AO22X9 U2433 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2454), .C(n2452), 
        .D(\registers[12][12] ), .Z(n1798) );
  HS65_LH_AO22X9 U2434 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2454), .C(n2452), 
        .D(\registers[12][13] ), .Z(n1799) );
  HS65_LH_AO22X9 U2435 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2454), .C(n2452), 
        .D(\registers[12][14] ), .Z(n1800) );
  HS65_LH_AO22X9 U2436 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2454), .C(n2452), 
        .D(\registers[12][15] ), .Z(n1801) );
  HS65_LH_AO22X9 U2437 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2454), .C(n2452), 
        .D(\registers[12][16] ), .Z(n1802) );
  HS65_LH_AO22X9 U2438 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2454), .C(n2452), 
        .D(\registers[12][17] ), .Z(n1803) );
  HS65_LH_AO22X9 U2439 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2454), .C(n2452), 
        .D(\registers[12][18] ), .Z(n1804) );
  HS65_LH_AO22X9 U2440 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2454), .C(n2451), 
        .D(\registers[12][19] ), .Z(n1805) );
  HS65_LH_AO22X9 U2441 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2454), .C(n2451), 
        .D(\registers[12][20] ), .Z(n1806) );
  HS65_LH_AO22X9 U2442 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2454), .C(n2451), 
        .D(\registers[12][21] ), .Z(n1807) );
  HS65_LH_AO22X9 U2443 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2454), .C(n2451), 
        .D(\registers[12][22] ), .Z(n1808) );
  HS65_LH_AO22X9 U2444 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2454), .C(n2451), 
        .D(\registers[12][23] ), .Z(n1809) );
  HS65_LH_AO22X9 U2445 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2454), .C(n2451), 
        .D(\registers[12][24] ), .Z(n1810) );
  HS65_LH_AO22X9 U2446 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2454), .C(n2451), 
        .D(\registers[12][25] ), .Z(n1811) );
  HS65_LH_AO22X9 U2447 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2454), .C(n2451), 
        .D(\registers[12][26] ), .Z(n1812) );
  HS65_LH_AO22X9 U2448 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2454), .C(n2451), 
        .D(\registers[12][27] ), .Z(n1813) );
  HS65_LH_AO22X9 U2449 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2454), .C(n2451), 
        .D(\registers[12][28] ), .Z(n1814) );
  HS65_LH_AO22X9 U2450 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2454), .C(n2451), 
        .D(\registers[12][29] ), .Z(n1815) );
  HS65_LH_AO22X9 U2451 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2454), .C(n2451), 
        .D(\registers[12][30] ), .Z(n1816) );
  HS65_LH_AO22X9 U2452 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2453), .C(n2451), 
        .D(\registers[12][31] ), .Z(n1817) );
  HS65_LH_AO22X9 U2453 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n326), .C(n323), 
        .D(\registers[24][0] ), .Z(n2170) );
  HS65_LH_AO22X9 U2454 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n326), .C(n323), 
        .D(\registers[24][1] ), .Z(n2171) );
  HS65_LH_AO22X9 U2455 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n326), .C(n323), 
        .D(\registers[24][2] ), .Z(n2172) );
  HS65_LH_AO22X9 U2456 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n326), .C(n323), 
        .D(\registers[24][3] ), .Z(n2173) );
  HS65_LH_AO22X9 U2457 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n326), .C(n323), 
        .D(\registers[24][4] ), .Z(n2174) );
  HS65_LH_AO22X9 U2458 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n326), .C(n323), 
        .D(\registers[24][5] ), .Z(n2175) );
  HS65_LH_AO22X9 U2459 ( .A(n2709), .B(n326), .C(n323), .D(\registers[24][6] ), 
        .Z(n2176) );
  HS65_LH_AO22X9 U2460 ( .A(n2711), .B(n326), .C(n323), .D(\registers[24][7] ), 
        .Z(n2177) );
  HS65_LH_AO22X9 U2461 ( .A(n2713), .B(n326), .C(n323), .D(\registers[24][8] ), 
        .Z(n2178) );
  HS65_LH_AO22X9 U2462 ( .A(n2715), .B(n326), .C(n323), .D(\registers[24][9] ), 
        .Z(n2179) );
  HS65_LH_AO22X9 U2463 ( .A(n2717), .B(n326), .C(n323), .D(\registers[24][10] ), .Z(n2180) );
  HS65_LH_AO22X9 U2464 ( .A(n2719), .B(n325), .C(n323), .D(\registers[24][11] ), .Z(n2181) );
  HS65_LH_AO22X9 U2465 ( .A(n2721), .B(n325), .C(n323), .D(\registers[24][12] ), .Z(n2182) );
  HS65_LH_AO22X9 U2466 ( .A(n2723), .B(n325), .C(n323), .D(\registers[24][13] ), .Z(n2183) );
  HS65_LH_AO22X9 U2467 ( .A(n2725), .B(n325), .C(n323), .D(\registers[24][14] ), .Z(n2184) );
  HS65_LH_AO22X9 U2468 ( .A(n2727), .B(n325), .C(n323), .D(\registers[24][15] ), .Z(n2185) );
  HS65_LH_AO22X9 U2469 ( .A(n2729), .B(n325), .C(n323), .D(\registers[24][16] ), .Z(n2186) );
  HS65_LH_AO22X9 U2470 ( .A(n2731), .B(n325), .C(n323), .D(\registers[24][17] ), .Z(n2187) );
  HS65_LH_AO22X9 U2471 ( .A(n2733), .B(n325), .C(n323), .D(\registers[24][18] ), .Z(n2188) );
  HS65_LH_AO22X9 U2472 ( .A(n2735), .B(n325), .C(n323), .D(\registers[24][19] ), .Z(n2189) );
  HS65_LH_AO22X9 U2473 ( .A(n2737), .B(n325), .C(n1425), .D(
        \registers[24][20] ), .Z(n2190) );
  HS65_LH_AO22X9 U2474 ( .A(n2739), .B(n325), .C(n1425), .D(
        \registers[24][21] ), .Z(n2191) );
  HS65_LH_AO22X9 U2475 ( .A(n2741), .B(n325), .C(n1425), .D(
        \registers[24][22] ), .Z(n2192) );
  HS65_LH_AO22X9 U2476 ( .A(n2743), .B(n325), .C(n1425), .D(
        \registers[24][23] ), .Z(n2193) );
  HS65_LH_AO22X9 U2477 ( .A(n2745), .B(n325), .C(n1425), .D(
        \registers[24][24] ), .Z(n2194) );
  HS65_LH_AO22X9 U2478 ( .A(n2747), .B(n325), .C(n1425), .D(
        \registers[24][25] ), .Z(n2195) );
  HS65_LH_AO22X9 U2479 ( .A(n2749), .B(n325), .C(n1425), .D(
        \registers[24][26] ), .Z(n2196) );
  HS65_LH_AO22X9 U2480 ( .A(n2751), .B(n325), .C(n1425), .D(
        \registers[24][27] ), .Z(n2197) );
  HS65_LH_AO22X9 U2481 ( .A(n2753), .B(n325), .C(n1425), .D(
        \registers[24][28] ), .Z(n2198) );
  HS65_LH_AO22X9 U2482 ( .A(n2755), .B(n325), .C(n1425), .D(
        \registers[24][29] ), .Z(n2199) );
  HS65_LH_AO22X9 U2483 ( .A(n2757), .B(n325), .C(n1425), .D(
        \registers[24][30] ), .Z(n2200) );
  HS65_LH_AO22X9 U2484 ( .A(n2759), .B(n324), .C(n1425), .D(
        \registers[24][31] ), .Z(n2201) );
  HS65_LH_AO22X9 U2485 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n297), .C(n294), 
        .D(\registers[30][0] ), .Z(n2362) );
  HS65_LH_AO22X9 U2486 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n297), .C(n293), 
        .D(\registers[30][1] ), .Z(n2363) );
  HS65_LH_AO22X9 U2487 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n297), .C(n294), 
        .D(\registers[30][2] ), .Z(n2364) );
  HS65_LH_AO22X9 U2488 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n297), .C(n293), 
        .D(\registers[30][3] ), .Z(n2365) );
  HS65_LH_AO22X9 U2489 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n297), .C(n294), 
        .D(\registers[30][4] ), .Z(n2366) );
  HS65_LH_AO22X9 U2490 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n297), .C(n293), 
        .D(\registers[30][5] ), .Z(n2367) );
  HS65_LH_AO22X9 U2491 ( .A(n2709), .B(n297), .C(n294), .D(\registers[30][6] ), 
        .Z(n2368) );
  HS65_LH_AO22X9 U2492 ( .A(n2711), .B(n297), .C(n294), .D(\registers[30][7] ), 
        .Z(n2369) );
  HS65_LH_AO22X9 U2493 ( .A(n2713), .B(n297), .C(n294), .D(\registers[30][8] ), 
        .Z(n2370) );
  HS65_LH_AO22X9 U2494 ( .A(n2715), .B(n297), .C(n294), .D(\registers[30][9] ), 
        .Z(n2371) );
  HS65_LH_AO22X9 U2495 ( .A(n2717), .B(n297), .C(n294), .D(\registers[30][10] ), .Z(n2372) );
  HS65_LH_AO22X9 U2496 ( .A(n2719), .B(n296), .C(n294), .D(\registers[30][11] ), .Z(n2373) );
  HS65_LH_AO22X9 U2497 ( .A(n2721), .B(n296), .C(n294), .D(\registers[30][12] ), .Z(n2374) );
  HS65_LH_AO22X9 U2498 ( .A(n2723), .B(n296), .C(n294), .D(\registers[30][13] ), .Z(n2375) );
  HS65_LH_AO22X9 U2499 ( .A(n2725), .B(n296), .C(n294), .D(\registers[30][14] ), .Z(n2376) );
  HS65_LH_AO22X9 U2500 ( .A(n2727), .B(n296), .C(n294), .D(\registers[30][15] ), .Z(n2377) );
  HS65_LH_AO22X9 U2501 ( .A(n2729), .B(n296), .C(n294), .D(\registers[30][16] ), .Z(n2378) );
  HS65_LH_AO22X9 U2502 ( .A(n2731), .B(n296), .C(n294), .D(\registers[30][17] ), .Z(n2379) );
  HS65_LH_AO22X9 U2503 ( .A(n2733), .B(n296), .C(n294), .D(\registers[30][18] ), .Z(n2380) );
  HS65_LH_AO22X9 U2504 ( .A(n2735), .B(n296), .C(n293), .D(\registers[30][19] ), .Z(n2381) );
  HS65_LH_AO22X9 U2505 ( .A(n2737), .B(n296), .C(n293), .D(\registers[30][20] ), .Z(n2382) );
  HS65_LH_AO22X9 U2506 ( .A(n2739), .B(n296), .C(n293), .D(\registers[30][21] ), .Z(n2383) );
  HS65_LH_AO22X9 U2507 ( .A(n2741), .B(n296), .C(n293), .D(\registers[30][22] ), .Z(n2384) );
  HS65_LH_AO22X9 U2508 ( .A(n2743), .B(n296), .C(n293), .D(\registers[30][23] ), .Z(n2385) );
  HS65_LH_AO22X9 U2509 ( .A(n2745), .B(n296), .C(n293), .D(\registers[30][24] ), .Z(n2386) );
  HS65_LH_AO22X9 U2510 ( .A(n2747), .B(n296), .C(n293), .D(\registers[30][25] ), .Z(n2387) );
  HS65_LH_AO22X9 U2511 ( .A(n2749), .B(n296), .C(n293), .D(\registers[30][26] ), .Z(n2388) );
  HS65_LH_AO22X9 U2512 ( .A(n2751), .B(n296), .C(n293), .D(\registers[30][27] ), .Z(n2389) );
  HS65_LH_AO22X9 U2513 ( .A(n2753), .B(n296), .C(n293), .D(\registers[30][28] ), .Z(n2390) );
  HS65_LH_AO22X9 U2514 ( .A(n2755), .B(n296), .C(n293), .D(\registers[30][29] ), .Z(n2391) );
  HS65_LH_AO22X9 U2515 ( .A(n2757), .B(n296), .C(n293), .D(\registers[30][30] ), .Z(n2392) );
  HS65_LH_AO22X9 U2516 ( .A(n2759), .B(n295), .C(n293), .D(\registers[30][31] ), .Z(n2393) );
  HS65_LH_AO22X9 U2517 ( .A(n2697), .B(n2480), .C(n2477), .D(\registers[7][0] ), .Z(n1626) );
  HS65_LH_AO22X9 U2518 ( .A(n2699), .B(n2480), .C(n2476), .D(\registers[7][1] ), .Z(n1627) );
  HS65_LH_AO22X9 U2519 ( .A(n2701), .B(n2480), .C(n2477), .D(\registers[7][2] ), .Z(n1628) );
  HS65_LH_AO22X9 U2520 ( .A(n2703), .B(n2480), .C(n2476), .D(\registers[7][3] ), .Z(n1629) );
  HS65_LH_AO22X9 U2521 ( .A(n2705), .B(n2480), .C(n2477), .D(\registers[7][4] ), .Z(n1630) );
  HS65_LH_AO22X9 U2522 ( .A(n2707), .B(n2480), .C(n2476), .D(\registers[7][5] ), .Z(n1631) );
  HS65_LH_AO22X9 U2523 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2480), .C(n2477), 
        .D(\registers[7][6] ), .Z(n1632) );
  HS65_LH_AO22X9 U2524 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2480), .C(n2477), 
        .D(\registers[7][7] ), .Z(n1633) );
  HS65_LH_AO22X9 U2525 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2480), .C(n2477), 
        .D(\registers[7][8] ), .Z(n1634) );
  HS65_LH_AO22X9 U2526 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2480), .C(n2477), 
        .D(\registers[7][9] ), .Z(n1635) );
  HS65_LH_AO22X9 U2527 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2480), .C(n2477), 
        .D(\registers[7][10] ), .Z(n1636) );
  HS65_LH_AO22X9 U2528 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2479), .C(n2477), 
        .D(\registers[7][11] ), .Z(n1637) );
  HS65_LH_AO22X9 U2529 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2479), .C(n2477), 
        .D(\registers[7][12] ), .Z(n1638) );
  HS65_LH_AO22X9 U2530 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2479), .C(n2477), 
        .D(\registers[7][13] ), .Z(n1639) );
  HS65_LH_AO22X9 U2531 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2479), .C(n2477), 
        .D(\registers[7][14] ), .Z(n1640) );
  HS65_LH_AO22X9 U2532 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2479), .C(n2477), 
        .D(\registers[7][15] ), .Z(n1641) );
  HS65_LH_AO22X9 U2533 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2479), .C(n2477), 
        .D(\registers[7][16] ), .Z(n1642) );
  HS65_LH_AO22X9 U2534 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2479), .C(n2477), 
        .D(\registers[7][17] ), .Z(n1643) );
  HS65_LH_AO22X9 U2535 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2479), .C(n2477), 
        .D(\registers[7][18] ), .Z(n1644) );
  HS65_LH_AO22X9 U2536 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2479), .C(n2476), 
        .D(\registers[7][19] ), .Z(n1645) );
  HS65_LH_AO22X9 U2537 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2479), .C(n2476), 
        .D(\registers[7][20] ), .Z(n1646) );
  HS65_LH_AO22X9 U2538 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2479), .C(n2476), 
        .D(\registers[7][21] ), .Z(n1647) );
  HS65_LH_AO22X9 U2539 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2479), .C(n2476), 
        .D(\registers[7][22] ), .Z(n1648) );
  HS65_LH_AO22X9 U2540 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2479), .C(n2476), 
        .D(\registers[7][23] ), .Z(n1649) );
  HS65_LH_AO22X9 U2541 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2479), .C(n2476), 
        .D(\registers[7][24] ), .Z(n1650) );
  HS65_LH_AO22X9 U2542 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2479), .C(n2476), 
        .D(\registers[7][25] ), .Z(n1651) );
  HS65_LH_AO22X9 U2543 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2479), .C(n2476), 
        .D(\registers[7][26] ), .Z(n1652) );
  HS65_LH_AO22X9 U2544 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2479), .C(n2476), 
        .D(\registers[7][27] ), .Z(n1653) );
  HS65_LH_AO22X9 U2545 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2479), .C(n2476), 
        .D(\registers[7][28] ), .Z(n1654) );
  HS65_LH_AO22X9 U2546 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2479), .C(n2476), 
        .D(\registers[7][29] ), .Z(n1655) );
  HS65_LH_AO22X9 U2547 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2479), .C(n2476), 
        .D(\registers[7][30] ), .Z(n1656) );
  HS65_LH_AO22X9 U2548 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2478), .C(n2476), 
        .D(\registers[7][31] ), .Z(n1657) );
  HS65_LH_AO22X9 U2549 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n1422), .C(n1419), 
        .D(\registers[19][0] ), .Z(n2010) );
  HS65_LH_AO22X9 U2550 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n1422), .C(n1418), 
        .D(\registers[19][1] ), .Z(n2011) );
  HS65_LH_AO22X9 U2551 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n1422), .C(n1419), 
        .D(\registers[19][2] ), .Z(n2012) );
  HS65_LH_AO22X9 U2552 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n1422), .C(n1418), 
        .D(\registers[19][3] ), .Z(n2013) );
  HS65_LH_AO22X9 U2553 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n1422), .C(n1419), 
        .D(\registers[19][4] ), .Z(n2014) );
  HS65_LH_AO22X9 U2554 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n1422), .C(n1418), 
        .D(\registers[19][5] ), .Z(n2015) );
  HS65_LH_AO22X9 U2555 ( .A(n2709), .B(n1422), .C(n1419), .D(
        \registers[19][6] ), .Z(n2016) );
  HS65_LH_AO22X9 U2556 ( .A(n2711), .B(n1422), .C(n1419), .D(
        \registers[19][7] ), .Z(n2017) );
  HS65_LH_AO22X9 U2557 ( .A(n2713), .B(n1422), .C(n1419), .D(
        \registers[19][8] ), .Z(n2018) );
  HS65_LH_AO22X9 U2558 ( .A(n2715), .B(n1422), .C(n1419), .D(
        \registers[19][9] ), .Z(n2019) );
  HS65_LH_AO22X9 U2559 ( .A(n2717), .B(n1422), .C(n1419), .D(
        \registers[19][10] ), .Z(n2020) );
  HS65_LH_AO22X9 U2560 ( .A(n2719), .B(n1421), .C(n1419), .D(
        \registers[19][11] ), .Z(n2021) );
  HS65_LH_AO22X9 U2561 ( .A(n2721), .B(n1421), .C(n1419), .D(
        \registers[19][12] ), .Z(n2022) );
  HS65_LH_AO22X9 U2562 ( .A(n2723), .B(n1421), .C(n1419), .D(
        \registers[19][13] ), .Z(n2023) );
  HS65_LH_AO22X9 U2563 ( .A(n2725), .B(n1421), .C(n1419), .D(
        \registers[19][14] ), .Z(n2024) );
  HS65_LH_AO22X9 U2564 ( .A(n2727), .B(n1421), .C(n1419), .D(
        \registers[19][15] ), .Z(n2025) );
  HS65_LH_AO22X9 U2565 ( .A(n2729), .B(n1421), .C(n1419), .D(
        \registers[19][16] ), .Z(n2026) );
  HS65_LH_AO22X9 U2566 ( .A(n2731), .B(n1421), .C(n1419), .D(
        \registers[19][17] ), .Z(n2027) );
  HS65_LH_AO22X9 U2567 ( .A(n2733), .B(n1421), .C(n1419), .D(
        \registers[19][18] ), .Z(n2028) );
  HS65_LH_AO22X9 U2568 ( .A(n2735), .B(n1421), .C(n1418), .D(
        \registers[19][19] ), .Z(n2029) );
  HS65_LH_AO22X9 U2569 ( .A(n2737), .B(n1421), .C(n1418), .D(
        \registers[19][20] ), .Z(n2030) );
  HS65_LH_AO22X9 U2570 ( .A(n2739), .B(n1421), .C(n1418), .D(
        \registers[19][21] ), .Z(n2031) );
  HS65_LH_AO22X9 U2571 ( .A(n2741), .B(n1421), .C(n1418), .D(
        \registers[19][22] ), .Z(n2032) );
  HS65_LH_AO22X9 U2572 ( .A(n2743), .B(n1421), .C(n1418), .D(
        \registers[19][23] ), .Z(n2033) );
  HS65_LH_AO22X9 U2573 ( .A(n2745), .B(n1421), .C(n1418), .D(
        \registers[19][24] ), .Z(n2034) );
  HS65_LH_AO22X9 U2574 ( .A(n2747), .B(n1421), .C(n1418), .D(
        \registers[19][25] ), .Z(n2035) );
  HS65_LH_AO22X9 U2575 ( .A(n2749), .B(n1421), .C(n1418), .D(
        \registers[19][26] ), .Z(n2036) );
  HS65_LH_AO22X9 U2576 ( .A(n2751), .B(n1421), .C(n1418), .D(
        \registers[19][27] ), .Z(n2037) );
  HS65_LH_AO22X9 U2577 ( .A(n2753), .B(n1421), .C(n1418), .D(
        \registers[19][28] ), .Z(n2038) );
  HS65_LH_AO22X9 U2578 ( .A(n2755), .B(n1421), .C(n1418), .D(
        \registers[19][29] ), .Z(n2039) );
  HS65_LH_AO22X9 U2579 ( .A(n2757), .B(n1421), .C(n1418), .D(
        \registers[19][30] ), .Z(n2040) );
  HS65_LH_AO22X9 U2580 ( .A(n2759), .B(n1420), .C(n1418), .D(
        \registers[19][31] ), .Z(n2041) );
  HS65_LH_AO22X9 U2581 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n332), .C(n329), 
        .D(\registers[23][0] ), .Z(n2138) );
  HS65_LH_AO22X9 U2582 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n332), .C(n328), 
        .D(\registers[23][1] ), .Z(n2139) );
  HS65_LH_AO22X9 U2583 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n332), .C(n329), 
        .D(\registers[23][2] ), .Z(n2140) );
  HS65_LH_AO22X9 U2584 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n332), .C(n328), 
        .D(\registers[23][3] ), .Z(n2141) );
  HS65_LH_AO22X9 U2585 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n332), .C(n329), 
        .D(\registers[23][4] ), .Z(n2142) );
  HS65_LH_AO22X9 U2586 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n332), .C(n328), 
        .D(\registers[23][5] ), .Z(n2143) );
  HS65_LH_AO22X9 U2587 ( .A(n2709), .B(n332), .C(n329), .D(\registers[23][6] ), 
        .Z(n2144) );
  HS65_LH_AO22X9 U2588 ( .A(n2711), .B(n332), .C(n329), .D(\registers[23][7] ), 
        .Z(n2145) );
  HS65_LH_AO22X9 U2589 ( .A(n2713), .B(n332), .C(n329), .D(\registers[23][8] ), 
        .Z(n2146) );
  HS65_LH_AO22X9 U2590 ( .A(n2715), .B(n332), .C(n329), .D(\registers[23][9] ), 
        .Z(n2147) );
  HS65_LH_AO22X9 U2591 ( .A(n2717), .B(n332), .C(n329), .D(\registers[23][10] ), .Z(n2148) );
  HS65_LH_AO22X9 U2592 ( .A(n2719), .B(n331), .C(n329), .D(\registers[23][11] ), .Z(n2149) );
  HS65_LH_AO22X9 U2593 ( .A(n2721), .B(n331), .C(n329), .D(\registers[23][12] ), .Z(n2150) );
  HS65_LH_AO22X9 U2594 ( .A(n2723), .B(n331), .C(n329), .D(\registers[23][13] ), .Z(n2151) );
  HS65_LH_AO22X9 U2595 ( .A(n2725), .B(n331), .C(n329), .D(\registers[23][14] ), .Z(n2152) );
  HS65_LH_AO22X9 U2596 ( .A(n2727), .B(n331), .C(n329), .D(\registers[23][15] ), .Z(n2153) );
  HS65_LH_AO22X9 U2597 ( .A(n2729), .B(n331), .C(n329), .D(\registers[23][16] ), .Z(n2154) );
  HS65_LH_AO22X9 U2598 ( .A(n2731), .B(n331), .C(n329), .D(\registers[23][17] ), .Z(n2155) );
  HS65_LH_AO22X9 U2599 ( .A(n2733), .B(n331), .C(n329), .D(\registers[23][18] ), .Z(n2156) );
  HS65_LH_AO22X9 U2600 ( .A(n2735), .B(n331), .C(n328), .D(\registers[23][19] ), .Z(n2157) );
  HS65_LH_AO22X9 U2601 ( .A(n2737), .B(n331), .C(n328), .D(\registers[23][20] ), .Z(n2158) );
  HS65_LH_AO22X9 U2602 ( .A(n2739), .B(n331), .C(n328), .D(\registers[23][21] ), .Z(n2159) );
  HS65_LH_AO22X9 U2603 ( .A(n2741), .B(n331), .C(n328), .D(\registers[23][22] ), .Z(n2160) );
  HS65_LH_AO22X9 U2604 ( .A(n2743), .B(n331), .C(n328), .D(\registers[23][23] ), .Z(n2161) );
  HS65_LH_AO22X9 U2605 ( .A(n2745), .B(n331), .C(n328), .D(\registers[23][24] ), .Z(n2162) );
  HS65_LH_AO22X9 U2606 ( .A(n2747), .B(n331), .C(n328), .D(\registers[23][25] ), .Z(n2163) );
  HS65_LH_AO22X9 U2607 ( .A(n2749), .B(n331), .C(n328), .D(\registers[23][26] ), .Z(n2164) );
  HS65_LH_AO22X9 U2608 ( .A(n2751), .B(n331), .C(n328), .D(\registers[23][27] ), .Z(n2165) );
  HS65_LH_AO22X9 U2609 ( .A(n2753), .B(n331), .C(n328), .D(\registers[23][28] ), .Z(n2166) );
  HS65_LH_AO22X9 U2610 ( .A(n2755), .B(n331), .C(n328), .D(\registers[23][29] ), .Z(n2167) );
  HS65_LH_AO22X9 U2611 ( .A(n2757), .B(n331), .C(n328), .D(\registers[23][30] ), .Z(n2168) );
  HS65_LH_AO22X9 U2612 ( .A(n2759), .B(n330), .C(n328), .D(\registers[23][31] ), .Z(n2169) );
  HS65_LH_AO22X9 U2613 ( .A(n2697), .B(n2490), .C(n2487), .D(\registers[5][0] ), .Z(n1562) );
  HS65_LH_AO22X9 U2614 ( .A(n2699), .B(n2490), .C(n2486), .D(\registers[5][1] ), .Z(n1563) );
  HS65_LH_AO22X9 U2615 ( .A(n2701), .B(n2490), .C(n2487), .D(\registers[5][2] ), .Z(n1564) );
  HS65_LH_AO22X9 U2616 ( .A(n2703), .B(n2490), .C(n2486), .D(\registers[5][3] ), .Z(n1565) );
  HS65_LH_AO22X9 U2617 ( .A(n2705), .B(n2490), .C(n2487), .D(\registers[5][4] ), .Z(n1566) );
  HS65_LH_AO22X9 U2618 ( .A(n2707), .B(n2490), .C(n2486), .D(\registers[5][5] ), .Z(n1567) );
  HS65_LH_AO22X9 U2619 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2490), .C(n2487), 
        .D(\registers[5][6] ), .Z(n1568) );
  HS65_LH_AO22X9 U2620 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2490), .C(n2487), 
        .D(\registers[5][7] ), .Z(n1569) );
  HS65_LH_AO22X9 U2621 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2490), .C(n2487), 
        .D(\registers[5][8] ), .Z(n1570) );
  HS65_LH_AO22X9 U2622 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2490), .C(n2487), 
        .D(\registers[5][9] ), .Z(n1571) );
  HS65_LH_AO22X9 U2623 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2490), .C(n2487), 
        .D(\registers[5][10] ), .Z(n1572) );
  HS65_LH_AO22X9 U2624 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2489), .C(n2487), 
        .D(\registers[5][11] ), .Z(n1573) );
  HS65_LH_AO22X9 U2625 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2489), .C(n2487), 
        .D(\registers[5][12] ), .Z(n1574) );
  HS65_LH_AO22X9 U2626 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2489), .C(n2487), 
        .D(\registers[5][13] ), .Z(n1575) );
  HS65_LH_AO22X9 U2627 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2489), .C(n2487), 
        .D(\registers[5][14] ), .Z(n1576) );
  HS65_LH_AO22X9 U2628 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2489), .C(n2487), 
        .D(\registers[5][15] ), .Z(n1577) );
  HS65_LH_AO22X9 U2629 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2489), .C(n2487), 
        .D(\registers[5][16] ), .Z(n1578) );
  HS65_LH_AO22X9 U2630 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2489), .C(n2487), 
        .D(\registers[5][17] ), .Z(n1579) );
  HS65_LH_AO22X9 U2631 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2489), .C(n2487), 
        .D(\registers[5][18] ), .Z(n1580) );
  HS65_LH_AO22X9 U2632 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2489), .C(n2486), 
        .D(\registers[5][19] ), .Z(n1581) );
  HS65_LH_AO22X9 U2633 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2489), .C(n2486), 
        .D(\registers[5][20] ), .Z(n1582) );
  HS65_LH_AO22X9 U2634 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2489), .C(n2486), 
        .D(\registers[5][21] ), .Z(n1583) );
  HS65_LH_AO22X9 U2635 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2489), .C(n2486), 
        .D(\registers[5][22] ), .Z(n1584) );
  HS65_LH_AO22X9 U2636 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2489), .C(n2486), 
        .D(\registers[5][23] ), .Z(n1585) );
  HS65_LH_AO22X9 U2637 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2489), .C(n2486), 
        .D(\registers[5][24] ), .Z(n1586) );
  HS65_LH_AO22X9 U2638 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2489), .C(n2486), 
        .D(\registers[5][25] ), .Z(n1587) );
  HS65_LH_AO22X9 U2639 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2489), .C(n2486), 
        .D(\registers[5][26] ), .Z(n1588) );
  HS65_LH_AO22X9 U2640 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2489), .C(n2486), 
        .D(\registers[5][27] ), .Z(n1589) );
  HS65_LH_AO22X9 U2641 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2489), .C(n2486), 
        .D(\registers[5][28] ), .Z(n1590) );
  HS65_LH_AO22X9 U2642 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2489), .C(n2486), 
        .D(\registers[5][29] ), .Z(n1591) );
  HS65_LH_AO22X9 U2643 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2489), .C(n2486), 
        .D(\registers[5][30] ), .Z(n1592) );
  HS65_LH_AO22X9 U2644 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2488), .C(n2486), 
        .D(\registers[5][31] ), .Z(n1593) );
  HS65_LH_AO22X9 U2645 ( .A(n2697), .B(n2485), .C(n2482), .D(\registers[6][0] ), .Z(n1594) );
  HS65_LH_AO22X9 U2646 ( .A(n2699), .B(n2485), .C(n2481), .D(\registers[6][1] ), .Z(n1595) );
  HS65_LH_AO22X9 U2647 ( .A(n2701), .B(n2485), .C(n2482), .D(\registers[6][2] ), .Z(n1596) );
  HS65_LH_AO22X9 U2648 ( .A(n2703), .B(n2485), .C(n2481), .D(\registers[6][3] ), .Z(n1597) );
  HS65_LH_AO22X9 U2649 ( .A(n2705), .B(n2485), .C(n2482), .D(\registers[6][4] ), .Z(n1598) );
  HS65_LH_AO22X9 U2650 ( .A(n2707), .B(n2485), .C(n2481), .D(\registers[6][5] ), .Z(n1599) );
  HS65_LH_AO22X9 U2651 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2485), .C(n2482), 
        .D(\registers[6][6] ), .Z(n1600) );
  HS65_LH_AO22X9 U2652 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2485), .C(n2482), 
        .D(\registers[6][7] ), .Z(n1601) );
  HS65_LH_AO22X9 U2653 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2485), .C(n2482), 
        .D(\registers[6][8] ), .Z(n1602) );
  HS65_LH_AO22X9 U2654 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2485), .C(n2482), 
        .D(\registers[6][9] ), .Z(n1603) );
  HS65_LH_AO22X9 U2655 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2485), .C(n2482), 
        .D(\registers[6][10] ), .Z(n1604) );
  HS65_LH_AO22X9 U2656 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2484), .C(n2482), 
        .D(\registers[6][11] ), .Z(n1605) );
  HS65_LH_AO22X9 U2657 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2484), .C(n2482), 
        .D(\registers[6][12] ), .Z(n1606) );
  HS65_LH_AO22X9 U2658 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2484), .C(n2482), 
        .D(\registers[6][13] ), .Z(n1607) );
  HS65_LH_AO22X9 U2659 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2484), .C(n2482), 
        .D(\registers[6][14] ), .Z(n1608) );
  HS65_LH_AO22X9 U2660 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2484), .C(n2482), 
        .D(\registers[6][15] ), .Z(n1609) );
  HS65_LH_AO22X9 U2661 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2484), .C(n2482), 
        .D(\registers[6][16] ), .Z(n1610) );
  HS65_LH_AO22X9 U2662 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2484), .C(n2482), 
        .D(\registers[6][17] ), .Z(n1611) );
  HS65_LH_AO22X9 U2663 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2484), .C(n2482), 
        .D(\registers[6][18] ), .Z(n1612) );
  HS65_LH_AO22X9 U2664 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2484), .C(n2481), 
        .D(\registers[6][19] ), .Z(n1613) );
  HS65_LH_AO22X9 U2665 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2484), .C(n2481), 
        .D(\registers[6][20] ), .Z(n1614) );
  HS65_LH_AO22X9 U2666 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2484), .C(n2481), 
        .D(\registers[6][21] ), .Z(n1615) );
  HS65_LH_AO22X9 U2667 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2484), .C(n2481), 
        .D(\registers[6][22] ), .Z(n1616) );
  HS65_LH_AO22X9 U2668 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2484), .C(n2481), 
        .D(\registers[6][23] ), .Z(n1617) );
  HS65_LH_AO22X9 U2669 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2484), .C(n2481), 
        .D(\registers[6][24] ), .Z(n1618) );
  HS65_LH_AO22X9 U2670 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2484), .C(n2481), 
        .D(\registers[6][25] ), .Z(n1619) );
  HS65_LH_AO22X9 U2671 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2484), .C(n2481), 
        .D(\registers[6][26] ), .Z(n1620) );
  HS65_LH_AO22X9 U2672 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2484), .C(n2481), 
        .D(\registers[6][27] ), .Z(n1621) );
  HS65_LH_AO22X9 U2673 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2484), .C(n2481), 
        .D(\registers[6][28] ), .Z(n1622) );
  HS65_LH_AO22X9 U2674 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2484), .C(n2481), 
        .D(\registers[6][29] ), .Z(n1623) );
  HS65_LH_AO22X9 U2675 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2484), .C(n2481), 
        .D(\registers[6][30] ), .Z(n1624) );
  HS65_LH_AO22X9 U2676 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2483), .C(n2481), 
        .D(\registers[6][31] ), .Z(n1625) );
  HS65_LH_AO22X9 U2677 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n2430), .C(n2427), 
        .D(\registers[17][0] ), .Z(n1946) );
  HS65_LH_AO22X9 U2678 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n2430), .C(n2426), 
        .D(\registers[17][1] ), .Z(n1947) );
  HS65_LH_AO22X9 U2679 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n2430), .C(n2427), 
        .D(\registers[17][2] ), .Z(n1948) );
  HS65_LH_AO22X9 U2680 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n2430), .C(n2426), 
        .D(\registers[17][3] ), .Z(n1949) );
  HS65_LH_AO22X9 U2681 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n2430), .C(n2427), 
        .D(\registers[17][4] ), .Z(n1950) );
  HS65_LH_AO22X9 U2682 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n2430), .C(n2426), 
        .D(\registers[17][5] ), .Z(n1951) );
  HS65_LH_AO22X9 U2683 ( .A(n2709), .B(n2430), .C(n2427), .D(
        \registers[17][6] ), .Z(n1952) );
  HS65_LH_AO22X9 U2684 ( .A(n2711), .B(n2430), .C(n2427), .D(
        \registers[17][7] ), .Z(n1953) );
  HS65_LH_AO22X9 U2685 ( .A(n2713), .B(n2430), .C(n2427), .D(
        \registers[17][8] ), .Z(n1954) );
  HS65_LH_AO22X9 U2686 ( .A(n2715), .B(n2430), .C(n2427), .D(
        \registers[17][9] ), .Z(n1955) );
  HS65_LH_AO22X9 U2687 ( .A(n2717), .B(n2430), .C(n2427), .D(
        \registers[17][10] ), .Z(n1956) );
  HS65_LH_AO22X9 U2688 ( .A(n2719), .B(n2429), .C(n2427), .D(
        \registers[17][11] ), .Z(n1957) );
  HS65_LH_AO22X9 U2689 ( .A(n2721), .B(n2429), .C(n2427), .D(
        \registers[17][12] ), .Z(n1958) );
  HS65_LH_AO22X9 U2690 ( .A(n2723), .B(n2429), .C(n2427), .D(
        \registers[17][13] ), .Z(n1959) );
  HS65_LH_AO22X9 U2691 ( .A(n2725), .B(n2429), .C(n2427), .D(
        \registers[17][14] ), .Z(n1960) );
  HS65_LH_AO22X9 U2692 ( .A(n2727), .B(n2429), .C(n2427), .D(
        \registers[17][15] ), .Z(n1961) );
  HS65_LH_AO22X9 U2693 ( .A(n2729), .B(n2429), .C(n2427), .D(
        \registers[17][16] ), .Z(n1962) );
  HS65_LH_AO22X9 U2694 ( .A(n2731), .B(n2429), .C(n2427), .D(
        \registers[17][17] ), .Z(n1963) );
  HS65_LH_AO22X9 U2695 ( .A(n2733), .B(n2429), .C(n2427), .D(
        \registers[17][18] ), .Z(n1964) );
  HS65_LH_AO22X9 U2696 ( .A(n2735), .B(n2429), .C(n2426), .D(
        \registers[17][19] ), .Z(n1965) );
  HS65_LH_AO22X9 U2697 ( .A(n2737), .B(n2429), .C(n2426), .D(
        \registers[17][20] ), .Z(n1966) );
  HS65_LH_AO22X9 U2698 ( .A(n2739), .B(n2429), .C(n2426), .D(
        \registers[17][21] ), .Z(n1967) );
  HS65_LH_AO22X9 U2699 ( .A(n2741), .B(n2429), .C(n2426), .D(
        \registers[17][22] ), .Z(n1968) );
  HS65_LH_AO22X9 U2700 ( .A(n2743), .B(n2429), .C(n2426), .D(
        \registers[17][23] ), .Z(n1969) );
  HS65_LH_AO22X9 U2701 ( .A(n2745), .B(n2429), .C(n2426), .D(
        \registers[17][24] ), .Z(n1970) );
  HS65_LH_AO22X9 U2702 ( .A(n2747), .B(n2429), .C(n2426), .D(
        \registers[17][25] ), .Z(n1971) );
  HS65_LH_AO22X9 U2703 ( .A(n2749), .B(n2429), .C(n2426), .D(
        \registers[17][26] ), .Z(n1972) );
  HS65_LH_AO22X9 U2704 ( .A(n2751), .B(n2429), .C(n2426), .D(
        \registers[17][27] ), .Z(n1973) );
  HS65_LH_AO22X9 U2705 ( .A(n2753), .B(n2429), .C(n2426), .D(
        \registers[17][28] ), .Z(n1974) );
  HS65_LH_AO22X9 U2706 ( .A(n2755), .B(n2429), .C(n2426), .D(
        \registers[17][29] ), .Z(n1975) );
  HS65_LH_AO22X9 U2707 ( .A(n2757), .B(n2429), .C(n2426), .D(
        \registers[17][30] ), .Z(n1976) );
  HS65_LH_AO22X9 U2708 ( .A(n2759), .B(n2428), .C(n2426), .D(
        \registers[17][31] ), .Z(n1977) );
  HS65_LH_AO22X9 U2709 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n1433), .C(n1424), 
        .D(\registers[18][0] ), .Z(n1978) );
  HS65_LH_AO22X9 U2710 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n1433), .C(n1423), 
        .D(\registers[18][1] ), .Z(n1979) );
  HS65_LH_AO22X9 U2711 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n1433), .C(n1424), 
        .D(\registers[18][2] ), .Z(n1980) );
  HS65_LH_AO22X9 U2712 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n1433), .C(n1423), 
        .D(\registers[18][3] ), .Z(n1981) );
  HS65_LH_AO22X9 U2713 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n1433), .C(n1424), 
        .D(\registers[18][4] ), .Z(n1982) );
  HS65_LH_AO22X9 U2714 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n1433), .C(n1423), 
        .D(\registers[18][5] ), .Z(n1983) );
  HS65_LH_AO22X9 U2715 ( .A(n2709), .B(n1433), .C(n1424), .D(
        \registers[18][6] ), .Z(n1984) );
  HS65_LH_AO22X9 U2716 ( .A(n2711), .B(n1433), .C(n1424), .D(
        \registers[18][7] ), .Z(n1985) );
  HS65_LH_AO22X9 U2717 ( .A(n2713), .B(n1433), .C(n1424), .D(
        \registers[18][8] ), .Z(n1986) );
  HS65_LH_AO22X9 U2718 ( .A(n2715), .B(n1433), .C(n1424), .D(
        \registers[18][9] ), .Z(n1987) );
  HS65_LH_AO22X9 U2719 ( .A(n2717), .B(n1433), .C(n1424), .D(
        \registers[18][10] ), .Z(n1988) );
  HS65_LH_AO22X9 U2720 ( .A(n2719), .B(n1432), .C(n1424), .D(
        \registers[18][11] ), .Z(n1989) );
  HS65_LH_AO22X9 U2721 ( .A(n2721), .B(n1432), .C(n1424), .D(
        \registers[18][12] ), .Z(n1990) );
  HS65_LH_AO22X9 U2722 ( .A(n2723), .B(n1432), .C(n1424), .D(
        \registers[18][13] ), .Z(n1991) );
  HS65_LH_AO22X9 U2723 ( .A(n2725), .B(n1432), .C(n1424), .D(
        \registers[18][14] ), .Z(n1992) );
  HS65_LH_AO22X9 U2724 ( .A(n2727), .B(n1432), .C(n1424), .D(
        \registers[18][15] ), .Z(n1993) );
  HS65_LH_AO22X9 U2725 ( .A(n2729), .B(n1432), .C(n1424), .D(
        \registers[18][16] ), .Z(n1994) );
  HS65_LH_AO22X9 U2726 ( .A(n2731), .B(n1432), .C(n1424), .D(
        \registers[18][17] ), .Z(n1995) );
  HS65_LH_AO22X9 U2727 ( .A(n2733), .B(n1432), .C(n1424), .D(
        \registers[18][18] ), .Z(n1996) );
  HS65_LH_AO22X9 U2728 ( .A(n2735), .B(n1432), .C(n1423), .D(
        \registers[18][19] ), .Z(n1997) );
  HS65_LH_AO22X9 U2729 ( .A(n2737), .B(n1432), .C(n1423), .D(
        \registers[18][20] ), .Z(n1998) );
  HS65_LH_AO22X9 U2730 ( .A(n2739), .B(n1432), .C(n1423), .D(
        \registers[18][21] ), .Z(n1999) );
  HS65_LH_AO22X9 U2731 ( .A(n2741), .B(n1432), .C(n1423), .D(
        \registers[18][22] ), .Z(n2000) );
  HS65_LH_AO22X9 U2732 ( .A(n2743), .B(n1432), .C(n1423), .D(
        \registers[18][23] ), .Z(n2001) );
  HS65_LH_AO22X9 U2733 ( .A(n2745), .B(n1432), .C(n1423), .D(
        \registers[18][24] ), .Z(n2002) );
  HS65_LH_AO22X9 U2734 ( .A(n2747), .B(n1432), .C(n1423), .D(
        \registers[18][25] ), .Z(n2003) );
  HS65_LH_AO22X9 U2735 ( .A(n2749), .B(n1432), .C(n1423), .D(
        \registers[18][26] ), .Z(n2004) );
  HS65_LH_AO22X9 U2736 ( .A(n2751), .B(n1432), .C(n1423), .D(
        \registers[18][27] ), .Z(n2005) );
  HS65_LH_AO22X9 U2737 ( .A(n2753), .B(n1432), .C(n1423), .D(
        \registers[18][28] ), .Z(n2006) );
  HS65_LH_AO22X9 U2738 ( .A(n2755), .B(n1432), .C(n1423), .D(
        \registers[18][29] ), .Z(n2007) );
  HS65_LH_AO22X9 U2739 ( .A(n2757), .B(n1432), .C(n1423), .D(
        \registers[18][30] ), .Z(n2008) );
  HS65_LH_AO22X9 U2740 ( .A(n2759), .B(n1427), .C(n1423), .D(
        \registers[18][31] ), .Z(n2009) );
  HS65_LH_AO22X9 U2741 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n1403), .C(n1397), 
        .D(\registers[21][0] ), .Z(n2074) );
  HS65_LH_AO22X9 U2742 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n1403), .C(n1395), 
        .D(\registers[21][1] ), .Z(n2075) );
  HS65_LH_AO22X9 U2743 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n1403), .C(n1397), 
        .D(\registers[21][2] ), .Z(n2076) );
  HS65_LH_AO22X9 U2744 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n1403), .C(n1395), 
        .D(\registers[21][3] ), .Z(n2077) );
  HS65_LH_AO22X9 U2745 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n1403), .C(n1397), 
        .D(\registers[21][4] ), .Z(n2078) );
  HS65_LH_AO22X9 U2746 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n1403), .C(n1395), 
        .D(\registers[21][5] ), .Z(n2079) );
  HS65_LH_AO22X9 U2747 ( .A(n2709), .B(n1403), .C(n1397), .D(
        \registers[21][6] ), .Z(n2080) );
  HS65_LH_AO22X9 U2748 ( .A(n2711), .B(n1403), .C(n1397), .D(
        \registers[21][7] ), .Z(n2081) );
  HS65_LH_AO22X9 U2749 ( .A(n2713), .B(n1403), .C(n1397), .D(
        \registers[21][8] ), .Z(n2082) );
  HS65_LH_AO22X9 U2750 ( .A(n2715), .B(n1403), .C(n1397), .D(
        \registers[21][9] ), .Z(n2083) );
  HS65_LH_AO22X9 U2751 ( .A(n2717), .B(n1403), .C(n1397), .D(
        \registers[21][10] ), .Z(n2084) );
  HS65_LH_AO22X9 U2752 ( .A(n2719), .B(n1401), .C(n1397), .D(
        \registers[21][11] ), .Z(n2085) );
  HS65_LH_AO22X9 U2753 ( .A(n2721), .B(n1401), .C(n1397), .D(
        \registers[21][12] ), .Z(n2086) );
  HS65_LH_AO22X9 U2754 ( .A(n2723), .B(n1401), .C(n1397), .D(
        \registers[21][13] ), .Z(n2087) );
  HS65_LH_AO22X9 U2755 ( .A(n2725), .B(n1401), .C(n1397), .D(
        \registers[21][14] ), .Z(n2088) );
  HS65_LH_AO22X9 U2756 ( .A(n2727), .B(n1401), .C(n1397), .D(
        \registers[21][15] ), .Z(n2089) );
  HS65_LH_AO22X9 U2757 ( .A(n2729), .B(n1401), .C(n1397), .D(
        \registers[21][16] ), .Z(n2090) );
  HS65_LH_AO22X9 U2758 ( .A(n2731), .B(n1401), .C(n1397), .D(
        \registers[21][17] ), .Z(n2091) );
  HS65_LH_AO22X9 U2759 ( .A(n2733), .B(n1401), .C(n1397), .D(
        \registers[21][18] ), .Z(n2092) );
  HS65_LH_AO22X9 U2760 ( .A(n2735), .B(n1401), .C(n1395), .D(
        \registers[21][19] ), .Z(n2093) );
  HS65_LH_AO22X9 U2761 ( .A(n2737), .B(n1401), .C(n1395), .D(
        \registers[21][20] ), .Z(n2094) );
  HS65_LH_AO22X9 U2762 ( .A(n2739), .B(n1401), .C(n1395), .D(
        \registers[21][21] ), .Z(n2095) );
  HS65_LH_AO22X9 U2763 ( .A(n2741), .B(n1401), .C(n1395), .D(
        \registers[21][22] ), .Z(n2096) );
  HS65_LH_AO22X9 U2764 ( .A(n2743), .B(n1401), .C(n1395), .D(
        \registers[21][23] ), .Z(n2097) );
  HS65_LH_AO22X9 U2765 ( .A(n2745), .B(n1401), .C(n1395), .D(
        \registers[21][24] ), .Z(n2098) );
  HS65_LH_AO22X9 U2766 ( .A(n2747), .B(n1401), .C(n1395), .D(
        \registers[21][25] ), .Z(n2099) );
  HS65_LH_AO22X9 U2767 ( .A(n2749), .B(n1401), .C(n1395), .D(
        \registers[21][26] ), .Z(n2100) );
  HS65_LH_AO22X9 U2768 ( .A(n2751), .B(n1401), .C(n1395), .D(
        \registers[21][27] ), .Z(n2101) );
  HS65_LH_AO22X9 U2769 ( .A(n2753), .B(n1401), .C(n1395), .D(
        \registers[21][28] ), .Z(n2102) );
  HS65_LH_AO22X9 U2770 ( .A(n2755), .B(n1401), .C(n1395), .D(
        \registers[21][29] ), .Z(n2103) );
  HS65_LH_AO22X9 U2771 ( .A(n2757), .B(n1401), .C(n1395), .D(
        \registers[21][30] ), .Z(n2104) );
  HS65_LH_AO22X9 U2772 ( .A(n2759), .B(n1399), .C(n1395), .D(
        \registers[21][31] ), .Z(n2105) );
  HS65_LH_AO22X9 U2773 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n1392), .C(n334), 
        .D(\registers[22][0] ), .Z(n2106) );
  HS65_LH_AO22X9 U2774 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n1392), .C(n333), 
        .D(\registers[22][1] ), .Z(n2107) );
  HS65_LH_AO22X9 U2775 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n1392), .C(n334), 
        .D(\registers[22][2] ), .Z(n2108) );
  HS65_LH_AO22X9 U2776 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n1392), .C(n333), 
        .D(\registers[22][3] ), .Z(n2109) );
  HS65_LH_AO22X9 U2777 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n1392), .C(n334), 
        .D(\registers[22][4] ), .Z(n2110) );
  HS65_LH_AO22X9 U2778 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n1392), .C(n333), 
        .D(\registers[22][5] ), .Z(n2111) );
  HS65_LH_AO22X9 U2779 ( .A(n2709), .B(n1392), .C(n334), .D(\registers[22][6] ), .Z(n2112) );
  HS65_LH_AO22X9 U2780 ( .A(n2711), .B(n1392), .C(n334), .D(\registers[22][7] ), .Z(n2113) );
  HS65_LH_AO22X9 U2781 ( .A(n2713), .B(n1392), .C(n334), .D(\registers[22][8] ), .Z(n2114) );
  HS65_LH_AO22X9 U2782 ( .A(n2715), .B(n1392), .C(n334), .D(\registers[22][9] ), .Z(n2115) );
  HS65_LH_AO22X9 U2783 ( .A(n2717), .B(n1392), .C(n334), .D(
        \registers[22][10] ), .Z(n2116) );
  HS65_LH_AO22X9 U2784 ( .A(n2719), .B(n880), .C(n334), .D(\registers[22][11] ), .Z(n2117) );
  HS65_LH_AO22X9 U2785 ( .A(n2721), .B(n880), .C(n334), .D(\registers[22][12] ), .Z(n2118) );
  HS65_LH_AO22X9 U2786 ( .A(n2723), .B(n880), .C(n334), .D(\registers[22][13] ), .Z(n2119) );
  HS65_LH_AO22X9 U2787 ( .A(n2725), .B(n880), .C(n334), .D(\registers[22][14] ), .Z(n2120) );
  HS65_LH_AO22X9 U2788 ( .A(n2727), .B(n880), .C(n334), .D(\registers[22][15] ), .Z(n2121) );
  HS65_LH_AO22X9 U2789 ( .A(n2729), .B(n880), .C(n334), .D(\registers[22][16] ), .Z(n2122) );
  HS65_LH_AO22X9 U2790 ( .A(n2731), .B(n880), .C(n334), .D(\registers[22][17] ), .Z(n2123) );
  HS65_LH_AO22X9 U2791 ( .A(n2733), .B(n880), .C(n334), .D(\registers[22][18] ), .Z(n2124) );
  HS65_LH_AO22X9 U2792 ( .A(n2735), .B(n880), .C(n333), .D(\registers[22][19] ), .Z(n2125) );
  HS65_LH_AO22X9 U2793 ( .A(n2737), .B(n880), .C(n333), .D(\registers[22][20] ), .Z(n2126) );
  HS65_LH_AO22X9 U2794 ( .A(n2739), .B(n880), .C(n333), .D(\registers[22][21] ), .Z(n2127) );
  HS65_LH_AO22X9 U2795 ( .A(n2741), .B(n880), .C(n333), .D(\registers[22][22] ), .Z(n2128) );
  HS65_LH_AO22X9 U2796 ( .A(n2743), .B(n880), .C(n333), .D(\registers[22][23] ), .Z(n2129) );
  HS65_LH_AO22X9 U2797 ( .A(n2745), .B(n880), .C(n333), .D(\registers[22][24] ), .Z(n2130) );
  HS65_LH_AO22X9 U2798 ( .A(n2747), .B(n880), .C(n333), .D(\registers[22][25] ), .Z(n2131) );
  HS65_LH_AO22X9 U2799 ( .A(n2749), .B(n880), .C(n333), .D(\registers[22][26] ), .Z(n2132) );
  HS65_LH_AO22X9 U2800 ( .A(n2751), .B(n880), .C(n333), .D(\registers[22][27] ), .Z(n2133) );
  HS65_LH_AO22X9 U2801 ( .A(n2753), .B(n880), .C(n333), .D(\registers[22][28] ), .Z(n2134) );
  HS65_LH_AO22X9 U2802 ( .A(n2755), .B(n880), .C(n333), .D(\registers[22][29] ), .Z(n2135) );
  HS65_LH_AO22X9 U2803 ( .A(n2757), .B(n880), .C(n333), .D(\registers[22][30] ), .Z(n2136) );
  HS65_LH_AO22X9 U2804 ( .A(n2759), .B(n352), .C(n333), .D(\registers[22][31] ), .Z(n2137) );
  HS65_LH_AO22X9 U2805 ( .A(n2697), .B(n2495), .C(n2492), .D(\registers[4][0] ), .Z(n1530) );
  HS65_LH_AO22X9 U2806 ( .A(n2699), .B(n2495), .C(n2491), .D(\registers[4][1] ), .Z(n1531) );
  HS65_LH_AO22X9 U2807 ( .A(n2701), .B(n2495), .C(n2492), .D(\registers[4][2] ), .Z(n1532) );
  HS65_LH_AO22X9 U2808 ( .A(n2703), .B(n2495), .C(n2491), .D(\registers[4][3] ), .Z(n1533) );
  HS65_LH_AO22X9 U2809 ( .A(n2705), .B(n2495), .C(n2492), .D(\registers[4][4] ), .Z(n1534) );
  HS65_LH_AO22X9 U2810 ( .A(n2707), .B(n2495), .C(n2491), .D(\registers[4][5] ), .Z(n1535) );
  HS65_LH_AO22X9 U2811 ( .A(\regfile_i[WRITE_DATA][6] ), .B(n2495), .C(n2492), 
        .D(\registers[4][6] ), .Z(n1536) );
  HS65_LH_AO22X9 U2812 ( .A(\regfile_i[WRITE_DATA][7] ), .B(n2495), .C(n2492), 
        .D(\registers[4][7] ), .Z(n1537) );
  HS65_LH_AO22X9 U2813 ( .A(\regfile_i[WRITE_DATA][8] ), .B(n2495), .C(n2492), 
        .D(\registers[4][8] ), .Z(n1538) );
  HS65_LH_AO22X9 U2814 ( .A(\regfile_i[WRITE_DATA][9] ), .B(n2495), .C(n2492), 
        .D(\registers[4][9] ), .Z(n1539) );
  HS65_LH_AO22X9 U2815 ( .A(\regfile_i[WRITE_DATA][10] ), .B(n2495), .C(n2492), 
        .D(\registers[4][10] ), .Z(n1540) );
  HS65_LH_AO22X9 U2816 ( .A(\regfile_i[WRITE_DATA][11] ), .B(n2494), .C(n2492), 
        .D(\registers[4][11] ), .Z(n1541) );
  HS65_LH_AO22X9 U2817 ( .A(\regfile_i[WRITE_DATA][12] ), .B(n2494), .C(n2492), 
        .D(\registers[4][12] ), .Z(n1542) );
  HS65_LH_AO22X9 U2818 ( .A(\regfile_i[WRITE_DATA][13] ), .B(n2494), .C(n2492), 
        .D(\registers[4][13] ), .Z(n1543) );
  HS65_LH_AO22X9 U2819 ( .A(\regfile_i[WRITE_DATA][14] ), .B(n2494), .C(n2492), 
        .D(\registers[4][14] ), .Z(n1544) );
  HS65_LH_AO22X9 U2820 ( .A(\regfile_i[WRITE_DATA][15] ), .B(n2494), .C(n2492), 
        .D(\registers[4][15] ), .Z(n1545) );
  HS65_LH_AO22X9 U2821 ( .A(\regfile_i[WRITE_DATA][16] ), .B(n2494), .C(n2492), 
        .D(\registers[4][16] ), .Z(n1546) );
  HS65_LH_AO22X9 U2822 ( .A(\regfile_i[WRITE_DATA][17] ), .B(n2494), .C(n2492), 
        .D(\registers[4][17] ), .Z(n1547) );
  HS65_LH_AO22X9 U2823 ( .A(\regfile_i[WRITE_DATA][18] ), .B(n2494), .C(n2492), 
        .D(\registers[4][18] ), .Z(n1548) );
  HS65_LH_AO22X9 U2824 ( .A(\regfile_i[WRITE_DATA][19] ), .B(n2494), .C(n2491), 
        .D(\registers[4][19] ), .Z(n1549) );
  HS65_LH_AO22X9 U2825 ( .A(\regfile_i[WRITE_DATA][20] ), .B(n2494), .C(n2491), 
        .D(\registers[4][20] ), .Z(n1550) );
  HS65_LH_AO22X9 U2826 ( .A(\regfile_i[WRITE_DATA][21] ), .B(n2494), .C(n2491), 
        .D(\registers[4][21] ), .Z(n1551) );
  HS65_LH_AO22X9 U2827 ( .A(\regfile_i[WRITE_DATA][22] ), .B(n2494), .C(n2491), 
        .D(\registers[4][22] ), .Z(n1552) );
  HS65_LH_AO22X9 U2828 ( .A(\regfile_i[WRITE_DATA][23] ), .B(n2494), .C(n2491), 
        .D(\registers[4][23] ), .Z(n1553) );
  HS65_LH_AO22X9 U2829 ( .A(\regfile_i[WRITE_DATA][24] ), .B(n2494), .C(n2491), 
        .D(\registers[4][24] ), .Z(n1554) );
  HS65_LH_AO22X9 U2830 ( .A(\regfile_i[WRITE_DATA][25] ), .B(n2494), .C(n2491), 
        .D(\registers[4][25] ), .Z(n1555) );
  HS65_LH_AO22X9 U2831 ( .A(\regfile_i[WRITE_DATA][26] ), .B(n2494), .C(n2491), 
        .D(\registers[4][26] ), .Z(n1556) );
  HS65_LH_AO22X9 U2832 ( .A(\regfile_i[WRITE_DATA][27] ), .B(n2494), .C(n2491), 
        .D(\registers[4][27] ), .Z(n1557) );
  HS65_LH_AO22X9 U2833 ( .A(\regfile_i[WRITE_DATA][28] ), .B(n2494), .C(n2491), 
        .D(\registers[4][28] ), .Z(n1558) );
  HS65_LH_AO22X9 U2834 ( .A(\regfile_i[WRITE_DATA][29] ), .B(n2494), .C(n2491), 
        .D(\registers[4][29] ), .Z(n1559) );
  HS65_LH_AO22X9 U2835 ( .A(\regfile_i[WRITE_DATA][30] ), .B(n2494), .C(n2491), 
        .D(\registers[4][30] ), .Z(n1560) );
  HS65_LH_AO22X9 U2836 ( .A(\regfile_i[WRITE_DATA][31] ), .B(n2493), .C(n2491), 
        .D(\registers[4][31] ), .Z(n1561) );
  HS65_LH_AO22X9 U2837 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n2434), .C(n2431), 
        .D(\registers[16][0] ), .Z(n1914) );
  HS65_LH_AO22X9 U2838 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n2434), .C(n2431), 
        .D(\registers[16][1] ), .Z(n1915) );
  HS65_LH_AO22X9 U2839 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n2434), .C(n2431), 
        .D(\registers[16][2] ), .Z(n1916) );
  HS65_LH_AO22X9 U2840 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n2434), .C(n2431), 
        .D(\registers[16][3] ), .Z(n1917) );
  HS65_LH_AO22X9 U2841 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n2434), .C(n2431), 
        .D(\registers[16][4] ), .Z(n1918) );
  HS65_LH_AO22X9 U2842 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n2434), .C(n2431), 
        .D(\registers[16][5] ), .Z(n1919) );
  HS65_LH_AO22X9 U2843 ( .A(n2709), .B(n2434), .C(n2431), .D(
        \registers[16][6] ), .Z(n1920) );
  HS65_LH_AO22X9 U2844 ( .A(n2711), .B(n2434), .C(n2431), .D(
        \registers[16][7] ), .Z(n1921) );
  HS65_LH_AO22X9 U2845 ( .A(n2713), .B(n2434), .C(n2431), .D(
        \registers[16][8] ), .Z(n1922) );
  HS65_LH_AO22X9 U2846 ( .A(n2715), .B(n2434), .C(n2431), .D(
        \registers[16][9] ), .Z(n1923) );
  HS65_LH_AO22X9 U2847 ( .A(n2717), .B(n2434), .C(n2431), .D(
        \registers[16][10] ), .Z(n1924) );
  HS65_LH_AO22X9 U2848 ( .A(n2719), .B(n2433), .C(n2431), .D(
        \registers[16][11] ), .Z(n1925) );
  HS65_LH_AO22X9 U2849 ( .A(n2721), .B(n2433), .C(n2431), .D(
        \registers[16][12] ), .Z(n1926) );
  HS65_LH_AO22X9 U2850 ( .A(n2723), .B(n2433), .C(n2431), .D(
        \registers[16][13] ), .Z(n1927) );
  HS65_LH_AO22X9 U2851 ( .A(n2725), .B(n2433), .C(n2431), .D(
        \registers[16][14] ), .Z(n1928) );
  HS65_LH_AO22X9 U2852 ( .A(n2727), .B(n2433), .C(n2431), .D(
        \registers[16][15] ), .Z(n1929) );
  HS65_LH_AO22X9 U2853 ( .A(n2729), .B(n2433), .C(n2431), .D(
        \registers[16][16] ), .Z(n1930) );
  HS65_LH_AO22X9 U2854 ( .A(n2731), .B(n2433), .C(n2431), .D(
        \registers[16][17] ), .Z(n1931) );
  HS65_LH_AO22X9 U2855 ( .A(n2733), .B(n2433), .C(n2431), .D(
        \registers[16][18] ), .Z(n1932) );
  HS65_LH_AO22X9 U2856 ( .A(n2735), .B(n2433), .C(n2431), .D(
        \registers[16][19] ), .Z(n1933) );
  HS65_LH_AO22X9 U2857 ( .A(n2737), .B(n2433), .C(n1416), .D(
        \registers[16][20] ), .Z(n1934) );
  HS65_LH_AO22X9 U2858 ( .A(n2739), .B(n2433), .C(n1416), .D(
        \registers[16][21] ), .Z(n1935) );
  HS65_LH_AO22X9 U2859 ( .A(n2741), .B(n2433), .C(n1416), .D(
        \registers[16][22] ), .Z(n1936) );
  HS65_LH_AO22X9 U2860 ( .A(n2743), .B(n2433), .C(n1416), .D(
        \registers[16][23] ), .Z(n1937) );
  HS65_LH_AO22X9 U2861 ( .A(n2745), .B(n2433), .C(n1416), .D(
        \registers[16][24] ), .Z(n1938) );
  HS65_LH_AO22X9 U2862 ( .A(n2747), .B(n2433), .C(n1416), .D(
        \registers[16][25] ), .Z(n1939) );
  HS65_LH_AO22X9 U2863 ( .A(n2749), .B(n2433), .C(n1416), .D(
        \registers[16][26] ), .Z(n1940) );
  HS65_LH_AO22X9 U2864 ( .A(n2751), .B(n2433), .C(n1416), .D(
        \registers[16][27] ), .Z(n1941) );
  HS65_LH_AO22X9 U2865 ( .A(n2753), .B(n2433), .C(n1416), .D(
        \registers[16][28] ), .Z(n1942) );
  HS65_LH_AO22X9 U2866 ( .A(n2755), .B(n2433), .C(n1416), .D(
        \registers[16][29] ), .Z(n1943) );
  HS65_LH_AO22X9 U2867 ( .A(n2757), .B(n2433), .C(n1416), .D(
        \registers[16][30] ), .Z(n1944) );
  HS65_LH_AO22X9 U2868 ( .A(n2759), .B(n2432), .C(n1416), .D(
        \registers[16][31] ), .Z(n1945) );
  HS65_LH_AO22X9 U2869 ( .A(\regfile_i[WRITE_DATA][0] ), .B(n1413), .C(n1410), 
        .D(\registers[20][0] ), .Z(n2042) );
  HS65_LH_AO22X9 U2870 ( .A(\regfile_i[WRITE_DATA][1] ), .B(n1413), .C(n1405), 
        .D(\registers[20][1] ), .Z(n2043) );
  HS65_LH_AO22X9 U2871 ( .A(\regfile_i[WRITE_DATA][2] ), .B(n1413), .C(n1410), 
        .D(\registers[20][2] ), .Z(n2044) );
  HS65_LH_AO22X9 U2872 ( .A(\regfile_i[WRITE_DATA][3] ), .B(n1413), .C(n1405), 
        .D(\registers[20][3] ), .Z(n2045) );
  HS65_LH_AO22X9 U2873 ( .A(\regfile_i[WRITE_DATA][4] ), .B(n1413), .C(n1410), 
        .D(\registers[20][4] ), .Z(n2046) );
  HS65_LH_AO22X9 U2874 ( .A(\regfile_i[WRITE_DATA][5] ), .B(n1413), .C(n1405), 
        .D(\registers[20][5] ), .Z(n2047) );
  HS65_LH_AO22X9 U2875 ( .A(n2709), .B(n1413), .C(n1410), .D(
        \registers[20][6] ), .Z(n2048) );
  HS65_LH_AO22X9 U2876 ( .A(n2711), .B(n1413), .C(n1410), .D(
        \registers[20][7] ), .Z(n2049) );
  HS65_LH_AO22X9 U2877 ( .A(n2713), .B(n1413), .C(n1410), .D(
        \registers[20][8] ), .Z(n2050) );
  HS65_LH_AO22X9 U2878 ( .A(n2715), .B(n1413), .C(n1410), .D(
        \registers[20][9] ), .Z(n2051) );
  HS65_LH_AO22X9 U2879 ( .A(n2717), .B(n1413), .C(n1410), .D(
        \registers[20][10] ), .Z(n2052) );
  HS65_LH_AO22X9 U2880 ( .A(n2719), .B(n1412), .C(n1410), .D(
        \registers[20][11] ), .Z(n2053) );
  HS65_LH_AO22X9 U2881 ( .A(n2721), .B(n1412), .C(n1410), .D(
        \registers[20][12] ), .Z(n2054) );
  HS65_LH_AO22X9 U2882 ( .A(n2723), .B(n1412), .C(n1410), .D(
        \registers[20][13] ), .Z(n2055) );
  HS65_LH_AO22X9 U2883 ( .A(n2725), .B(n1412), .C(n1410), .D(
        \registers[20][14] ), .Z(n2056) );
  HS65_LH_AO22X9 U2884 ( .A(n2727), .B(n1412), .C(n1410), .D(
        \registers[20][15] ), .Z(n2057) );
  HS65_LH_AO22X9 U2885 ( .A(n2729), .B(n1412), .C(n1410), .D(
        \registers[20][16] ), .Z(n2058) );
  HS65_LH_AO22X9 U2886 ( .A(n2731), .B(n1412), .C(n1410), .D(
        \registers[20][17] ), .Z(n2059) );
  HS65_LH_AO22X9 U2887 ( .A(n2733), .B(n1412), .C(n1410), .D(
        \registers[20][18] ), .Z(n2060) );
  HS65_LH_AO22X9 U2888 ( .A(n2735), .B(n1412), .C(n1405), .D(
        \registers[20][19] ), .Z(n2061) );
  HS65_LH_AO22X9 U2889 ( .A(n2737), .B(n1412), .C(n1405), .D(
        \registers[20][20] ), .Z(n2062) );
  HS65_LH_AO22X9 U2890 ( .A(n2739), .B(n1412), .C(n1405), .D(
        \registers[20][21] ), .Z(n2063) );
  HS65_LH_AO22X9 U2891 ( .A(n2741), .B(n1412), .C(n1405), .D(
        \registers[20][22] ), .Z(n2064) );
  HS65_LH_AO22X9 U2892 ( .A(n2743), .B(n1412), .C(n1405), .D(
        \registers[20][23] ), .Z(n2065) );
  HS65_LH_AO22X9 U2893 ( .A(n2745), .B(n1412), .C(n1405), .D(
        \registers[20][24] ), .Z(n2066) );
  HS65_LH_AO22X9 U2894 ( .A(n2747), .B(n1412), .C(n1405), .D(
        \registers[20][25] ), .Z(n2067) );
  HS65_LH_AO22X9 U2895 ( .A(n2749), .B(n1412), .C(n1405), .D(
        \registers[20][26] ), .Z(n2068) );
  HS65_LH_AO22X9 U2896 ( .A(n2751), .B(n1412), .C(n1405), .D(
        \registers[20][27] ), .Z(n2069) );
  HS65_LH_AO22X9 U2897 ( .A(n2753), .B(n1412), .C(n1405), .D(
        \registers[20][28] ), .Z(n2070) );
  HS65_LH_AO22X9 U2898 ( .A(n2755), .B(n1412), .C(n1405), .D(
        \registers[20][29] ), .Z(n2071) );
  HS65_LH_AO22X9 U2899 ( .A(n2757), .B(n1412), .C(n1405), .D(
        \registers[20][30] ), .Z(n2072) );
  HS65_LH_AO22X9 U2900 ( .A(n2759), .B(n1411), .C(n1405), .D(
        \registers[20][31] ), .Z(n2073) );
  HS65_LH_NOR3X4 U2901 ( .A(\regfile_i[ADRWRITE][0] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(n2896), .Z(n1396) );
  HS65_LH_NOR3X4 U2902 ( .A(n2897), .B(\regfile_i[ADRWRITE][2] ), .C(n2896), 
        .Z(n1398) );
  HS65_LH_NOR3X4 U2903 ( .A(\regfile_i[ADRWRITE][1] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(n2897), .Z(n1393) );
  HS65_LH_IVX9 U2904 ( .A(\regfile_i[ADRWRITE][0] ), .Z(n2897) );
  HS65_LH_IVX9 U2905 ( .A(\regfile_i[ADRWRITE][1] ), .Z(n2896) );
  HS65_LH_IVX9 U2906 ( .A(\regfile_i[ADRWRITE][3] ), .Z(n2895) );
  HS65_LH_NOR3X4 U2907 ( .A(\regfile_i[ADRWRITE][1] ), .B(
        \regfile_i[ADRWRITE][2] ), .C(\regfile_i[ADRWRITE][0] ), .Z(n1391) );
  HS65_LH_AND3X9 U2908 ( .A(\regfile_i[WR_EN] ), .B(n2895), .C(
        \regfile_i[ADRWRITE][4] ), .Z(n1417) );
  HS65_LH_AND3X9 U2909 ( .A(\regfile_i[ADRWRITE][3] ), .B(\regfile_i[WR_EN] ), 
        .C(\regfile_i[ADRWRITE][4] ), .Z(n1426) );
endmodule


module id_top ( clk, rst_n, .id_top_i({\id_top_i[INSTRUCTION][31] , 
        \id_top_i[INSTRUCTION][30] , \id_top_i[INSTRUCTION][29] , 
        \id_top_i[INSTRUCTION][28] , \id_top_i[INSTRUCTION][27] , 
        \id_top_i[INSTRUCTION][26] , \id_top_i[INSTRUCTION][25] , 
        \id_top_i[INSTRUCTION][24] , \id_top_i[INSTRUCTION][23] , 
        \id_top_i[INSTRUCTION][22] , \id_top_i[INSTRUCTION][21] , 
        \id_top_i[INSTRUCTION][20] , \id_top_i[INSTRUCTION][19] , 
        \id_top_i[INSTRUCTION][18] , \id_top_i[INSTRUCTION][17] , 
        \id_top_i[INSTRUCTION][16] , \id_top_i[INSTRUCTION][15] , 
        \id_top_i[INSTRUCTION][14] , \id_top_i[INSTRUCTION][13] , 
        \id_top_i[INSTRUCTION][12] , \id_top_i[INSTRUCTION][11] , 
        \id_top_i[INSTRUCTION][10] , \id_top_i[INSTRUCTION][9] , 
        \id_top_i[INSTRUCTION][8] , \id_top_i[INSTRUCTION][7] , 
        \id_top_i[INSTRUCTION][6] , \id_top_i[INSTRUCTION][5] , 
        \id_top_i[INSTRUCTION][4] , \id_top_i[INSTRUCTION][3] , 
        \id_top_i[INSTRUCTION][2] , \id_top_i[INSTRUCTION][1] , 
        \id_top_i[INSTRUCTION][0] , \id_top_i[WRITEBACK_DATA][31] , 
        \id_top_i[WRITEBACK_DATA][30] , \id_top_i[WRITEBACK_DATA][29] , 
        \id_top_i[WRITEBACK_DATA][28] , \id_top_i[WRITEBACK_DATA][27] , 
        \id_top_i[WRITEBACK_DATA][26] , \id_top_i[WRITEBACK_DATA][25] , 
        \id_top_i[WRITEBACK_DATA][24] , \id_top_i[WRITEBACK_DATA][23] , 
        \id_top_i[WRITEBACK_DATA][22] , \id_top_i[WRITEBACK_DATA][21] , 
        \id_top_i[WRITEBACK_DATA][20] , \id_top_i[WRITEBACK_DATA][19] , 
        \id_top_i[WRITEBACK_DATA][18] , \id_top_i[WRITEBACK_DATA][17] , 
        \id_top_i[WRITEBACK_DATA][16] , \id_top_i[WRITEBACK_DATA][15] , 
        \id_top_i[WRITEBACK_DATA][14] , \id_top_i[WRITEBACK_DATA][13] , 
        \id_top_i[WRITEBACK_DATA][12] , \id_top_i[WRITEBACK_DATA][11] , 
        \id_top_i[WRITEBACK_DATA][10] , \id_top_i[WRITEBACK_DATA][9] , 
        \id_top_i[WRITEBACK_DATA][8] , \id_top_i[WRITEBACK_DATA][7] , 
        \id_top_i[WRITEBACK_DATA][6] , \id_top_i[WRITEBACK_DATA][5] , 
        \id_top_i[WRITEBACK_DATA][4] , \id_top_i[WRITEBACK_DATA][3] , 
        \id_top_i[WRITEBACK_DATA][2] , \id_top_i[WRITEBACK_DATA][1] , 
        \id_top_i[WRITEBACK_DATA][0] , \id_top_i[FORWARD_A] , 
        \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] , \id_top_i[WRITE_REG][4] , 
        \id_top_i[WRITE_REG][3] , \id_top_i[WRITE_REG][2] , 
        \id_top_i[WRITE_REG][1] , \id_top_i[WRITE_REG][0] }), .id_top_o({
        \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] , 
        \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] , 
        \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] , 
        \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] , 
        \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] , 
        \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] , 
        \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] , 
        \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] , 
        \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] , 
        \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] , 
        \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] , 
        \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] , 
        \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] , 
        \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] , 
        \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] , 
        \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] , 
        \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] , 
        \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] , 
        \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] , 
        \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] , 
        \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] , 
        \id_top_o[REG_B][0] , \id_top_o[INSTR_31_26][5] , 
        \id_top_o[INSTR_31_26][4] , \id_top_o[INSTR_31_26][3] , 
        \id_top_o[INSTR_31_26][2] , \id_top_o[INSTR_31_26][1] , 
        \id_top_o[INSTR_31_26][0] , \id_top_o[RS][4] , \id_top_o[RS][3] , 
        \id_top_o[RS][2] , \id_top_o[RS][1] , \id_top_o[RS][0] , 
        \id_top_o[RT][4] , \id_top_o[RT][3] , \id_top_o[RT][2] , 
        \id_top_o[RT][1] , \id_top_o[RT][0] , \id_top_o[RD][4] , 
        \id_top_o[RD][3] , \id_top_o[RD][2] , \id_top_o[RD][1] , 
        \id_top_o[RD][0] , \id_top_o[INSTR_10_6][4] , 
        \id_top_o[INSTR_10_6][3] , \id_top_o[INSTR_10_6][2] , 
        \id_top_o[INSTR_10_6][1] , \id_top_o[INSTR_10_6][0] , 
        \id_top_o[INSTR_5_0][5] , \id_top_o[INSTR_5_0][4] , 
        \id_top_o[INSTR_5_0][3] , \id_top_o[INSTR_5_0][2] , 
        \id_top_o[INSTR_5_0][1] , \id_top_o[INSTR_5_0][0] , 
        \id_top_o[SIGN_EXTEND][31] , \id_top_o[SIGN_EXTEND][30] , 
        \id_top_o[SIGN_EXTEND][29] , \id_top_o[SIGN_EXTEND][28] , 
        \id_top_o[SIGN_EXTEND][27] , \id_top_o[SIGN_EXTEND][26] , 
        \id_top_o[SIGN_EXTEND][25] , \id_top_o[SIGN_EXTEND][24] , 
        \id_top_o[SIGN_EXTEND][23] , \id_top_o[SIGN_EXTEND][22] , 
        \id_top_o[SIGN_EXTEND][21] , \id_top_o[SIGN_EXTEND][20] , 
        \id_top_o[SIGN_EXTEND][19] , \id_top_o[SIGN_EXTEND][18] , 
        \id_top_o[SIGN_EXTEND][17] , \id_top_o[SIGN_EXTEND][16] , 
        \id_top_o[SIGN_EXTEND][15] , \id_top_o[SIGN_EXTEND][14] , 
        \id_top_o[SIGN_EXTEND][13] , \id_top_o[SIGN_EXTEND][12] , 
        \id_top_o[SIGN_EXTEND][11] , \id_top_o[SIGN_EXTEND][10] , 
        \id_top_o[SIGN_EXTEND][9] , \id_top_o[SIGN_EXTEND][8] , 
        \id_top_o[SIGN_EXTEND][7] , \id_top_o[SIGN_EXTEND][6] , 
        \id_top_o[SIGN_EXTEND][5] , \id_top_o[SIGN_EXTEND][4] , 
        \id_top_o[SIGN_EXTEND][3] , \id_top_o[SIGN_EXTEND][2] , 
        \id_top_o[SIGN_EXTEND][1] , \id_top_o[SIGN_EXTEND][0] }) );
  input clk, rst_n, \id_top_i[INSTRUCTION][31] , \id_top_i[INSTRUCTION][30] ,
         \id_top_i[INSTRUCTION][29] , \id_top_i[INSTRUCTION][28] ,
         \id_top_i[INSTRUCTION][27] , \id_top_i[INSTRUCTION][26] ,
         \id_top_i[INSTRUCTION][25] , \id_top_i[INSTRUCTION][24] ,
         \id_top_i[INSTRUCTION][23] , \id_top_i[INSTRUCTION][22] ,
         \id_top_i[INSTRUCTION][21] , \id_top_i[INSTRUCTION][20] ,
         \id_top_i[INSTRUCTION][19] , \id_top_i[INSTRUCTION][18] ,
         \id_top_i[INSTRUCTION][17] , \id_top_i[INSTRUCTION][16] ,
         \id_top_i[INSTRUCTION][15] , \id_top_i[INSTRUCTION][14] ,
         \id_top_i[INSTRUCTION][13] , \id_top_i[INSTRUCTION][12] ,
         \id_top_i[INSTRUCTION][11] , \id_top_i[INSTRUCTION][10] ,
         \id_top_i[INSTRUCTION][9] , \id_top_i[INSTRUCTION][8] ,
         \id_top_i[INSTRUCTION][7] , \id_top_i[INSTRUCTION][6] ,
         \id_top_i[INSTRUCTION][5] , \id_top_i[INSTRUCTION][4] ,
         \id_top_i[INSTRUCTION][3] , \id_top_i[INSTRUCTION][2] ,
         \id_top_i[INSTRUCTION][1] , \id_top_i[INSTRUCTION][0] ,
         \id_top_i[WRITEBACK_DATA][31] , \id_top_i[WRITEBACK_DATA][30] ,
         \id_top_i[WRITEBACK_DATA][29] , \id_top_i[WRITEBACK_DATA][28] ,
         \id_top_i[WRITEBACK_DATA][27] , \id_top_i[WRITEBACK_DATA][26] ,
         \id_top_i[WRITEBACK_DATA][25] , \id_top_i[WRITEBACK_DATA][24] ,
         \id_top_i[WRITEBACK_DATA][23] , \id_top_i[WRITEBACK_DATA][22] ,
         \id_top_i[WRITEBACK_DATA][21] , \id_top_i[WRITEBACK_DATA][20] ,
         \id_top_i[WRITEBACK_DATA][19] , \id_top_i[WRITEBACK_DATA][18] ,
         \id_top_i[WRITEBACK_DATA][17] , \id_top_i[WRITEBACK_DATA][16] ,
         \id_top_i[WRITEBACK_DATA][15] , \id_top_i[WRITEBACK_DATA][14] ,
         \id_top_i[WRITEBACK_DATA][13] , \id_top_i[WRITEBACK_DATA][12] ,
         \id_top_i[WRITEBACK_DATA][11] , \id_top_i[WRITEBACK_DATA][10] ,
         \id_top_i[WRITEBACK_DATA][9] , \id_top_i[WRITEBACK_DATA][8] ,
         \id_top_i[WRITEBACK_DATA][7] , \id_top_i[WRITEBACK_DATA][6] ,
         \id_top_i[WRITEBACK_DATA][5] , \id_top_i[WRITEBACK_DATA][4] ,
         \id_top_i[WRITEBACK_DATA][3] , \id_top_i[WRITEBACK_DATA][2] ,
         \id_top_i[WRITEBACK_DATA][1] , \id_top_i[WRITEBACK_DATA][0] ,
         \id_top_i[FORWARD_A] , \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] ,
         \id_top_i[WRITE_REG][4] , \id_top_i[WRITE_REG][3] ,
         \id_top_i[WRITE_REG][2] , \id_top_i[WRITE_REG][1] ,
         \id_top_i[WRITE_REG][0] ;
  output \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] ,
         \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] ,
         \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] ,
         \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] ,
         \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] ,
         \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] ,
         \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] ,
         \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] ,
         \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] ,
         \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] ,
         \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] ,
         \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] ,
         \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] ,
         \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] ,
         \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] ,
         \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] ,
         \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] ,
         \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] ,
         \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] ,
         \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] ,
         \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] ,
         \id_top_o[REG_B][0] , \id_top_o[INSTR_31_26][5] ,
         \id_top_o[INSTR_31_26][4] , \id_top_o[INSTR_31_26][3] ,
         \id_top_o[INSTR_31_26][2] , \id_top_o[INSTR_31_26][1] ,
         \id_top_o[INSTR_31_26][0] , \id_top_o[RS][4] , \id_top_o[RS][3] ,
         \id_top_o[RS][2] , \id_top_o[RS][1] , \id_top_o[RS][0] ,
         \id_top_o[RT][4] , \id_top_o[RT][3] , \id_top_o[RT][2] ,
         \id_top_o[RT][1] , \id_top_o[RT][0] , \id_top_o[RD][4] ,
         \id_top_o[RD][3] , \id_top_o[RD][2] , \id_top_o[RD][1] ,
         \id_top_o[RD][0] , \id_top_o[INSTR_10_6][4] ,
         \id_top_o[INSTR_10_6][3] , \id_top_o[INSTR_10_6][2] ,
         \id_top_o[INSTR_10_6][1] , \id_top_o[INSTR_10_6][0] ,
         \id_top_o[INSTR_5_0][5] , \id_top_o[INSTR_5_0][4] ,
         \id_top_o[INSTR_5_0][3] , \id_top_o[INSTR_5_0][2] ,
         \id_top_o[INSTR_5_0][1] , \id_top_o[INSTR_5_0][0] ,
         \id_top_o[SIGN_EXTEND][31] , \id_top_o[SIGN_EXTEND][30] ,
         \id_top_o[SIGN_EXTEND][29] , \id_top_o[SIGN_EXTEND][28] ,
         \id_top_o[SIGN_EXTEND][27] , \id_top_o[SIGN_EXTEND][26] ,
         \id_top_o[SIGN_EXTEND][25] , \id_top_o[SIGN_EXTEND][24] ,
         \id_top_o[SIGN_EXTEND][23] , \id_top_o[SIGN_EXTEND][22] ,
         \id_top_o[SIGN_EXTEND][21] , \id_top_o[SIGN_EXTEND][20] ,
         \id_top_o[SIGN_EXTEND][19] , \id_top_o[SIGN_EXTEND][18] ,
         \id_top_o[SIGN_EXTEND][17] , \id_top_o[SIGN_EXTEND][16] ,
         \id_top_o[SIGN_EXTEND][15] , \id_top_o[SIGN_EXTEND][14] ,
         \id_top_o[SIGN_EXTEND][13] , \id_top_o[SIGN_EXTEND][12] ,
         \id_top_o[SIGN_EXTEND][11] , \id_top_o[SIGN_EXTEND][10] ,
         \id_top_o[SIGN_EXTEND][9] , \id_top_o[SIGN_EXTEND][8] ,
         \id_top_o[SIGN_EXTEND][7] , \id_top_o[SIGN_EXTEND][6] ,
         \id_top_o[SIGN_EXTEND][5] , \id_top_o[SIGN_EXTEND][4] ,
         \id_top_o[SIGN_EXTEND][3] , \id_top_o[SIGN_EXTEND][2] ,
         \id_top_o[SIGN_EXTEND][1] , \id_top_o[SIGN_EXTEND][0] ;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96;

  regfile regfile_inst ( .clk(clk), .rst_n(rst_n), .regfile_i({
        \id_top_i[INSTRUCTION][25] , \id_top_i[INSTRUCTION][24] , 
        \id_top_i[INSTRUCTION][23] , \id_top_i[INSTRUCTION][22] , 
        \id_top_i[INSTRUCTION][21] , \id_top_i[INSTRUCTION][20] , 
        \id_top_i[INSTRUCTION][19] , \id_top_i[INSTRUCTION][18] , 
        \id_top_i[INSTRUCTION][17] , \id_top_i[INSTRUCTION][16] , 
        \id_top_i[WRITE_REG][4] , \id_top_i[WRITE_REG][3] , 
        \id_top_i[WRITE_REG][2] , \id_top_i[WRITE_REG][1] , 
        \id_top_i[WRITE_REG][0] , n96, n95, n94, n93, n92, n91, n90, n89, n88, 
        n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, 
        n73, n72, n71, n70, n69, n68, n67, n66, n65, \id_top_i[FORWARD_A] , 
        \id_top_i[FORWARD_B] , \id_top_i[REGWRITE] }), .regfile_o({
        \id_top_o[REG_A][31] , \id_top_o[REG_A][30] , \id_top_o[REG_A][29] , 
        \id_top_o[REG_A][28] , \id_top_o[REG_A][27] , \id_top_o[REG_A][26] , 
        \id_top_o[REG_A][25] , \id_top_o[REG_A][24] , \id_top_o[REG_A][23] , 
        \id_top_o[REG_A][22] , \id_top_o[REG_A][21] , \id_top_o[REG_A][20] , 
        \id_top_o[REG_A][19] , \id_top_o[REG_A][18] , \id_top_o[REG_A][17] , 
        \id_top_o[REG_A][16] , \id_top_o[REG_A][15] , \id_top_o[REG_A][14] , 
        \id_top_o[REG_A][13] , \id_top_o[REG_A][12] , \id_top_o[REG_A][11] , 
        \id_top_o[REG_A][10] , \id_top_o[REG_A][9] , \id_top_o[REG_A][8] , 
        \id_top_o[REG_A][7] , \id_top_o[REG_A][6] , \id_top_o[REG_A][5] , 
        \id_top_o[REG_A][4] , \id_top_o[REG_A][3] , \id_top_o[REG_A][2] , 
        \id_top_o[REG_A][1] , \id_top_o[REG_A][0] , \id_top_o[REG_B][31] , 
        \id_top_o[REG_B][30] , \id_top_o[REG_B][29] , \id_top_o[REG_B][28] , 
        \id_top_o[REG_B][27] , \id_top_o[REG_B][26] , \id_top_o[REG_B][25] , 
        \id_top_o[REG_B][24] , \id_top_o[REG_B][23] , \id_top_o[REG_B][22] , 
        \id_top_o[REG_B][21] , \id_top_o[REG_B][20] , \id_top_o[REG_B][19] , 
        \id_top_o[REG_B][18] , \id_top_o[REG_B][17] , \id_top_o[REG_B][16] , 
        \id_top_o[REG_B][15] , \id_top_o[REG_B][14] , \id_top_o[REG_B][13] , 
        \id_top_o[REG_B][12] , \id_top_o[REG_B][11] , \id_top_o[REG_B][10] , 
        \id_top_o[REG_B][9] , \id_top_o[REG_B][8] , \id_top_o[REG_B][7] , 
        \id_top_o[REG_B][6] , \id_top_o[REG_B][5] , \id_top_o[REG_B][4] , 
        \id_top_o[REG_B][3] , \id_top_o[REG_B][2] , \id_top_o[REG_B][1] , 
        \id_top_o[REG_B][0] }) );
  HS65_LH_BFX9 U1 ( .A(\id_top_i[WRITEBACK_DATA][0] ), .Z(n65) );
  HS65_LH_BFX9 U2 ( .A(\id_top_i[WRITEBACK_DATA][1] ), .Z(n66) );
  HS65_LH_BFX9 U3 ( .A(\id_top_i[WRITEBACK_DATA][2] ), .Z(n67) );
  HS65_LH_BFX9 U4 ( .A(\id_top_i[WRITEBACK_DATA][3] ), .Z(n68) );
  HS65_LH_BFX9 U5 ( .A(\id_top_i[WRITEBACK_DATA][4] ), .Z(n69) );
  HS65_LH_BFX9 U6 ( .A(\id_top_i[WRITEBACK_DATA][5] ), .Z(n70) );
  HS65_LH_BFX9 U7 ( .A(\id_top_i[WRITEBACK_DATA][6] ), .Z(n71) );
  HS65_LH_BFX9 U8 ( .A(\id_top_i[WRITEBACK_DATA][7] ), .Z(n72) );
  HS65_LH_BFX9 U9 ( .A(\id_top_i[WRITEBACK_DATA][8] ), .Z(n73) );
  HS65_LH_BFX9 U10 ( .A(\id_top_i[WRITEBACK_DATA][9] ), .Z(n74) );
  HS65_LH_BFX9 U11 ( .A(\id_top_i[WRITEBACK_DATA][10] ), .Z(n75) );
  HS65_LH_BFX9 U12 ( .A(\id_top_i[WRITEBACK_DATA][11] ), .Z(n76) );
  HS65_LH_BFX9 U13 ( .A(\id_top_i[WRITEBACK_DATA][12] ), .Z(n77) );
  HS65_LH_BFX9 U14 ( .A(\id_top_i[WRITEBACK_DATA][13] ), .Z(n78) );
  HS65_LH_BFX9 U15 ( .A(\id_top_i[WRITEBACK_DATA][14] ), .Z(n79) );
  HS65_LH_BFX9 U16 ( .A(\id_top_i[WRITEBACK_DATA][15] ), .Z(n80) );
  HS65_LH_BFX9 U17 ( .A(\id_top_i[WRITEBACK_DATA][16] ), .Z(n81) );
  HS65_LH_BFX9 U18 ( .A(\id_top_i[WRITEBACK_DATA][17] ), .Z(n82) );
  HS65_LH_BFX9 U19 ( .A(\id_top_i[WRITEBACK_DATA][18] ), .Z(n83) );
  HS65_LH_BFX9 U20 ( .A(\id_top_i[WRITEBACK_DATA][19] ), .Z(n84) );
  HS65_LH_BFX9 U21 ( .A(\id_top_i[WRITEBACK_DATA][20] ), .Z(n85) );
  HS65_LH_BFX9 U22 ( .A(\id_top_i[WRITEBACK_DATA][21] ), .Z(n86) );
  HS65_LH_BFX9 U23 ( .A(\id_top_i[WRITEBACK_DATA][22] ), .Z(n87) );
  HS65_LH_BFX9 U24 ( .A(\id_top_i[WRITEBACK_DATA][23] ), .Z(n88) );
  HS65_LH_BFX9 U25 ( .A(\id_top_i[WRITEBACK_DATA][24] ), .Z(n89) );
  HS65_LH_BFX9 U26 ( .A(\id_top_i[WRITEBACK_DATA][25] ), .Z(n90) );
  HS65_LH_BFX9 U27 ( .A(\id_top_i[WRITEBACK_DATA][26] ), .Z(n91) );
  HS65_LH_BFX9 U28 ( .A(\id_top_i[WRITEBACK_DATA][27] ), .Z(n92) );
  HS65_LH_BFX9 U29 ( .A(\id_top_i[WRITEBACK_DATA][28] ), .Z(n93) );
  HS65_LH_BFX9 U30 ( .A(\id_top_i[WRITEBACK_DATA][29] ), .Z(n94) );
  HS65_LH_BFX9 U31 ( .A(\id_top_i[WRITEBACK_DATA][30] ), .Z(n95) );
  HS65_LH_BFX9 U32 ( .A(\id_top_i[WRITEBACK_DATA][31] ), .Z(n96) );
  HS65_LH_BFX9 U33 ( .A(\id_top_i[INSTRUCTION][11] ), .Z(\id_top_o[RD][0] ) );
  HS65_LH_BFX9 U34 ( .A(\id_top_i[INSTRUCTION][12] ), .Z(\id_top_o[RD][1] ) );
  HS65_LH_BFX9 U35 ( .A(\id_top_i[INSTRUCTION][13] ), .Z(\id_top_o[RD][2] ) );
  HS65_LH_BFX9 U36 ( .A(\id_top_i[INSTRUCTION][14] ), .Z(\id_top_o[RD][3] ) );
  HS65_LH_BFX9 U37 ( .A(\id_top_i[INSTRUCTION][0] ), .Z(
        \id_top_o[SIGN_EXTEND][0] ) );
  HS65_LH_BFX9 U38 ( .A(\id_top_i[INSTRUCTION][1] ), .Z(
        \id_top_o[SIGN_EXTEND][1] ) );
  HS65_LH_BFX9 U39 ( .A(\id_top_i[INSTRUCTION][2] ), .Z(
        \id_top_o[SIGN_EXTEND][2] ) );
  HS65_LH_BFX9 U40 ( .A(\id_top_i[INSTRUCTION][3] ), .Z(
        \id_top_o[SIGN_EXTEND][3] ) );
  HS65_LH_BFX9 U41 ( .A(\id_top_i[INSTRUCTION][4] ), .Z(
        \id_top_o[SIGN_EXTEND][4] ) );
  HS65_LH_BFX9 U42 ( .A(\id_top_i[INSTRUCTION][5] ), .Z(
        \id_top_o[SIGN_EXTEND][5] ) );
  HS65_LH_BFX9 U43 ( .A(\id_top_i[INSTRUCTION][6] ), .Z(
        \id_top_o[SIGN_EXTEND][6] ) );
  HS65_LH_BFX9 U44 ( .A(\id_top_i[INSTRUCTION][7] ), .Z(
        \id_top_o[SIGN_EXTEND][7] ) );
  HS65_LH_BFX9 U45 ( .A(\id_top_i[INSTRUCTION][8] ), .Z(
        \id_top_o[SIGN_EXTEND][8] ) );
  HS65_LH_BFX9 U46 ( .A(\id_top_i[INSTRUCTION][9] ), .Z(
        \id_top_o[SIGN_EXTEND][9] ) );
  HS65_LH_BFX9 U47 ( .A(\id_top_i[INSTRUCTION][10] ), .Z(
        \id_top_o[SIGN_EXTEND][10] ) );
  HS65_LH_BFX9 U48 ( .A(\id_top_i[INSTRUCTION][11] ), .Z(
        \id_top_o[SIGN_EXTEND][11] ) );
  HS65_LH_BFX9 U49 ( .A(\id_top_i[INSTRUCTION][12] ), .Z(
        \id_top_o[SIGN_EXTEND][12] ) );
  HS65_LH_BFX9 U50 ( .A(\id_top_i[INSTRUCTION][13] ), .Z(
        \id_top_o[SIGN_EXTEND][13] ) );
  HS65_LH_BFX9 U51 ( .A(\id_top_i[INSTRUCTION][14] ), .Z(
        \id_top_o[SIGN_EXTEND][14] ) );
  HS65_LH_BFX9 U52 ( .A(\id_top_i[INSTRUCTION][0] ), .Z(
        \id_top_o[INSTR_5_0][0] ) );
  HS65_LH_BFX9 U53 ( .A(\id_top_i[INSTRUCTION][1] ), .Z(
        \id_top_o[INSTR_5_0][1] ) );
  HS65_LH_BFX9 U54 ( .A(\id_top_i[INSTRUCTION][2] ), .Z(
        \id_top_o[INSTR_5_0][2] ) );
  HS65_LH_BFX9 U55 ( .A(\id_top_i[INSTRUCTION][3] ), .Z(
        \id_top_o[INSTR_5_0][3] ) );
  HS65_LH_BFX9 U56 ( .A(\id_top_i[INSTRUCTION][4] ), .Z(
        \id_top_o[INSTR_5_0][4] ) );
  HS65_LH_BFX9 U57 ( .A(\id_top_i[INSTRUCTION][5] ), .Z(
        \id_top_o[INSTR_5_0][5] ) );
  HS65_LH_BFX9 U58 ( .A(\id_top_i[INSTRUCTION][6] ), .Z(
        \id_top_o[INSTR_10_6][0] ) );
  HS65_LH_BFX9 U59 ( .A(\id_top_i[INSTRUCTION][7] ), .Z(
        \id_top_o[INSTR_10_6][1] ) );
  HS65_LH_BFX9 U60 ( .A(\id_top_i[INSTRUCTION][8] ), .Z(
        \id_top_o[INSTR_10_6][2] ) );
  HS65_LH_BFX9 U61 ( .A(\id_top_i[INSTRUCTION][9] ), .Z(
        \id_top_o[INSTR_10_6][3] ) );
  HS65_LH_BFX9 U62 ( .A(\id_top_i[INSTRUCTION][10] ), .Z(
        \id_top_o[INSTR_10_6][4] ) );
  HS65_LH_BFX9 U63 ( .A(\id_top_i[INSTRUCTION][31] ), .Z(
        \id_top_o[INSTR_31_26][5] ) );
  HS65_LH_BFX9 U64 ( .A(\id_top_i[INSTRUCTION][30] ), .Z(
        \id_top_o[INSTR_31_26][4] ) );
  HS65_LH_BFX9 U65 ( .A(\id_top_i[INSTRUCTION][29] ), .Z(
        \id_top_o[INSTR_31_26][3] ) );
  HS65_LH_BFX9 U66 ( .A(\id_top_i[INSTRUCTION][28] ), .Z(
        \id_top_o[INSTR_31_26][2] ) );
  HS65_LH_BFX9 U67 ( .A(\id_top_i[INSTRUCTION][27] ), .Z(
        \id_top_o[INSTR_31_26][1] ) );
  HS65_LH_BFX9 U68 ( .A(\id_top_i[INSTRUCTION][26] ), .Z(
        \id_top_o[INSTR_31_26][0] ) );
  HS65_LH_BFX9 U69 ( .A(\id_top_i[INSTRUCTION][25] ), .Z(\id_top_o[RS][4] ) );
  HS65_LH_BFX9 U70 ( .A(\id_top_i[INSTRUCTION][24] ), .Z(\id_top_o[RS][3] ) );
  HS65_LH_BFX9 U71 ( .A(\id_top_i[INSTRUCTION][23] ), .Z(\id_top_o[RS][2] ) );
  HS65_LH_BFX9 U72 ( .A(\id_top_i[INSTRUCTION][22] ), .Z(\id_top_o[RS][1] ) );
  HS65_LH_BFX9 U73 ( .A(\id_top_i[INSTRUCTION][21] ), .Z(\id_top_o[RS][0] ) );
  HS65_LH_BFX9 U74 ( .A(\id_top_i[INSTRUCTION][20] ), .Z(\id_top_o[RT][4] ) );
  HS65_LH_BFX9 U75 ( .A(\id_top_i[INSTRUCTION][19] ), .Z(\id_top_o[RT][3] ) );
  HS65_LH_BFX9 U76 ( .A(\id_top_i[INSTRUCTION][18] ), .Z(\id_top_o[RT][2] ) );
  HS65_LH_BFX9 U77 ( .A(\id_top_i[INSTRUCTION][17] ), .Z(\id_top_o[RT][1] ) );
  HS65_LH_BFX9 U78 ( .A(\id_top_i[INSTRUCTION][16] ), .Z(\id_top_o[RT][0] ) );
  HS65_LH_BFX9 U79 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][16] ) );
  HS65_LH_BFX9 U80 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][17] ) );
  HS65_LH_BFX9 U81 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][18] ) );
  HS65_LH_BFX9 U82 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][19] ) );
  HS65_LH_BFX9 U83 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][20] ) );
  HS65_LH_BFX9 U84 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][21] ) );
  HS65_LH_BFX9 U85 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][22] ) );
  HS65_LH_BFX9 U86 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][23] ) );
  HS65_LH_BFX9 U87 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][24] ) );
  HS65_LH_BFX9 U88 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][25] ) );
  HS65_LH_BFX9 U89 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][26] ) );
  HS65_LH_BFX9 U90 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][27] ) );
  HS65_LH_BFX9 U91 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][28] ) );
  HS65_LH_BFX9 U92 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][29] ) );
  HS65_LH_BFX9 U93 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][30] ) );
  HS65_LH_BFX9 U94 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][31] ) );
  HS65_LH_BFX9 U95 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(\id_top_o[RD][4] ) );
  HS65_LH_BFX9 U96 ( .A(\id_top_i[INSTRUCTION][15] ), .Z(
        \id_top_o[SIGN_EXTEND][15] ) );
endmodule


module id_exe ( clk, rst_n, halt_i, .ID_EXE_i({\ID_EXE_i[REGA][31] , 
        \ID_EXE_i[REGA][30] , \ID_EXE_i[REGA][29] , \ID_EXE_i[REGA][28] , 
        \ID_EXE_i[REGA][27] , \ID_EXE_i[REGA][26] , \ID_EXE_i[REGA][25] , 
        \ID_EXE_i[REGA][24] , \ID_EXE_i[REGA][23] , \ID_EXE_i[REGA][22] , 
        \ID_EXE_i[REGA][21] , \ID_EXE_i[REGA][20] , \ID_EXE_i[REGA][19] , 
        \ID_EXE_i[REGA][18] , \ID_EXE_i[REGA][17] , \ID_EXE_i[REGA][16] , 
        \ID_EXE_i[REGA][15] , \ID_EXE_i[REGA][14] , \ID_EXE_i[REGA][13] , 
        \ID_EXE_i[REGA][12] , \ID_EXE_i[REGA][11] , \ID_EXE_i[REGA][10] , 
        \ID_EXE_i[REGA][9] , \ID_EXE_i[REGA][8] , \ID_EXE_i[REGA][7] , 
        \ID_EXE_i[REGA][6] , \ID_EXE_i[REGA][5] , \ID_EXE_i[REGA][4] , 
        \ID_EXE_i[REGA][3] , \ID_EXE_i[REGA][2] , \ID_EXE_i[REGA][1] , 
        \ID_EXE_i[REGA][0] , \ID_EXE_i[REGB][31] , \ID_EXE_i[REGB][30] , 
        \ID_EXE_i[REGB][29] , \ID_EXE_i[REGB][28] , \ID_EXE_i[REGB][27] , 
        \ID_EXE_i[REGB][26] , \ID_EXE_i[REGB][25] , \ID_EXE_i[REGB][24] , 
        \ID_EXE_i[REGB][23] , \ID_EXE_i[REGB][22] , \ID_EXE_i[REGB][21] , 
        \ID_EXE_i[REGB][20] , \ID_EXE_i[REGB][19] , \ID_EXE_i[REGB][18] , 
        \ID_EXE_i[REGB][17] , \ID_EXE_i[REGB][16] , \ID_EXE_i[REGB][15] , 
        \ID_EXE_i[REGB][14] , \ID_EXE_i[REGB][13] , \ID_EXE_i[REGB][12] , 
        \ID_EXE_i[REGB][11] , \ID_EXE_i[REGB][10] , \ID_EXE_i[REGB][9] , 
        \ID_EXE_i[REGB][8] , \ID_EXE_i[REGB][7] , \ID_EXE_i[REGB][6] , 
        \ID_EXE_i[REGB][5] , \ID_EXE_i[REGB][4] , \ID_EXE_i[REGB][3] , 
        \ID_EXE_i[REGB][2] , \ID_EXE_i[REGB][1] , \ID_EXE_i[REGB][0] , 
        \ID_EXE_i[SHAMT][4] , \ID_EXE_i[SHAMT][3] , \ID_EXE_i[SHAMT][2] , 
        \ID_EXE_i[SHAMT][1] , \ID_EXE_i[SHAMT][0] , \ID_EXE_i[FUNCT][5] , 
        \ID_EXE_i[FUNCT][4] , \ID_EXE_i[FUNCT][3] , \ID_EXE_i[FUNCT][2] , 
        \ID_EXE_i[FUNCT][1] , \ID_EXE_i[FUNCT][0] , 
        \ID_EXE_i[SIGN_EXTEND][31] , \ID_EXE_i[SIGN_EXTEND][30] , 
        \ID_EXE_i[SIGN_EXTEND][29] , \ID_EXE_i[SIGN_EXTEND][28] , 
        \ID_EXE_i[SIGN_EXTEND][27] , \ID_EXE_i[SIGN_EXTEND][26] , 
        \ID_EXE_i[SIGN_EXTEND][25] , \ID_EXE_i[SIGN_EXTEND][24] , 
        \ID_EXE_i[SIGN_EXTEND][23] , \ID_EXE_i[SIGN_EXTEND][22] , 
        \ID_EXE_i[SIGN_EXTEND][21] , \ID_EXE_i[SIGN_EXTEND][20] , 
        \ID_EXE_i[SIGN_EXTEND][19] , \ID_EXE_i[SIGN_EXTEND][18] , 
        \ID_EXE_i[SIGN_EXTEND][17] , \ID_EXE_i[SIGN_EXTEND][16] , 
        \ID_EXE_i[SIGN_EXTEND][15] , \ID_EXE_i[SIGN_EXTEND][14] , 
        \ID_EXE_i[SIGN_EXTEND][13] , \ID_EXE_i[SIGN_EXTEND][12] , 
        \ID_EXE_i[SIGN_EXTEND][11] , \ID_EXE_i[SIGN_EXTEND][10] , 
        \ID_EXE_i[SIGN_EXTEND][9] , \ID_EXE_i[SIGN_EXTEND][8] , 
        \ID_EXE_i[SIGN_EXTEND][7] , \ID_EXE_i[SIGN_EXTEND][6] , 
        \ID_EXE_i[SIGN_EXTEND][5] , \ID_EXE_i[SIGN_EXTEND][4] , 
        \ID_EXE_i[SIGN_EXTEND][3] , \ID_EXE_i[SIGN_EXTEND][2] , 
        \ID_EXE_i[SIGN_EXTEND][1] , \ID_EXE_i[SIGN_EXTEND][0] , 
        \ID_EXE_i[PC_PLUS1][11] , \ID_EXE_i[PC_PLUS1][10] , 
        \ID_EXE_i[PC_PLUS1][9] , \ID_EXE_i[PC_PLUS1][8] , 
        \ID_EXE_i[PC_PLUS1][7] , \ID_EXE_i[PC_PLUS1][6] , 
        \ID_EXE_i[PC_PLUS1][5] , \ID_EXE_i[PC_PLUS1][4] , 
        \ID_EXE_i[PC_PLUS1][3] , \ID_EXE_i[PC_PLUS1][2] , 
        \ID_EXE_i[PC_PLUS1][1] , \ID_EXE_i[PC_PLUS1][0] , \ID_EXE_i[RS][4] , 
        \ID_EXE_i[RS][3] , \ID_EXE_i[RS][2] , \ID_EXE_i[RS][1] , 
        \ID_EXE_i[RS][0] , \ID_EXE_i[RT][4] , \ID_EXE_i[RT][3] , 
        \ID_EXE_i[RT][2] , \ID_EXE_i[RT][1] , \ID_EXE_i[RT][0] , 
        \ID_EXE_i[RD][4] , \ID_EXE_i[RD][3] , \ID_EXE_i[RD][2] , 
        \ID_EXE_i[RD][1] , \ID_EXE_i[RD][0] , \ID_EXE_i[ALUSRC_B] , 
        \ID_EXE_i[MEMTOREG] , \ID_EXE_i[REGWRITE] , \ID_EXE_i[MEMWEN_N] , 
        \ID_EXE_i[CALU_OP][3] , \ID_EXE_i[CALU_OP][2] , \ID_EXE_i[CALU_OP][1] , 
        \ID_EXE_i[CALU_OP][0] , \ID_EXE_i[REGDST] }), .ID_EXE_o({
        \ID_EXE_o[REGA][31] , \ID_EXE_o[REGA][30] , \ID_EXE_o[REGA][29] , 
        \ID_EXE_o[REGA][28] , \ID_EXE_o[REGA][27] , \ID_EXE_o[REGA][26] , 
        \ID_EXE_o[REGA][25] , \ID_EXE_o[REGA][24] , \ID_EXE_o[REGA][23] , 
        \ID_EXE_o[REGA][22] , \ID_EXE_o[REGA][21] , \ID_EXE_o[REGA][20] , 
        \ID_EXE_o[REGA][19] , \ID_EXE_o[REGA][18] , \ID_EXE_o[REGA][17] , 
        \ID_EXE_o[REGA][16] , \ID_EXE_o[REGA][15] , \ID_EXE_o[REGA][14] , 
        \ID_EXE_o[REGA][13] , \ID_EXE_o[REGA][12] , \ID_EXE_o[REGA][11] , 
        \ID_EXE_o[REGA][10] , \ID_EXE_o[REGA][9] , \ID_EXE_o[REGA][8] , 
        \ID_EXE_o[REGA][7] , \ID_EXE_o[REGA][6] , \ID_EXE_o[REGA][5] , 
        \ID_EXE_o[REGA][4] , \ID_EXE_o[REGA][3] , \ID_EXE_o[REGA][2] , 
        \ID_EXE_o[REGA][1] , \ID_EXE_o[REGA][0] , \ID_EXE_o[REGB][31] , 
        \ID_EXE_o[REGB][30] , \ID_EXE_o[REGB][29] , \ID_EXE_o[REGB][28] , 
        \ID_EXE_o[REGB][27] , \ID_EXE_o[REGB][26] , \ID_EXE_o[REGB][25] , 
        \ID_EXE_o[REGB][24] , \ID_EXE_o[REGB][23] , \ID_EXE_o[REGB][22] , 
        \ID_EXE_o[REGB][21] , \ID_EXE_o[REGB][20] , \ID_EXE_o[REGB][19] , 
        \ID_EXE_o[REGB][18] , \ID_EXE_o[REGB][17] , \ID_EXE_o[REGB][16] , 
        \ID_EXE_o[REGB][15] , \ID_EXE_o[REGB][14] , \ID_EXE_o[REGB][13] , 
        \ID_EXE_o[REGB][12] , \ID_EXE_o[REGB][11] , \ID_EXE_o[REGB][10] , 
        \ID_EXE_o[REGB][9] , \ID_EXE_o[REGB][8] , \ID_EXE_o[REGB][7] , 
        \ID_EXE_o[REGB][6] , \ID_EXE_o[REGB][5] , \ID_EXE_o[REGB][4] , 
        \ID_EXE_o[REGB][3] , \ID_EXE_o[REGB][2] , \ID_EXE_o[REGB][1] , 
        \ID_EXE_o[REGB][0] , \ID_EXE_o[SHAMT][4] , \ID_EXE_o[SHAMT][3] , 
        \ID_EXE_o[SHAMT][2] , \ID_EXE_o[SHAMT][1] , \ID_EXE_o[SHAMT][0] , 
        \ID_EXE_o[FUNCT][5] , \ID_EXE_o[FUNCT][4] , \ID_EXE_o[FUNCT][3] , 
        \ID_EXE_o[FUNCT][2] , \ID_EXE_o[FUNCT][1] , \ID_EXE_o[FUNCT][0] , 
        \ID_EXE_o[SIGN_EXTEND][31] , \ID_EXE_o[SIGN_EXTEND][30] , 
        \ID_EXE_o[SIGN_EXTEND][29] , \ID_EXE_o[SIGN_EXTEND][28] , 
        \ID_EXE_o[SIGN_EXTEND][27] , \ID_EXE_o[SIGN_EXTEND][26] , 
        \ID_EXE_o[SIGN_EXTEND][25] , \ID_EXE_o[SIGN_EXTEND][24] , 
        \ID_EXE_o[SIGN_EXTEND][23] , \ID_EXE_o[SIGN_EXTEND][22] , 
        \ID_EXE_o[SIGN_EXTEND][21] , \ID_EXE_o[SIGN_EXTEND][20] , 
        \ID_EXE_o[SIGN_EXTEND][19] , \ID_EXE_o[SIGN_EXTEND][18] , 
        \ID_EXE_o[SIGN_EXTEND][17] , \ID_EXE_o[SIGN_EXTEND][16] , 
        \ID_EXE_o[SIGN_EXTEND][15] , \ID_EXE_o[SIGN_EXTEND][14] , 
        \ID_EXE_o[SIGN_EXTEND][13] , \ID_EXE_o[SIGN_EXTEND][12] , 
        \ID_EXE_o[SIGN_EXTEND][11] , \ID_EXE_o[SIGN_EXTEND][10] , 
        \ID_EXE_o[SIGN_EXTEND][9] , \ID_EXE_o[SIGN_EXTEND][8] , 
        \ID_EXE_o[SIGN_EXTEND][7] , \ID_EXE_o[SIGN_EXTEND][6] , 
        \ID_EXE_o[SIGN_EXTEND][5] , \ID_EXE_o[SIGN_EXTEND][4] , 
        \ID_EXE_o[SIGN_EXTEND][3] , \ID_EXE_o[SIGN_EXTEND][2] , 
        \ID_EXE_o[SIGN_EXTEND][1] , \ID_EXE_o[SIGN_EXTEND][0] , 
        \ID_EXE_o[PC_PLUS1][11] , \ID_EXE_o[PC_PLUS1][10] , 
        \ID_EXE_o[PC_PLUS1][9] , \ID_EXE_o[PC_PLUS1][8] , 
        \ID_EXE_o[PC_PLUS1][7] , \ID_EXE_o[PC_PLUS1][6] , 
        \ID_EXE_o[PC_PLUS1][5] , \ID_EXE_o[PC_PLUS1][4] , 
        \ID_EXE_o[PC_PLUS1][3] , \ID_EXE_o[PC_PLUS1][2] , 
        \ID_EXE_o[PC_PLUS1][1] , \ID_EXE_o[PC_PLUS1][0] , \ID_EXE_o[RS][4] , 
        \ID_EXE_o[RS][3] , \ID_EXE_o[RS][2] , \ID_EXE_o[RS][1] , 
        \ID_EXE_o[RS][0] , \ID_EXE_o[RT][4] , \ID_EXE_o[RT][3] , 
        \ID_EXE_o[RT][2] , \ID_EXE_o[RT][1] , \ID_EXE_o[RT][0] , 
        \ID_EXE_o[RD][4] , \ID_EXE_o[RD][3] , \ID_EXE_o[RD][2] , 
        \ID_EXE_o[RD][1] , \ID_EXE_o[RD][0] , \ID_EXE_o[ALUSRC_B] , 
        \ID_EXE_o[MEMTOREG] , \ID_EXE_o[REGWRITE] , \ID_EXE_o[MEMWEN_N] , 
        \ID_EXE_o[CALU_OP][3] , \ID_EXE_o[CALU_OP][2] , \ID_EXE_o[CALU_OP][1] , 
        \ID_EXE_o[CALU_OP][0] , \ID_EXE_o[REGDST] }) );
  input clk, rst_n, halt_i, \ID_EXE_i[REGA][31] , \ID_EXE_i[REGA][30] ,
         \ID_EXE_i[REGA][29] , \ID_EXE_i[REGA][28] , \ID_EXE_i[REGA][27] ,
         \ID_EXE_i[REGA][26] , \ID_EXE_i[REGA][25] , \ID_EXE_i[REGA][24] ,
         \ID_EXE_i[REGA][23] , \ID_EXE_i[REGA][22] , \ID_EXE_i[REGA][21] ,
         \ID_EXE_i[REGA][20] , \ID_EXE_i[REGA][19] , \ID_EXE_i[REGA][18] ,
         \ID_EXE_i[REGA][17] , \ID_EXE_i[REGA][16] , \ID_EXE_i[REGA][15] ,
         \ID_EXE_i[REGA][14] , \ID_EXE_i[REGA][13] , \ID_EXE_i[REGA][12] ,
         \ID_EXE_i[REGA][11] , \ID_EXE_i[REGA][10] , \ID_EXE_i[REGA][9] ,
         \ID_EXE_i[REGA][8] , \ID_EXE_i[REGA][7] , \ID_EXE_i[REGA][6] ,
         \ID_EXE_i[REGA][5] , \ID_EXE_i[REGA][4] , \ID_EXE_i[REGA][3] ,
         \ID_EXE_i[REGA][2] , \ID_EXE_i[REGA][1] , \ID_EXE_i[REGA][0] ,
         \ID_EXE_i[REGB][31] , \ID_EXE_i[REGB][30] , \ID_EXE_i[REGB][29] ,
         \ID_EXE_i[REGB][28] , \ID_EXE_i[REGB][27] , \ID_EXE_i[REGB][26] ,
         \ID_EXE_i[REGB][25] , \ID_EXE_i[REGB][24] , \ID_EXE_i[REGB][23] ,
         \ID_EXE_i[REGB][22] , \ID_EXE_i[REGB][21] , \ID_EXE_i[REGB][20] ,
         \ID_EXE_i[REGB][19] , \ID_EXE_i[REGB][18] , \ID_EXE_i[REGB][17] ,
         \ID_EXE_i[REGB][16] , \ID_EXE_i[REGB][15] , \ID_EXE_i[REGB][14] ,
         \ID_EXE_i[REGB][13] , \ID_EXE_i[REGB][12] , \ID_EXE_i[REGB][11] ,
         \ID_EXE_i[REGB][10] , \ID_EXE_i[REGB][9] , \ID_EXE_i[REGB][8] ,
         \ID_EXE_i[REGB][7] , \ID_EXE_i[REGB][6] , \ID_EXE_i[REGB][5] ,
         \ID_EXE_i[REGB][4] , \ID_EXE_i[REGB][3] , \ID_EXE_i[REGB][2] ,
         \ID_EXE_i[REGB][1] , \ID_EXE_i[REGB][0] , \ID_EXE_i[SHAMT][4] ,
         \ID_EXE_i[SHAMT][3] , \ID_EXE_i[SHAMT][2] , \ID_EXE_i[SHAMT][1] ,
         \ID_EXE_i[SHAMT][0] , \ID_EXE_i[FUNCT][5] , \ID_EXE_i[FUNCT][4] ,
         \ID_EXE_i[FUNCT][3] , \ID_EXE_i[FUNCT][2] , \ID_EXE_i[FUNCT][1] ,
         \ID_EXE_i[FUNCT][0] , \ID_EXE_i[SIGN_EXTEND][31] ,
         \ID_EXE_i[SIGN_EXTEND][30] , \ID_EXE_i[SIGN_EXTEND][29] ,
         \ID_EXE_i[SIGN_EXTEND][28] , \ID_EXE_i[SIGN_EXTEND][27] ,
         \ID_EXE_i[SIGN_EXTEND][26] , \ID_EXE_i[SIGN_EXTEND][25] ,
         \ID_EXE_i[SIGN_EXTEND][24] , \ID_EXE_i[SIGN_EXTEND][23] ,
         \ID_EXE_i[SIGN_EXTEND][22] , \ID_EXE_i[SIGN_EXTEND][21] ,
         \ID_EXE_i[SIGN_EXTEND][20] , \ID_EXE_i[SIGN_EXTEND][19] ,
         \ID_EXE_i[SIGN_EXTEND][18] , \ID_EXE_i[SIGN_EXTEND][17] ,
         \ID_EXE_i[SIGN_EXTEND][16] , \ID_EXE_i[SIGN_EXTEND][15] ,
         \ID_EXE_i[SIGN_EXTEND][14] , \ID_EXE_i[SIGN_EXTEND][13] ,
         \ID_EXE_i[SIGN_EXTEND][12] , \ID_EXE_i[SIGN_EXTEND][11] ,
         \ID_EXE_i[SIGN_EXTEND][10] , \ID_EXE_i[SIGN_EXTEND][9] ,
         \ID_EXE_i[SIGN_EXTEND][8] , \ID_EXE_i[SIGN_EXTEND][7] ,
         \ID_EXE_i[SIGN_EXTEND][6] , \ID_EXE_i[SIGN_EXTEND][5] ,
         \ID_EXE_i[SIGN_EXTEND][4] , \ID_EXE_i[SIGN_EXTEND][3] ,
         \ID_EXE_i[SIGN_EXTEND][2] , \ID_EXE_i[SIGN_EXTEND][1] ,
         \ID_EXE_i[SIGN_EXTEND][0] , \ID_EXE_i[PC_PLUS1][11] ,
         \ID_EXE_i[PC_PLUS1][10] , \ID_EXE_i[PC_PLUS1][9] ,
         \ID_EXE_i[PC_PLUS1][8] , \ID_EXE_i[PC_PLUS1][7] ,
         \ID_EXE_i[PC_PLUS1][6] , \ID_EXE_i[PC_PLUS1][5] ,
         \ID_EXE_i[PC_PLUS1][4] , \ID_EXE_i[PC_PLUS1][3] ,
         \ID_EXE_i[PC_PLUS1][2] , \ID_EXE_i[PC_PLUS1][1] ,
         \ID_EXE_i[PC_PLUS1][0] , \ID_EXE_i[RS][4] , \ID_EXE_i[RS][3] ,
         \ID_EXE_i[RS][2] , \ID_EXE_i[RS][1] , \ID_EXE_i[RS][0] ,
         \ID_EXE_i[RT][4] , \ID_EXE_i[RT][3] , \ID_EXE_i[RT][2] ,
         \ID_EXE_i[RT][1] , \ID_EXE_i[RT][0] , \ID_EXE_i[RD][4] ,
         \ID_EXE_i[RD][3] , \ID_EXE_i[RD][2] , \ID_EXE_i[RD][1] ,
         \ID_EXE_i[RD][0] , \ID_EXE_i[ALUSRC_B] , \ID_EXE_i[MEMTOREG] ,
         \ID_EXE_i[REGWRITE] , \ID_EXE_i[MEMWEN_N] , \ID_EXE_i[CALU_OP][3] ,
         \ID_EXE_i[CALU_OP][2] , \ID_EXE_i[CALU_OP][1] ,
         \ID_EXE_i[CALU_OP][0] , \ID_EXE_i[REGDST] ;
  output \ID_EXE_o[REGA][31] , \ID_EXE_o[REGA][30] , \ID_EXE_o[REGA][29] ,
         \ID_EXE_o[REGA][28] , \ID_EXE_o[REGA][27] , \ID_EXE_o[REGA][26] ,
         \ID_EXE_o[REGA][25] , \ID_EXE_o[REGA][24] , \ID_EXE_o[REGA][23] ,
         \ID_EXE_o[REGA][22] , \ID_EXE_o[REGA][21] , \ID_EXE_o[REGA][20] ,
         \ID_EXE_o[REGA][19] , \ID_EXE_o[REGA][18] , \ID_EXE_o[REGA][17] ,
         \ID_EXE_o[REGA][16] , \ID_EXE_o[REGA][15] , \ID_EXE_o[REGA][14] ,
         \ID_EXE_o[REGA][13] , \ID_EXE_o[REGA][12] , \ID_EXE_o[REGA][11] ,
         \ID_EXE_o[REGA][10] , \ID_EXE_o[REGA][9] , \ID_EXE_o[REGA][8] ,
         \ID_EXE_o[REGA][7] , \ID_EXE_o[REGA][6] , \ID_EXE_o[REGA][5] ,
         \ID_EXE_o[REGA][4] , \ID_EXE_o[REGA][3] , \ID_EXE_o[REGA][2] ,
         \ID_EXE_o[REGA][1] , \ID_EXE_o[REGA][0] , \ID_EXE_o[REGB][31] ,
         \ID_EXE_o[REGB][30] , \ID_EXE_o[REGB][29] , \ID_EXE_o[REGB][28] ,
         \ID_EXE_o[REGB][27] , \ID_EXE_o[REGB][26] , \ID_EXE_o[REGB][25] ,
         \ID_EXE_o[REGB][24] , \ID_EXE_o[REGB][23] , \ID_EXE_o[REGB][22] ,
         \ID_EXE_o[REGB][21] , \ID_EXE_o[REGB][20] , \ID_EXE_o[REGB][19] ,
         \ID_EXE_o[REGB][18] , \ID_EXE_o[REGB][17] , \ID_EXE_o[REGB][16] ,
         \ID_EXE_o[REGB][15] , \ID_EXE_o[REGB][14] , \ID_EXE_o[REGB][13] ,
         \ID_EXE_o[REGB][12] , \ID_EXE_o[REGB][11] , \ID_EXE_o[REGB][10] ,
         \ID_EXE_o[REGB][9] , \ID_EXE_o[REGB][8] , \ID_EXE_o[REGB][7] ,
         \ID_EXE_o[REGB][6] , \ID_EXE_o[REGB][5] , \ID_EXE_o[REGB][4] ,
         \ID_EXE_o[REGB][3] , \ID_EXE_o[REGB][2] , \ID_EXE_o[REGB][1] ,
         \ID_EXE_o[REGB][0] , \ID_EXE_o[SHAMT][4] , \ID_EXE_o[SHAMT][3] ,
         \ID_EXE_o[SHAMT][2] , \ID_EXE_o[SHAMT][1] , \ID_EXE_o[SHAMT][0] ,
         \ID_EXE_o[FUNCT][5] , \ID_EXE_o[FUNCT][4] , \ID_EXE_o[FUNCT][3] ,
         \ID_EXE_o[FUNCT][2] , \ID_EXE_o[FUNCT][1] , \ID_EXE_o[FUNCT][0] ,
         \ID_EXE_o[SIGN_EXTEND][31] , \ID_EXE_o[SIGN_EXTEND][30] ,
         \ID_EXE_o[SIGN_EXTEND][29] , \ID_EXE_o[SIGN_EXTEND][28] ,
         \ID_EXE_o[SIGN_EXTEND][27] , \ID_EXE_o[SIGN_EXTEND][26] ,
         \ID_EXE_o[SIGN_EXTEND][25] , \ID_EXE_o[SIGN_EXTEND][24] ,
         \ID_EXE_o[SIGN_EXTEND][23] , \ID_EXE_o[SIGN_EXTEND][22] ,
         \ID_EXE_o[SIGN_EXTEND][21] , \ID_EXE_o[SIGN_EXTEND][20] ,
         \ID_EXE_o[SIGN_EXTEND][19] , \ID_EXE_o[SIGN_EXTEND][18] ,
         \ID_EXE_o[SIGN_EXTEND][17] , \ID_EXE_o[SIGN_EXTEND][16] ,
         \ID_EXE_o[SIGN_EXTEND][15] , \ID_EXE_o[SIGN_EXTEND][14] ,
         \ID_EXE_o[SIGN_EXTEND][13] , \ID_EXE_o[SIGN_EXTEND][12] ,
         \ID_EXE_o[SIGN_EXTEND][11] , \ID_EXE_o[SIGN_EXTEND][10] ,
         \ID_EXE_o[SIGN_EXTEND][9] , \ID_EXE_o[SIGN_EXTEND][8] ,
         \ID_EXE_o[SIGN_EXTEND][7] , \ID_EXE_o[SIGN_EXTEND][6] ,
         \ID_EXE_o[SIGN_EXTEND][5] , \ID_EXE_o[SIGN_EXTEND][4] ,
         \ID_EXE_o[SIGN_EXTEND][3] , \ID_EXE_o[SIGN_EXTEND][2] ,
         \ID_EXE_o[SIGN_EXTEND][1] , \ID_EXE_o[SIGN_EXTEND][0] ,
         \ID_EXE_o[PC_PLUS1][11] , \ID_EXE_o[PC_PLUS1][10] ,
         \ID_EXE_o[PC_PLUS1][9] , \ID_EXE_o[PC_PLUS1][8] ,
         \ID_EXE_o[PC_PLUS1][7] , \ID_EXE_o[PC_PLUS1][6] ,
         \ID_EXE_o[PC_PLUS1][5] , \ID_EXE_o[PC_PLUS1][4] ,
         \ID_EXE_o[PC_PLUS1][3] , \ID_EXE_o[PC_PLUS1][2] ,
         \ID_EXE_o[PC_PLUS1][1] , \ID_EXE_o[PC_PLUS1][0] , \ID_EXE_o[RS][4] ,
         \ID_EXE_o[RS][3] , \ID_EXE_o[RS][2] , \ID_EXE_o[RS][1] ,
         \ID_EXE_o[RS][0] , \ID_EXE_o[RT][4] , \ID_EXE_o[RT][3] ,
         \ID_EXE_o[RT][2] , \ID_EXE_o[RT][1] , \ID_EXE_o[RT][0] ,
         \ID_EXE_o[RD][4] , \ID_EXE_o[RD][3] , \ID_EXE_o[RD][2] ,
         \ID_EXE_o[RD][1] , \ID_EXE_o[RD][0] , \ID_EXE_o[ALUSRC_B] ,
         \ID_EXE_o[MEMTOREG] , \ID_EXE_o[REGWRITE] , \ID_EXE_o[MEMWEN_N] ,
         \ID_EXE_o[CALU_OP][3] , \ID_EXE_o[CALU_OP][2] ,
         \ID_EXE_o[CALU_OP][1] , \ID_EXE_o[CALU_OP][0] , \ID_EXE_o[REGDST] ;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n1,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180;

  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][31]  ( .D(n144), .CP(clk), .RN(n164), 
        .Q(\ID_EXE_o[REGA][31] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][30]  ( .D(n143), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][30] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][29]  ( .D(n142), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][29] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][28]  ( .D(n141), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][28] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][27]  ( .D(n140), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][27] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][26]  ( .D(n139), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][26] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][25]  ( .D(n138), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][25] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][24]  ( .D(n137), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][24] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][23]  ( .D(n136), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][23] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][22]  ( .D(n135), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][22] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][21]  ( .D(n134), .CP(clk), .RN(n175), 
        .Q(\ID_EXE_o[REGA][21] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][20]  ( .D(n133), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][20] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][19]  ( .D(n132), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][19] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][18]  ( .D(n131), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][18] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][17]  ( .D(n130), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][17] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][16]  ( .D(n129), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][16] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][15]  ( .D(n128), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][15] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][14]  ( .D(n127), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][14] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][13]  ( .D(n126), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][13] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][12]  ( .D(n125), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][12] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][11]  ( .D(n124), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][11] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][10]  ( .D(n123), .CP(clk), .RN(n174), 
        .Q(\ID_EXE_o[REGA][10] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][9]  ( .D(n122), .CP(clk), .RN(n174), .Q(
        \ID_EXE_o[REGA][9] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][8]  ( .D(n121), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][8] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][7]  ( .D(n120), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][7] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][6]  ( .D(n119), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][6] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][5]  ( .D(n118), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][5] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][4]  ( .D(n117), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][3]  ( .D(n116), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][2]  ( .D(n115), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][1]  ( .D(n114), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGA][0]  ( .D(n113), .CP(clk), .RN(n173), .Q(
        \ID_EXE_o[REGA][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][31]  ( .D(n112), .CP(clk), .RN(n173), 
        .Q(\ID_EXE_o[REGB][31] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][30]  ( .D(n111), .CP(clk), .RN(n173), 
        .Q(\ID_EXE_o[REGB][30] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][29]  ( .D(n110), .CP(clk), .RN(n173), 
        .Q(\ID_EXE_o[REGB][29] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][28]  ( .D(n109), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][28] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][27]  ( .D(n108), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][27] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][26]  ( .D(n107), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][26] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][25]  ( .D(n106), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][25] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][24]  ( .D(n105), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][24] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][23]  ( .D(n104), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][23] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][22]  ( .D(n103), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][22] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][21]  ( .D(n102), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][21] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][20]  ( .D(n101), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][20] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][19]  ( .D(n100), .CP(clk), .RN(n172), 
        .Q(\ID_EXE_o[REGB][19] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][18]  ( .D(n99), .CP(clk), .RN(n172), .Q(
        \ID_EXE_o[REGB][18] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][17]  ( .D(n98), .CP(clk), .RN(n172), .Q(
        \ID_EXE_o[REGB][17] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][16]  ( .D(n97), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][16] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][15]  ( .D(n96), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][15] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][14]  ( .D(n95), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][14] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][13]  ( .D(n94), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][13] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][12]  ( .D(n93), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][12] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][11]  ( .D(n92), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][11] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][10]  ( .D(n91), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][10] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][9]  ( .D(n90), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][9] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][8]  ( .D(n89), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][8] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][7]  ( .D(n88), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][7] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][6]  ( .D(n87), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][6] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][5]  ( .D(n86), .CP(clk), .RN(n171), .Q(
        \ID_EXE_o[REGB][5] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][4]  ( .D(n85), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[REGB][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][3]  ( .D(n84), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[REGB][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][2]  ( .D(n83), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[REGB][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][1]  ( .D(n82), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[REGB][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGB][0]  ( .D(n81), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[REGB][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SHAMT][4]  ( .D(n80), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[SHAMT][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SHAMT][3]  ( .D(n79), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[SHAMT][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SHAMT][2]  ( .D(n78), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[SHAMT][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SHAMT][1]  ( .D(n77), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[SHAMT][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SHAMT][0]  ( .D(n76), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[SHAMT][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][5]  ( .D(n75), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[FUNCT][5] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][4]  ( .D(n74), .CP(clk), .RN(n170), .Q(
        \ID_EXE_o[FUNCT][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][3]  ( .D(n73), .CP(clk), .RN(n169), .Q(
        \ID_EXE_o[FUNCT][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][2]  ( .D(n72), .CP(clk), .RN(n169), .Q(
        \ID_EXE_o[FUNCT][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][1]  ( .D(n71), .CP(clk), .RN(n169), .Q(
        \ID_EXE_o[FUNCT][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[FUNCT][0]  ( .D(n70), .CP(clk), .RN(n169), .Q(
        \ID_EXE_o[FUNCT][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][31]  ( .D(n69), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][31] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][30]  ( .D(n68), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][30] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][29]  ( .D(n67), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][29] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][28]  ( .D(n66), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][28] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][27]  ( .D(n65), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][27] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][26]  ( .D(n64), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][26] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][25]  ( .D(n63), .CP(clk), .RN(
        n169), .Q(\ID_EXE_o[SIGN_EXTEND][25] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][24]  ( .D(n62), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][24] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][23]  ( .D(n61), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][23] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][22]  ( .D(n60), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][22] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][21]  ( .D(n59), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][21] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][20]  ( .D(n58), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][20] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][19]  ( .D(n57), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][19] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][18]  ( .D(n56), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][18] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][17]  ( .D(n55), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][17] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][16]  ( .D(n54), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][16] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][15]  ( .D(n53), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][15] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][14]  ( .D(n52), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][14] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][13]  ( .D(n51), .CP(clk), .RN(
        n168), .Q(\ID_EXE_o[SIGN_EXTEND][13] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][12]  ( .D(n50), .CP(clk), .RN(
        n167), .Q(\ID_EXE_o[SIGN_EXTEND][12] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][11]  ( .D(n49), .CP(clk), .RN(
        n167), .Q(\ID_EXE_o[SIGN_EXTEND][11] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][10]  ( .D(n48), .CP(clk), .RN(
        n167), .Q(\ID_EXE_o[SIGN_EXTEND][10] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][9]  ( .D(n47), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][9] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][8]  ( .D(n46), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][8] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][7]  ( .D(n45), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][7] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][6]  ( .D(n44), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][6] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][5]  ( .D(n43), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][5] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][4]  ( .D(n42), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][3]  ( .D(n41), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][2]  ( .D(n40), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][1]  ( .D(n39), .CP(clk), .RN(n167), .Q(\ID_EXE_o[SIGN_EXTEND][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[SIGN_EXTEND][0]  ( .D(n38), .CP(clk), .RN(n166), .Q(\ID_EXE_o[SIGN_EXTEND][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][11]  ( .D(n37), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][11] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][10]  ( .D(n36), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][10] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][9]  ( .D(n35), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][9] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][8]  ( .D(n34), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][8] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][7]  ( .D(n33), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][7] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][6]  ( .D(n32), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][6] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][5]  ( .D(n31), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][5] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][4]  ( .D(n30), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][3]  ( .D(n29), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][2]  ( .D(n28), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][1]  ( .D(n27), .CP(clk), .RN(n166), 
        .Q(\ID_EXE_o[PC_PLUS1][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[PC_PLUS1][0]  ( .D(n26), .CP(clk), .RN(n165), 
        .Q(\ID_EXE_o[PC_PLUS1][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RS][4]  ( .D(n25), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RS][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RS][3]  ( .D(n24), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RS][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RS][2]  ( .D(n23), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RS][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RS][1]  ( .D(n22), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RS][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RS][0]  ( .D(n21), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RS][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RT][4]  ( .D(n20), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RT][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RT][3]  ( .D(n19), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RT][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RT][2]  ( .D(n18), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RT][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RT][1]  ( .D(n17), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RT][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RT][0]  ( .D(n16), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RT][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RD][4]  ( .D(n15), .CP(clk), .RN(n165), .Q(
        \ID_EXE_o[RD][4] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RD][3]  ( .D(n14), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[RD][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RD][2]  ( .D(n13), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[RD][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RD][1]  ( .D(n12), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[RD][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[RD][0]  ( .D(n11), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[RD][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[ALUSRC_B]  ( .D(n10), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[ALUSRC_B] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[MEMTOREG]  ( .D(n9), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[MEMTOREG] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGWRITE]  ( .D(n8), .CP(clk), .RN(n164), .Q(
        \ID_EXE_o[REGWRITE] ) );
  HS65_LH_DFPSQX9 \id_exe_c_reg[MEMWEN_N]  ( .D(n7), .CP(clk), .SN(n175), .Q(
        \ID_EXE_o[MEMWEN_N] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[CALU_OP][3]  ( .D(n6), .CP(clk), .RN(n164), 
        .Q(\ID_EXE_o[CALU_OP][3] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[CALU_OP][2]  ( .D(n5), .CP(clk), .RN(n164), 
        .Q(\ID_EXE_o[CALU_OP][2] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[CALU_OP][1]  ( .D(n4), .CP(clk), .RN(n164), 
        .Q(\ID_EXE_o[CALU_OP][1] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[CALU_OP][0]  ( .D(n3), .CP(clk), .RN(n164), 
        .Q(\ID_EXE_o[CALU_OP][0] ) );
  HS65_LH_DFPRQX9 \id_exe_c_reg[REGDST]  ( .D(n2), .CP(clk), .RN(n169), .Q(
        \ID_EXE_o[REGDST] ) );
  HS65_LH_BFX9 U2 ( .A(n179), .Z(n165) );
  HS65_LH_BFX9 U3 ( .A(n179), .Z(n166) );
  HS65_LH_BFX9 U4 ( .A(n178), .Z(n167) );
  HS65_LH_BFX9 U5 ( .A(n178), .Z(n168) );
  HS65_LH_BFX9 U6 ( .A(n178), .Z(n169) );
  HS65_LH_BFX9 U7 ( .A(n177), .Z(n170) );
  HS65_LH_BFX9 U8 ( .A(n177), .Z(n171) );
  HS65_LH_BFX9 U9 ( .A(n177), .Z(n172) );
  HS65_LH_BFX9 U10 ( .A(n176), .Z(n173) );
  HS65_LH_BFX9 U11 ( .A(n176), .Z(n174) );
  HS65_LH_BFX9 U12 ( .A(n179), .Z(n164) );
  HS65_LH_BFX9 U13 ( .A(n176), .Z(n175) );
  HS65_LH_BFX9 U14 ( .A(n163), .Z(n178) );
  HS65_LH_BFX9 U15 ( .A(n162), .Z(n177) );
  HS65_LH_BFX9 U16 ( .A(n162), .Z(n176) );
  HS65_LH_BFX9 U17 ( .A(n163), .Z(n179) );
  HS65_LH_BFX9 U18 ( .A(n1), .Z(n150) );
  HS65_LH_BFX9 U19 ( .A(n1), .Z(n151) );
  HS65_LH_BFX9 U20 ( .A(n1), .Z(n152) );
  HS65_LH_BFX9 U21 ( .A(n145), .Z(n153) );
  HS65_LH_BFX9 U22 ( .A(n145), .Z(n154) );
  HS65_LH_BFX9 U23 ( .A(n145), .Z(n155) );
  HS65_LH_BFX9 U24 ( .A(n146), .Z(n156) );
  HS65_LH_BFX9 U25 ( .A(n146), .Z(n157) );
  HS65_LH_BFX9 U26 ( .A(n146), .Z(n158) );
  HS65_LH_BFX9 U27 ( .A(n147), .Z(n159) );
  HS65_LH_BFX9 U28 ( .A(n147), .Z(n160) );
  HS65_LH_BFX9 U29 ( .A(n147), .Z(n161) );
  HS65_LH_BFX9 U30 ( .A(rst_n), .Z(n162) );
  HS65_LH_BFX9 U31 ( .A(rst_n), .Z(n163) );
  HS65_LH_BFX9 U32 ( .A(n149), .Z(n1) );
  HS65_LH_BFX9 U33 ( .A(n149), .Z(n145) );
  HS65_LH_BFX9 U34 ( .A(n148), .Z(n146) );
  HS65_LH_BFX9 U35 ( .A(n148), .Z(n147) );
  HS65_LH_BFX9 U36 ( .A(n180), .Z(n149) );
  HS65_LH_BFX9 U37 ( .A(n180), .Z(n148) );
  HS65_LH_AO22X9 U38 ( .A(\ID_EXE_o[REGA][0] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][0] ), .D(n159), .Z(n113) );
  HS65_LH_AO22X9 U39 ( .A(\ID_EXE_o[REGA][1] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][1] ), .D(n159), .Z(n114) );
  HS65_LH_AO22X9 U40 ( .A(\ID_EXE_o[REGA][2] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][2] ), .D(n159), .Z(n115) );
  HS65_LH_AO22X9 U41 ( .A(\ID_EXE_o[REGA][3] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][3] ), .D(n159), .Z(n116) );
  HS65_LH_AO22X9 U42 ( .A(\ID_EXE_o[REGA][4] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][4] ), .D(n159), .Z(n117) );
  HS65_LH_AO22X9 U43 ( .A(\ID_EXE_o[REGA][5] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][5] ), .D(n159), .Z(n118) );
  HS65_LH_AO22X9 U44 ( .A(\ID_EXE_o[REGA][6] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][6] ), .D(n159), .Z(n119) );
  HS65_LH_AO22X9 U45 ( .A(\ID_EXE_o[REGA][7] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][7] ), .D(n159), .Z(n120) );
  HS65_LH_AO22X9 U46 ( .A(\ID_EXE_o[REGA][8] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][8] ), .D(n159), .Z(n121) );
  HS65_LH_AO22X9 U47 ( .A(\ID_EXE_o[REGA][9] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][9] ), .D(n160), .Z(n122) );
  HS65_LH_AO22X9 U48 ( .A(\ID_EXE_o[REGA][10] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][10] ), .D(n160), .Z(n123) );
  HS65_LH_AO22X9 U49 ( .A(\ID_EXE_o[REGA][11] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][11] ), .D(n160), .Z(n124) );
  HS65_LH_AO22X9 U50 ( .A(\ID_EXE_o[REGA][12] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][12] ), .D(n160), .Z(n125) );
  HS65_LH_AO22X9 U51 ( .A(\ID_EXE_o[REGA][13] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][13] ), .D(n160), .Z(n126) );
  HS65_LH_AO22X9 U52 ( .A(\ID_EXE_o[REGA][14] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][14] ), .D(n160), .Z(n127) );
  HS65_LH_AO22X9 U53 ( .A(\ID_EXE_o[REGA][15] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][15] ), .D(n160), .Z(n128) );
  HS65_LH_AO22X9 U54 ( .A(\ID_EXE_o[REGA][16] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][16] ), .D(n160), .Z(n129) );
  HS65_LH_AO22X9 U55 ( .A(\ID_EXE_o[REGA][17] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][17] ), .D(n160), .Z(n130) );
  HS65_LH_AO22X9 U56 ( .A(\ID_EXE_o[REGA][18] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][18] ), .D(n160), .Z(n131) );
  HS65_LH_AO22X9 U57 ( .A(\ID_EXE_o[REGA][19] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][19] ), .D(n160), .Z(n132) );
  HS65_LH_AO22X9 U58 ( .A(\ID_EXE_o[REGA][20] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][20] ), .D(n160), .Z(n133) );
  HS65_LH_AO22X9 U59 ( .A(\ID_EXE_o[REGA][21] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][21] ), .D(n161), .Z(n134) );
  HS65_LH_AO22X9 U60 ( .A(\ID_EXE_o[REGA][22] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][22] ), .D(n161), .Z(n135) );
  HS65_LH_AO22X9 U61 ( .A(\ID_EXE_o[REGA][23] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][23] ), .D(n161), .Z(n136) );
  HS65_LH_AO22X9 U62 ( .A(\ID_EXE_o[REGA][24] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][24] ), .D(n161), .Z(n137) );
  HS65_LH_AO22X9 U63 ( .A(\ID_EXE_o[REGA][25] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][25] ), .D(n161), .Z(n138) );
  HS65_LH_AO22X9 U64 ( .A(\ID_EXE_o[REGA][26] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][26] ), .D(n161), .Z(n139) );
  HS65_LH_AO22X9 U65 ( .A(\ID_EXE_o[REGA][27] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][27] ), .D(n161), .Z(n140) );
  HS65_LH_AO22X9 U66 ( .A(\ID_EXE_o[REGA][28] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][28] ), .D(n161), .Z(n141) );
  HS65_LH_AO22X9 U67 ( .A(\ID_EXE_o[REGA][29] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][29] ), .D(n161), .Z(n142) );
  HS65_LH_AO22X9 U68 ( .A(\ID_EXE_o[REGA][30] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][30] ), .D(n161), .Z(n143) );
  HS65_LH_AO22X9 U69 ( .A(\ID_EXE_o[REGA][31] ), .B(halt_i), .C(
        \ID_EXE_i[REGA][31] ), .D(n161), .Z(n144) );
  HS65_LH_AO22X9 U70 ( .A(\ID_EXE_o[REGB][0] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][0] ), .D(n156), .Z(n81) );
  HS65_LH_AO22X9 U71 ( .A(\ID_EXE_o[REGB][1] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][1] ), .D(n156), .Z(n82) );
  HS65_LH_AO22X9 U72 ( .A(\ID_EXE_o[REGB][2] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][2] ), .D(n156), .Z(n83) );
  HS65_LH_AO22X9 U73 ( .A(\ID_EXE_o[REGB][3] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][3] ), .D(n156), .Z(n84) );
  HS65_LH_AO22X9 U74 ( .A(\ID_EXE_o[REGB][4] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][4] ), .D(n156), .Z(n85) );
  HS65_LH_AO22X9 U75 ( .A(\ID_EXE_o[REGB][5] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][5] ), .D(n157), .Z(n86) );
  HS65_LH_AO22X9 U76 ( .A(\ID_EXE_o[REGB][6] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][6] ), .D(n157), .Z(n87) );
  HS65_LH_AO22X9 U77 ( .A(\ID_EXE_o[REGB][7] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][7] ), .D(n157), .Z(n88) );
  HS65_LH_AO22X9 U78 ( .A(\ID_EXE_o[REGB][8] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][8] ), .D(n157), .Z(n89) );
  HS65_LH_AO22X9 U79 ( .A(\ID_EXE_o[REGB][9] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][9] ), .D(n157), .Z(n90) );
  HS65_LH_AO22X9 U80 ( .A(\ID_EXE_o[REGB][11] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][11] ), .D(n157), .Z(n92) );
  HS65_LH_AO22X9 U81 ( .A(\ID_EXE_o[REGB][12] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][12] ), .D(n157), .Z(n93) );
  HS65_LH_AO22X9 U82 ( .A(\ID_EXE_o[REGB][13] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][13] ), .D(n157), .Z(n94) );
  HS65_LH_AO22X9 U83 ( .A(\ID_EXE_o[REGB][14] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][14] ), .D(n157), .Z(n95) );
  HS65_LH_AO22X9 U84 ( .A(\ID_EXE_o[REGB][15] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][15] ), .D(n157), .Z(n96) );
  HS65_LH_AO22X9 U85 ( .A(\ID_EXE_o[REGB][16] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][16] ), .D(n157), .Z(n97) );
  HS65_LH_AO22X9 U86 ( .A(\ID_EXE_o[REGB][17] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][17] ), .D(n158), .Z(n98) );
  HS65_LH_AO22X9 U87 ( .A(\ID_EXE_o[REGB][18] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][18] ), .D(n158), .Z(n99) );
  HS65_LH_AO22X9 U88 ( .A(\ID_EXE_o[REGB][19] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][19] ), .D(n158), .Z(n100) );
  HS65_LH_AO22X9 U89 ( .A(\ID_EXE_o[REGB][20] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][20] ), .D(n158), .Z(n101) );
  HS65_LH_AO22X9 U90 ( .A(\ID_EXE_o[REGB][21] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][21] ), .D(n158), .Z(n102) );
  HS65_LH_AO22X9 U91 ( .A(\ID_EXE_o[REGB][22] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][22] ), .D(n158), .Z(n103) );
  HS65_LH_AO22X9 U92 ( .A(\ID_EXE_o[REGB][23] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][23] ), .D(n158), .Z(n104) );
  HS65_LH_AO22X9 U93 ( .A(\ID_EXE_o[REGB][24] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][24] ), .D(n158), .Z(n105) );
  HS65_LH_AO22X9 U94 ( .A(\ID_EXE_o[REGB][25] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][25] ), .D(n158), .Z(n106) );
  HS65_LH_AO22X9 U95 ( .A(\ID_EXE_o[REGB][26] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][26] ), .D(n158), .Z(n107) );
  HS65_LH_AO22X9 U96 ( .A(\ID_EXE_o[REGB][27] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][27] ), .D(n158), .Z(n108) );
  HS65_LH_AO22X9 U97 ( .A(\ID_EXE_o[REGB][28] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][28] ), .D(n158), .Z(n109) );
  HS65_LH_AO22X9 U98 ( .A(\ID_EXE_o[REGB][29] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][29] ), .D(n159), .Z(n110) );
  HS65_LH_AO22X9 U99 ( .A(\ID_EXE_o[REGB][30] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][30] ), .D(n159), .Z(n111) );
  HS65_LH_AO22X9 U100 ( .A(\ID_EXE_o[REGB][31] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][31] ), .D(n159), .Z(n112) );
  HS65_LH_AO22X9 U101 ( .A(\ID_EXE_o[REGB][10] ), .B(halt_i), .C(
        \ID_EXE_i[REGB][10] ), .D(n157), .Z(n91) );
  HS65_LH_AO22X9 U102 ( .A(\ID_EXE_o[ALUSRC_B] ), .B(halt_i), .C(
        \ID_EXE_i[ALUSRC_B] ), .D(n150), .Z(n10) );
  HS65_LH_AO22X9 U103 ( .A(\ID_EXE_o[CALU_OP][0] ), .B(halt_i), .C(
        \ID_EXE_i[CALU_OP][0] ), .D(n150), .Z(n3) );
  HS65_LH_AO22X9 U104 ( .A(\ID_EXE_o[CALU_OP][2] ), .B(halt_i), .C(
        \ID_EXE_i[CALU_OP][2] ), .D(n150), .Z(n5) );
  HS65_LH_AO22X9 U105 ( .A(\ID_EXE_o[RT][0] ), .B(halt_i), .C(
        \ID_EXE_i[RT][0] ), .D(n151), .Z(n16) );
  HS65_LH_AO22X9 U106 ( .A(\ID_EXE_o[RS][0] ), .B(halt_i), .C(
        \ID_EXE_i[RS][0] ), .D(n151), .Z(n21) );
  HS65_LH_AO22X9 U107 ( .A(\ID_EXE_o[RT][1] ), .B(halt_i), .C(
        \ID_EXE_i[RT][1] ), .D(n151), .Z(n17) );
  HS65_LH_AO22X9 U108 ( .A(\ID_EXE_o[RT][2] ), .B(halt_i), .C(
        \ID_EXE_i[RT][2] ), .D(n151), .Z(n18) );
  HS65_LH_AO22X9 U109 ( .A(\ID_EXE_o[RT][3] ), .B(halt_i), .C(
        \ID_EXE_i[RT][3] ), .D(n151), .Z(n19) );
  HS65_LH_AO22X9 U110 ( .A(\ID_EXE_o[RS][1] ), .B(halt_i), .C(
        \ID_EXE_i[RS][1] ), .D(n151), .Z(n22) );
  HS65_LH_AO22X9 U111 ( .A(\ID_EXE_o[RS][2] ), .B(halt_i), .C(
        \ID_EXE_i[RS][2] ), .D(n151), .Z(n23) );
  HS65_LH_AO22X9 U112 ( .A(\ID_EXE_o[RS][3] ), .B(halt_i), .C(
        \ID_EXE_i[RS][3] ), .D(n151), .Z(n24) );
  HS65_LH_AO22X9 U113 ( .A(\ID_EXE_o[REGWRITE] ), .B(halt_i), .C(
        \ID_EXE_i[REGWRITE] ), .D(n150), .Z(n8) );
  HS65_LH_AO22X9 U114 ( .A(\ID_EXE_o[RT][4] ), .B(halt_i), .C(
        \ID_EXE_i[RT][4] ), .D(n151), .Z(n20) );
  HS65_LH_AO22X9 U115 ( .A(\ID_EXE_o[RS][4] ), .B(halt_i), .C(
        \ID_EXE_i[RS][4] ), .D(n151), .Z(n25) );
  HS65_LH_AO22X9 U116 ( .A(\ID_EXE_o[MEMWEN_N] ), .B(halt_i), .C(
        \ID_EXE_i[MEMWEN_N] ), .D(n150), .Z(n7) );
  HS65_LH_AO22X9 U117 ( .A(\ID_EXE_o[CALU_OP][1] ), .B(halt_i), .C(
        \ID_EXE_i[CALU_OP][1] ), .D(n150), .Z(n4) );
  HS65_LH_AO22X9 U118 ( .A(halt_i), .B(\ID_EXE_o[REGDST] ), .C(
        \ID_EXE_i[REGDST] ), .D(n150), .Z(n2) );
  HS65_LH_AO22X9 U119 ( .A(\ID_EXE_o[RD][4] ), .B(halt_i), .C(
        \ID_EXE_i[RD][4] ), .D(n151), .Z(n15) );
  HS65_LH_AO22X9 U120 ( .A(\ID_EXE_o[SIGN_EXTEND][15] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][15] ), .D(n154), .Z(n53) );
  HS65_LH_AO22X9 U121 ( .A(\ID_EXE_o[SIGN_EXTEND][16] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][16] ), .D(n154), .Z(n54) );
  HS65_LH_AO22X9 U122 ( .A(\ID_EXE_o[SIGN_EXTEND][17] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][17] ), .D(n154), .Z(n55) );
  HS65_LH_AO22X9 U123 ( .A(\ID_EXE_o[SIGN_EXTEND][18] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][18] ), .D(n154), .Z(n56) );
  HS65_LH_AO22X9 U124 ( .A(\ID_EXE_o[SIGN_EXTEND][19] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][19] ), .D(n154), .Z(n57) );
  HS65_LH_AO22X9 U125 ( .A(\ID_EXE_o[SIGN_EXTEND][20] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][20] ), .D(n154), .Z(n58) );
  HS65_LH_AO22X9 U126 ( .A(\ID_EXE_o[SIGN_EXTEND][21] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][21] ), .D(n154), .Z(n59) );
  HS65_LH_AO22X9 U127 ( .A(\ID_EXE_o[SIGN_EXTEND][22] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][22] ), .D(n154), .Z(n60) );
  HS65_LH_AO22X9 U128 ( .A(\ID_EXE_o[SIGN_EXTEND][23] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][23] ), .D(n154), .Z(n61) );
  HS65_LH_AO22X9 U129 ( .A(\ID_EXE_o[SIGN_EXTEND][24] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][24] ), .D(n155), .Z(n62) );
  HS65_LH_AO22X9 U130 ( .A(\ID_EXE_o[SIGN_EXTEND][25] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][25] ), .D(n155), .Z(n63) );
  HS65_LH_AO22X9 U131 ( .A(\ID_EXE_o[SIGN_EXTEND][26] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][26] ), .D(n155), .Z(n64) );
  HS65_LH_AO22X9 U132 ( .A(\ID_EXE_o[SIGN_EXTEND][27] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][27] ), .D(n155), .Z(n65) );
  HS65_LH_AO22X9 U133 ( .A(\ID_EXE_o[SIGN_EXTEND][28] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][28] ), .D(n155), .Z(n66) );
  HS65_LH_AO22X9 U134 ( .A(\ID_EXE_o[SIGN_EXTEND][29] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][29] ), .D(n155), .Z(n67) );
  HS65_LH_AO22X9 U135 ( .A(\ID_EXE_o[SIGN_EXTEND][30] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][30] ), .D(n155), .Z(n68) );
  HS65_LH_AO22X9 U136 ( .A(\ID_EXE_o[SIGN_EXTEND][31] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][31] ), .D(n155), .Z(n69) );
  HS65_LH_AO22X9 U137 ( .A(\ID_EXE_o[RD][0] ), .B(halt_i), .C(
        \ID_EXE_i[RD][0] ), .D(n150), .Z(n11) );
  HS65_LH_AO22X9 U138 ( .A(\ID_EXE_o[RD][1] ), .B(halt_i), .C(
        \ID_EXE_i[RD][1] ), .D(n150), .Z(n12) );
  HS65_LH_AO22X9 U139 ( .A(\ID_EXE_o[RD][2] ), .B(halt_i), .C(
        \ID_EXE_i[RD][2] ), .D(n150), .Z(n13) );
  HS65_LH_AO22X9 U140 ( .A(\ID_EXE_o[RD][3] ), .B(halt_i), .C(
        \ID_EXE_i[RD][3] ), .D(n151), .Z(n14) );
  HS65_LH_AO22X9 U141 ( .A(\ID_EXE_o[SIGN_EXTEND][0] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][0] ), .D(n153), .Z(n38) );
  HS65_LH_AO22X9 U142 ( .A(\ID_EXE_o[SIGN_EXTEND][1] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][1] ), .D(n153), .Z(n39) );
  HS65_LH_AO22X9 U143 ( .A(\ID_EXE_o[SIGN_EXTEND][2] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][2] ), .D(n153), .Z(n40) );
  HS65_LH_AO22X9 U144 ( .A(\ID_EXE_o[SIGN_EXTEND][3] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][3] ), .D(n153), .Z(n41) );
  HS65_LH_AO22X9 U145 ( .A(\ID_EXE_o[SIGN_EXTEND][4] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][4] ), .D(n153), .Z(n42) );
  HS65_LH_AO22X9 U146 ( .A(\ID_EXE_o[SIGN_EXTEND][5] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][5] ), .D(n153), .Z(n43) );
  HS65_LH_AO22X9 U147 ( .A(\ID_EXE_o[SIGN_EXTEND][6] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][6] ), .D(n153), .Z(n44) );
  HS65_LH_AO22X9 U148 ( .A(\ID_EXE_o[SIGN_EXTEND][7] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][7] ), .D(n153), .Z(n45) );
  HS65_LH_AO22X9 U149 ( .A(\ID_EXE_o[SIGN_EXTEND][8] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][8] ), .D(n153), .Z(n46) );
  HS65_LH_AO22X9 U150 ( .A(\ID_EXE_o[SIGN_EXTEND][9] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][9] ), .D(n153), .Z(n47) );
  HS65_LH_AO22X9 U151 ( .A(\ID_EXE_o[SIGN_EXTEND][10] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][10] ), .D(n153), .Z(n48) );
  HS65_LH_AO22X9 U152 ( .A(\ID_EXE_o[SIGN_EXTEND][11] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][11] ), .D(n153), .Z(n49) );
  HS65_LH_AO22X9 U153 ( .A(\ID_EXE_o[SIGN_EXTEND][12] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][12] ), .D(n154), .Z(n50) );
  HS65_LH_AO22X9 U154 ( .A(\ID_EXE_o[SIGN_EXTEND][13] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][13] ), .D(n154), .Z(n51) );
  HS65_LH_AO22X9 U155 ( .A(\ID_EXE_o[SIGN_EXTEND][14] ), .B(halt_i), .C(
        \ID_EXE_i[SIGN_EXTEND][14] ), .D(n154), .Z(n52) );
  HS65_LH_AO22X9 U156 ( .A(\ID_EXE_o[FUNCT][0] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][0] ), .D(n155), .Z(n70) );
  HS65_LH_AO22X9 U157 ( .A(\ID_EXE_o[FUNCT][1] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][1] ), .D(n155), .Z(n71) );
  HS65_LH_AO22X9 U158 ( .A(\ID_EXE_o[FUNCT][2] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][2] ), .D(n155), .Z(n72) );
  HS65_LH_AO22X9 U159 ( .A(\ID_EXE_o[FUNCT][3] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][3] ), .D(n155), .Z(n73) );
  HS65_LH_AO22X9 U160 ( .A(\ID_EXE_o[FUNCT][4] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][4] ), .D(n156), .Z(n74) );
  HS65_LH_AO22X9 U161 ( .A(\ID_EXE_o[FUNCT][5] ), .B(halt_i), .C(
        \ID_EXE_i[FUNCT][5] ), .D(n156), .Z(n75) );
  HS65_LH_AO22X9 U162 ( .A(\ID_EXE_o[SHAMT][0] ), .B(halt_i), .C(
        \ID_EXE_i[SHAMT][0] ), .D(n156), .Z(n76) );
  HS65_LH_AO22X9 U163 ( .A(\ID_EXE_o[SHAMT][1] ), .B(halt_i), .C(
        \ID_EXE_i[SHAMT][1] ), .D(n156), .Z(n77) );
  HS65_LH_AO22X9 U164 ( .A(\ID_EXE_o[SHAMT][2] ), .B(halt_i), .C(
        \ID_EXE_i[SHAMT][2] ), .D(n156), .Z(n78) );
  HS65_LH_AO22X9 U165 ( .A(\ID_EXE_o[SHAMT][3] ), .B(halt_i), .C(
        \ID_EXE_i[SHAMT][3] ), .D(n156), .Z(n79) );
  HS65_LH_AO22X9 U166 ( .A(\ID_EXE_o[SHAMT][4] ), .B(halt_i), .C(
        \ID_EXE_i[SHAMT][4] ), .D(n156), .Z(n80) );
  HS65_LH_AO22X9 U167 ( .A(\ID_EXE_o[MEMTOREG] ), .B(halt_i), .C(
        \ID_EXE_i[MEMTOREG] ), .D(n150), .Z(n9) );
  HS65_LH_AO22X9 U168 ( .A(\ID_EXE_o[PC_PLUS1][1] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][1] ), .D(n152), .Z(n27) );
  HS65_LH_AO22X9 U169 ( .A(\ID_EXE_o[PC_PLUS1][2] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][2] ), .D(n152), .Z(n28) );
  HS65_LH_AO22X9 U170 ( .A(\ID_EXE_o[PC_PLUS1][3] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][3] ), .D(n152), .Z(n29) );
  HS65_LH_AO22X9 U171 ( .A(\ID_EXE_o[PC_PLUS1][4] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][4] ), .D(n152), .Z(n30) );
  HS65_LH_AO22X9 U172 ( .A(\ID_EXE_o[PC_PLUS1][5] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][5] ), .D(n152), .Z(n31) );
  HS65_LH_AO22X9 U173 ( .A(\ID_EXE_o[PC_PLUS1][6] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][6] ), .D(n152), .Z(n32) );
  HS65_LH_AO22X9 U174 ( .A(\ID_EXE_o[PC_PLUS1][7] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][7] ), .D(n152), .Z(n33) );
  HS65_LH_AO22X9 U175 ( .A(\ID_EXE_o[PC_PLUS1][8] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][8] ), .D(n152), .Z(n34) );
  HS65_LH_AO22X9 U176 ( .A(\ID_EXE_o[PC_PLUS1][9] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][9] ), .D(n152), .Z(n35) );
  HS65_LH_AO22X9 U177 ( .A(\ID_EXE_o[PC_PLUS1][10] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][10] ), .D(n152), .Z(n36) );
  HS65_LH_AO22X9 U178 ( .A(\ID_EXE_o[PC_PLUS1][11] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][11] ), .D(n152), .Z(n37) );
  HS65_LH_AO22X9 U179 ( .A(\ID_EXE_o[PC_PLUS1][0] ), .B(halt_i), .C(
        \ID_EXE_i[PC_PLUS1][0] ), .D(n152), .Z(n26) );
  HS65_LH_AO22X9 U180 ( .A(\ID_EXE_o[CALU_OP][3] ), .B(halt_i), .C(
        \ID_EXE_i[CALU_OP][3] ), .D(n150), .Z(n6) );
  HS65_LH_IVX9 U181 ( .A(halt_i), .Z(n180) );
endmodule


module alu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328;

  HS65_LH_IVX9 U157 ( .A(n296), .Z(n247) );
  HS65_LH_IVX9 U158 ( .A(n305), .Z(n256) );
  HS65_LH_IVX9 U159 ( .A(n306), .Z(n260) );
  HS65_LH_OR2X9 U160 ( .A(B[11]), .B(n241), .Z(n327) );
  HS65_LH_IVX9 U161 ( .A(n279), .Z(n252) );
  HS65_LH_IVX9 U162 ( .A(n297), .Z(n246) );
  HS65_LH_IVX9 U163 ( .A(n284), .Z(n250) );
  HS65_LH_IVX9 U164 ( .A(n308), .Z(n263) );
  HS65_LH_IVX9 U165 ( .A(B[3]), .Z(n228) );
  HS65_LH_IVX9 U166 ( .A(B[4]), .Z(n229) );
  HS65_LH_IVX9 U167 ( .A(A[11]), .Z(n241) );
  HS65_LH_IVX9 U168 ( .A(A[17]), .Z(n243) );
  HS65_LH_IVX9 U169 ( .A(B[27]), .Z(n237) );
  HS65_LH_IVX9 U170 ( .A(B[2]), .Z(n227) );
  HS65_LH_IVX9 U171 ( .A(A[8]), .Z(n240) );
  HS65_LH_IVX9 U172 ( .A(A[14]), .Z(n242) );
  HS65_LH_IVX9 U173 ( .A(A[5]), .Z(n239) );
  HS65_LH_IVX9 U174 ( .A(A[20]), .Z(n244) );
  HS65_LH_IVX9 U175 ( .A(A[29]), .Z(n245) );
  HS65_LH_IVX9 U176 ( .A(n321), .Z(n257) );
  HS65_LH_IVX9 U177 ( .A(A[15]), .Z(n255) );
  HS65_LH_IVX9 U178 ( .A(A[7]), .Z(n264) );
  HS65_LH_IVX9 U179 ( .A(A[4]), .Z(n267) );
  HS65_LH_IVX9 U180 ( .A(n316), .Z(n266) );
  HS65_LH_IVX9 U181 ( .A(B[25]), .Z(n235) );
  HS65_LH_IVX9 U182 ( .A(A[1]), .Z(n268) );
  HS65_LH_IVX9 U183 ( .A(n320), .Z(n254) );
  HS65_LH_AND2X4 U184 ( .A(A[3]), .B(n228), .Z(n318) );
  HS65_LH_OR2X9 U185 ( .A(B[17]), .B(n243), .Z(n281) );
  HS65_LH_IVX9 U186 ( .A(A[9]), .Z(n262) );
  HS65_LH_IVX9 U187 ( .A(A[31]), .Z(n248) );
  HS65_LH_IVX9 U188 ( .A(A[16]), .Z(n253) );
  HS65_LH_IVX9 U189 ( .A(A[28]), .Z(n249) );
  HS65_LH_IVX9 U190 ( .A(A[21]), .Z(n251) );
  HS65_LH_IVX9 U191 ( .A(A[13]), .Z(n258) );
  HS65_LH_IVX9 U192 ( .A(A[12]), .Z(n259) );
  HS65_LH_IVX9 U193 ( .A(B[1]), .Z(n226) );
  HS65_LH_IVX9 U194 ( .A(B[23]), .Z(n233) );
  HS65_LH_IVX9 U195 ( .A(B[19]), .Z(n231) );
  HS65_LH_IVX9 U196 ( .A(B[26]), .Z(n236) );
  HS65_LH_IVX9 U197 ( .A(B[22]), .Z(n232) );
  HS65_LH_IVX9 U198 ( .A(B[18]), .Z(n230) );
  HS65_LH_IVX9 U199 ( .A(B[24]), .Z(n234) );
  HS65_LH_IVX9 U200 ( .A(B[30]), .Z(n238) );
  HS65_LH_IVX9 U201 ( .A(A[6]), .Z(n265) );
  HS65_LH_IVX9 U202 ( .A(A[10]), .Z(n261) );
  HS65_LH_OAI12X2 U203 ( .A(n269), .B(n270), .C(n271), .Z(GE_LT_GT_LE) );
  HS65_LH_OAI32X2 U204 ( .A(n272), .B(n273), .C(n274), .D(n275), .E(n272), .Z(
        n271) );
  HS65_LH_AOI212X2 U205 ( .A(n276), .B(n277), .C(n277), .D(n252), .E(n278), 
        .Z(n274) );
  HS65_LH_OA32X4 U206 ( .A(n230), .B(A[18]), .C(n280), .D(A[19]), .E(n231), 
        .Z(n277) );
  HS65_LH_AOI32X3 U207 ( .A(n281), .B(n253), .C(B[16]), .D(B[17]), .E(n243), 
        .Z(n276) );
  HS65_LH_AOI22X1 U208 ( .A(n282), .B(n283), .C(n283), .D(n250), .Z(n273) );
  HS65_LH_OA32X4 U209 ( .A(n232), .B(A[22]), .C(n285), .D(A[23]), .E(n233), 
        .Z(n283) );
  HS65_LH_AOI32X3 U210 ( .A(n286), .B(n244), .C(B[20]), .D(B[21]), .E(n251), 
        .Z(n282) );
  HS65_LH_CBI4I1X3 U211 ( .A(n247), .B(n246), .C(n287), .D(n288), .Z(n272) );
  HS65_LH_OAI212X3 U212 ( .A(n289), .B(n290), .C(n291), .D(n289), .E(n292), 
        .Z(n288) );
  HS65_LH_OAI32X2 U213 ( .A(n234), .B(A[24]), .C(n293), .D(A[25]), .E(n235), 
        .Z(n290) );
  HS65_LH_OAI32X2 U214 ( .A(n236), .B(A[26]), .C(n294), .D(A[27]), .E(n237), 
        .Z(n289) );
  HS65_LH_AOI312X2 U215 ( .A(n295), .B(n249), .C(B[28]), .D(B[29]), .E(n245), 
        .F(n296), .Z(n287) );
  HS65_LH_OAI32X2 U216 ( .A(n238), .B(A[30]), .C(n298), .D(B[31]), .E(n248), 
        .Z(n296) );
  HS65_LH_NAND3AX3 U217 ( .A(n278), .B(n279), .C(n275), .Z(n270) );
  HS65_LH_AND3X4 U218 ( .A(n291), .B(n292), .C(n299), .Z(n275) );
  HS65_LH_AOI12X2 U219 ( .A(A[24]), .B(n234), .C(n293), .Z(n299) );
  HS65_LH_NOR2AX3 U220 ( .A(A[25]), .B(B[25]), .Z(n293) );
  HS65_LH_OA112X4 U221 ( .A(B[28]), .B(n249), .C(n295), .D(n297), .Z(n292) );
  HS65_LH_AOI12X2 U222 ( .A(n238), .B(A[30]), .C(n298), .Z(n297) );
  HS65_LH_AND2X4 U223 ( .A(B[31]), .B(n248), .Z(n298) );
  HS65_LH_OR2X4 U224 ( .A(B[29]), .B(n245), .Z(n295) );
  HS65_LH_AOI12X2 U225 ( .A(n236), .B(A[26]), .C(n294), .Z(n291) );
  HS65_LH_AND2X4 U226 ( .A(A[27]), .B(n237), .Z(n294) );
  HS65_LH_AOI12X2 U227 ( .A(n230), .B(A[18]), .C(n280), .Z(n279) );
  HS65_LH_AND2X4 U228 ( .A(A[19]), .B(n231), .Z(n280) );
  HS65_LH_OAI112X1 U229 ( .A(B[20]), .B(n244), .C(n286), .D(n284), .Z(n278) );
  HS65_LH_AOI12X2 U230 ( .A(n232), .B(A[22]), .C(n285), .Z(n284) );
  HS65_LH_AND2X4 U231 ( .A(A[23]), .B(n233), .Z(n285) );
  HS65_LH_OR2X4 U232 ( .A(B[21]), .B(n251), .Z(n286) );
  HS65_LH_OAI212X3 U233 ( .A(n300), .B(n301), .C(n302), .D(n300), .E(n303), 
        .Z(n269) );
  HS65_LH_OA12X4 U234 ( .A(n253), .B(B[16]), .C(n281), .Z(n303) );
  HS65_LH_NOR3X1 U235 ( .A(n304), .B(n305), .C(n306), .Z(n302) );
  HS65_LH_OAI12X2 U236 ( .A(B[8]), .B(n240), .C(n307), .Z(n304) );
  HS65_LH_CBI4I1X3 U237 ( .A(n308), .B(n309), .C(n310), .D(n311), .Z(n301) );
  HS65_LH_NAND3AX3 U238 ( .A(n309), .B(n312), .C(n313), .Z(n311) );
  HS65_LH_AOI212X2 U239 ( .A(n314), .B(n315), .C(A[4]), .D(n229), .E(n316), 
        .Z(n313) );
  HS65_LH_AOI22X1 U240 ( .A(B[1]), .B(n268), .C(n317), .D(B[0]), .Z(n314) );
  HS65_LH_AOI12X2 U241 ( .A(A[1]), .B(n226), .C(A[0]), .Z(n317) );
  HS65_LH_CBI4I1X3 U242 ( .A(A[2]), .B(n227), .C(n318), .D(n315), .Z(n312) );
  HS65_LH_OA32X4 U243 ( .A(n227), .B(A[2]), .C(n318), .D(A[3]), .E(n228), .Z(
        n315) );
  HS65_LH_AOI312X2 U244 ( .A(n266), .B(n267), .C(B[4]), .D(B[5]), .E(n239), 
        .F(n263), .Z(n310) );
  HS65_LH_NOR2X2 U245 ( .A(n239), .B(B[5]), .Z(n316) );
  HS65_LH_OAI12X2 U246 ( .A(B[6]), .B(n265), .C(n319), .Z(n309) );
  HS65_LH_AOI32X3 U247 ( .A(B[6]), .B(n265), .C(n319), .D(n264), .E(B[7]), .Z(
        n308) );
  HS65_LH_NAND2AX4 U248 ( .A(B[7]), .B(A[7]), .Z(n319) );
  HS65_LH_CBI4I1X3 U249 ( .A(n320), .B(n321), .C(n322), .D(n323), .Z(n300) );
  HS65_LH_OAI212X3 U250 ( .A(n324), .B(n325), .C(n260), .D(n324), .E(n256), 
        .Z(n323) );
  HS65_LH_OAI112X1 U251 ( .A(B[12]), .B(n259), .C(n326), .D(n257), .Z(n305) );
  HS65_LH_OAI12X2 U252 ( .A(B[10]), .B(n261), .C(n327), .Z(n306) );
  HS65_LH_AO32X4 U253 ( .A(B[8]), .B(n240), .C(n307), .D(n262), .E(B[9]), .Z(
        n325) );
  HS65_LH_NAND2AX4 U254 ( .A(B[9]), .B(A[9]), .Z(n307) );
  HS65_LH_AO32X4 U255 ( .A(B[10]), .B(n261), .C(n327), .D(n241), .E(B[11]), 
        .Z(n324) );
  HS65_LH_AOI312X2 U256 ( .A(n326), .B(n259), .C(B[12]), .D(B[13]), .E(n258), 
        .F(n254), .Z(n322) );
  HS65_LH_OR2X4 U257 ( .A(B[13]), .B(n258), .Z(n326) );
  HS65_LH_OAI12X2 U258 ( .A(B[14]), .B(n242), .C(n328), .Z(n321) );
  HS65_LH_AOI32X3 U259 ( .A(B[14]), .B(n242), .C(n328), .D(n255), .E(B[15]), 
        .Z(n320) );
  HS65_LH_NAND2AX4 U260 ( .A(B[15]), .B(A[15]), .Z(n328) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  HS65_LH_FA1X4 U2_23 ( .A0(A[23]), .B0(n25), .CI(carry[23]), .CO(carry[24]), 
        .S0(DIFF[23]) );
  HS65_LH_FA1X4 U2_29 ( .A0(A[29]), .B0(n31), .CI(carry[29]), .CO(carry[30]), 
        .S0(DIFF[29]) );
  HS65_LH_FA1X4 U2_26 ( .A0(A[26]), .B0(n28), .CI(carry[26]), .CO(carry[27]), 
        .S0(DIFF[26]) );
  HS65_LH_FA1X4 U2_17 ( .A0(A[17]), .B0(n19), .CI(carry[17]), .CO(carry[18]), 
        .S0(DIFF[17]) );
  HS65_LH_FA1X4 U2_5 ( .A0(A[5]), .B0(n7), .CI(carry[5]), .CO(carry[6]), .S0(
        DIFF[5]) );
  HS65_LH_FA1X4 U2_14 ( .A0(A[14]), .B0(n16), .CI(carry[14]), .CO(carry[15]), 
        .S0(DIFF[14]) );
  HS65_LH_FA1X4 U2_8 ( .A0(A[8]), .B0(n10), .CI(carry[8]), .CO(carry[9]), .S0(
        DIFF[8]) );
  HS65_LH_FA1X4 U2_3 ( .A0(A[3]), .B0(n5), .CI(carry[3]), .CO(carry[4]), .S0(
        DIFF[3]) );
  HS65_LH_FA1X4 U2_1 ( .A0(A[1]), .B0(n3), .CI(carry[1]), .CO(carry[2]), .S0(
        DIFF[1]) );
  HS65_LH_FA1X4 U2_9 ( .A0(A[9]), .B0(n11), .CI(carry[9]), .CO(carry[10]), 
        .S0(DIFF[9]) );
  HS65_LH_FA1X4 U2_7 ( .A0(A[7]), .B0(n9), .CI(carry[7]), .CO(carry[8]), .S0(
        DIFF[7]) );
  HS65_LH_FA1X4 U2_10 ( .A0(A[10]), .B0(n12), .CI(carry[10]), .CO(carry[11]), 
        .S0(DIFF[10]) );
  HS65_LH_FA1X4 U2_6 ( .A0(A[6]), .B0(n8), .CI(carry[6]), .CO(carry[7]), .S0(
        DIFF[6]) );
  HS65_LH_FA1X4 U2_4 ( .A0(A[4]), .B0(n6), .CI(carry[4]), .CO(carry[5]), .S0(
        DIFF[4]) );
  HS65_LH_FA1X4 U2_30 ( .A0(A[30]), .B0(n32), .CI(carry[30]), .CO(carry[31]), 
        .S0(DIFF[30]) );
  HS65_LH_FA1X4 U2_25 ( .A0(A[25]), .B0(n27), .CI(carry[25]), .CO(carry[26]), 
        .S0(DIFF[25]) );
  HS65_LH_FA1X4 U2_19 ( .A0(A[19]), .B0(n21), .CI(carry[19]), .CO(carry[20]), 
        .S0(DIFF[19]) );
  HS65_LH_FA1X4 U2_27 ( .A0(A[27]), .B0(n29), .CI(carry[27]), .CO(carry[28]), 
        .S0(DIFF[27]) );
  HS65_LH_FA1X4 U2_24 ( .A0(A[24]), .B0(n26), .CI(carry[24]), .CO(carry[25]), 
        .S0(DIFF[24]) );
  HS65_LH_FA1X4 U2_21 ( .A0(A[21]), .B0(n23), .CI(carry[21]), .CO(carry[22]), 
        .S0(DIFF[21]) );
  HS65_LH_FA1X4 U2_18 ( .A0(A[18]), .B0(n20), .CI(carry[18]), .CO(carry[19]), 
        .S0(DIFF[18]) );
  HS65_LH_FA1X4 U2_13 ( .A0(A[13]), .B0(n15), .CI(carry[13]), .CO(carry[14]), 
        .S0(DIFF[13]) );
  HS65_LH_FA1X4 U2_12 ( .A0(A[12]), .B0(n14), .CI(carry[12]), .CO(carry[13]), 
        .S0(DIFF[12]) );
  HS65_LH_FA1X4 U2_22 ( .A0(A[22]), .B0(n24), .CI(carry[22]), .CO(carry[23]), 
        .S0(DIFF[22]) );
  HS65_LH_FA1X4 U2_15 ( .A0(A[15]), .B0(n17), .CI(carry[15]), .CO(carry[16]), 
        .S0(DIFF[15]) );
  HS65_LH_FA1X4 U2_28 ( .A0(A[28]), .B0(n30), .CI(carry[28]), .CO(carry[29]), 
        .S0(DIFF[28]) );
  HS65_LH_FA1X4 U2_16 ( .A0(A[16]), .B0(n18), .CI(carry[16]), .CO(carry[17]), 
        .S0(DIFF[16]) );
  HS65_LHS_XOR3X2 U2_31 ( .A(A[31]), .B(n33), .C(carry[31]), .Z(DIFF[31]) );
  HS65_LH_FA1X4 U2_2 ( .A0(A[2]), .B0(n4), .CI(carry[2]), .CO(carry[3]), .S0(
        DIFF[2]) );
  HS65_LH_FA1X4 U2_20 ( .A0(A[20]), .B0(n22), .CI(carry[20]), .CO(carry[21]), 
        .S0(DIFF[20]) );
  HS65_LH_FA1X4 U2_11 ( .A0(A[11]), .B0(n13), .CI(carry[11]), .CO(carry[12]), 
        .S0(DIFF[11]) );
  HS65_LH_IVX9 U1 ( .A(B[11]), .Z(n13) );
  HS65_LH_IVX9 U2 ( .A(B[20]), .Z(n22) );
  HS65_LH_IVX9 U3 ( .A(B[2]), .Z(n4) );
  HS65_LH_IVX9 U4 ( .A(B[31]), .Z(n33) );
  HS65_LH_IVX9 U5 ( .A(B[16]), .Z(n18) );
  HS65_LH_IVX9 U6 ( .A(B[28]), .Z(n30) );
  HS65_LH_IVX9 U7 ( .A(B[15]), .Z(n17) );
  HS65_LH_IVX9 U8 ( .A(B[22]), .Z(n24) );
  HS65_LH_IVX9 U9 ( .A(B[12]), .Z(n14) );
  HS65_LH_IVX9 U10 ( .A(B[13]), .Z(n15) );
  HS65_LH_IVX9 U11 ( .A(B[18]), .Z(n20) );
  HS65_LH_IVX9 U12 ( .A(B[21]), .Z(n23) );
  HS65_LH_IVX9 U13 ( .A(B[24]), .Z(n26) );
  HS65_LH_IVX9 U14 ( .A(B[27]), .Z(n29) );
  HS65_LH_IVX9 U15 ( .A(B[19]), .Z(n21) );
  HS65_LH_IVX9 U16 ( .A(B[25]), .Z(n27) );
  HS65_LH_IVX9 U17 ( .A(B[30]), .Z(n32) );
  HS65_LH_IVX9 U18 ( .A(B[4]), .Z(n6) );
  HS65_LH_IVX9 U19 ( .A(B[6]), .Z(n8) );
  HS65_LH_IVX9 U20 ( .A(B[10]), .Z(n12) );
  HS65_LH_IVX9 U21 ( .A(B[7]), .Z(n9) );
  HS65_LH_IVX9 U22 ( .A(B[9]), .Z(n11) );
  HS65_LH_IVX9 U23 ( .A(B[1]), .Z(n3) );
  HS65_LH_NAND2X7 U24 ( .A(n1), .B(B[0]), .Z(carry[1]) );
  HS65_LH_IVX9 U25 ( .A(B[3]), .Z(n5) );
  HS65_LH_IVX9 U26 ( .A(B[8]), .Z(n10) );
  HS65_LH_IVX9 U27 ( .A(B[14]), .Z(n16) );
  HS65_LH_IVX9 U28 ( .A(B[5]), .Z(n7) );
  HS65_LH_IVX9 U29 ( .A(B[17]), .Z(n19) );
  HS65_LH_IVX9 U30 ( .A(B[26]), .Z(n28) );
  HS65_LH_IVX9 U31 ( .A(B[29]), .Z(n31) );
  HS65_LH_IVX9 U32 ( .A(B[23]), .Z(n25) );
  HS65_LH_IVX9 U33 ( .A(A[0]), .Z(n1) );
  HS65_LH_IVX9 U34 ( .A(B[0]), .Z(n2) );
  HS65_LHS_XNOR2X6 U35 ( .A(A[0]), .B(n2), .Z(DIFF[0]) );
endmodule


module alu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114;

  HS65_LH_IVX9 U1 ( .A(n114), .Z(n39) );
  HS65_LH_IVX9 U2 ( .A(n53), .Z(n34) );
  HS65_LH_IVX9 U3 ( .A(n101), .Z(n37) );
  HS65_LH_IVX9 U4 ( .A(B[2]), .Z(n1) );
  HS65_LH_IVX9 U5 ( .A(A[14]), .Z(n21) );
  HS65_LH_IVX9 U6 ( .A(B[3]), .Z(n2) );
  HS65_LH_IVX9 U7 ( .A(B[11]), .Z(n6) );
  HS65_LH_IVX9 U8 ( .A(A[8]), .Z(n20) );
  HS65_LH_IVX9 U9 ( .A(A[26]), .Z(n22) );
  HS65_LH_IVX9 U10 ( .A(B[27]), .Z(n16) );
  HS65_LH_IVX9 U11 ( .A(B[20]), .Z(n12) );
  HS65_LH_IVX9 U12 ( .A(B[28]), .Z(n17) );
  HS65_LH_IVX9 U13 ( .A(B[31]), .Z(n19) );
  HS65_LH_IVX9 U14 ( .A(n66), .Z(n26) );
  HS65_LH_IVX9 U15 ( .A(n75), .Z(n23) );
  HS65_LH_IVX9 U16 ( .A(n59), .Z(n24) );
  HS65_LH_IVX9 U17 ( .A(A[22]), .Z(n29) );
  HS65_LH_IVX9 U18 ( .A(n70), .Z(n32) );
  HS65_LH_IVX9 U19 ( .A(n50), .Z(n36) );
  HS65_LH_IVX9 U20 ( .A(n63), .Z(n27) );
  HS65_LH_IVX9 U21 ( .A(A[6]), .Z(n38) );
  HS65_LH_IVX9 U22 ( .A(n69), .Z(n30) );
  HS65_LH_OR2X9 U23 ( .A(B[14]), .B(n21), .Z(n49) );
  HS65_LH_IVX9 U24 ( .A(B[12]), .Z(n7) );
  HS65_LH_IVX9 U25 ( .A(B[13]), .Z(n8) );
  HS65_LH_IVX9 U26 ( .A(B[15]), .Z(n9) );
  HS65_LH_IVX9 U27 ( .A(B[7]), .Z(n4) );
  HS65_LH_IVX9 U28 ( .A(B[5]), .Z(n3) );
  HS65_LH_IVX9 U29 ( .A(B[9]), .Z(n5) );
  HS65_LH_IVX9 U30 ( .A(A[1]), .Z(n41) );
  HS65_LH_IVX9 U31 ( .A(A[4]), .Z(n40) );
  HS65_LH_IVX9 U32 ( .A(A[10]), .Z(n35) );
  HS65_LH_OR2X9 U33 ( .A(B[26]), .B(n22), .Z(n65) );
  HS65_LH_IVX9 U34 ( .A(A[16]), .Z(n33) );
  HS65_LH_IVX9 U35 ( .A(A[24]), .Z(n28) );
  HS65_LH_IVX9 U36 ( .A(A[18]), .Z(n31) );
  HS65_LH_IVX9 U37 ( .A(B[23]), .Z(n14) );
  HS65_LH_IVX9 U38 ( .A(B[19]), .Z(n11) );
  HS65_LH_IVX9 U39 ( .A(B[25]), .Z(n15) );
  HS65_LH_IVX9 U40 ( .A(B[21]), .Z(n13) );
  HS65_LH_IVX9 U41 ( .A(B[17]), .Z(n10) );
  HS65_LH_IVX9 U42 ( .A(A[30]), .Z(n25) );
  HS65_LH_IVX9 U43 ( .A(B[29]), .Z(n18) );
  HS65_LH_CNIVX3 U44 ( .A(EQ), .Z(NE) );
  HS65_LH_NOR4ABX2 U45 ( .A(n42), .B(n43), .C(n44), .D(n45), .Z(EQ) );
  HS65_LH_NAND4X4 U46 ( .A(n46), .B(n47), .C(n48), .D(n49), .Z(n45) );
  HS65_LH_NAND4ABX3 U47 ( .A(n50), .B(n34), .C(n51), .D(n52), .Z(n44) );
  HS65_LH_NOR4ABX2 U48 ( .A(n54), .B(n55), .C(n56), .D(n57), .Z(n43) );
  HS65_LH_NAND4ABX3 U49 ( .A(n58), .B(n59), .C(n60), .D(n61), .Z(n57) );
  HS65_LH_AOI22X1 U50 ( .A(n41), .B(n62), .C(n62), .D(B[1]), .Z(n58) );
  HS65_LH_NAND2AX4 U51 ( .A(B[0]), .B(A[0]), .Z(n62) );
  HS65_LH_NAND4ABX3 U52 ( .A(n63), .B(n26), .C(n64), .D(n65), .Z(n56) );
  HS65_LH_NOR4ABX2 U53 ( .A(n67), .B(n68), .C(n69), .D(n70), .Z(n55) );
  HS65_LH_AND4X3 U54 ( .A(n71), .B(n72), .C(n73), .D(n74), .Z(n54) );
  HS65_LH_NOR4ABX2 U55 ( .A(n75), .B(n76), .C(n77), .D(LT), .Z(n42) );
  HS65_LH_OAI22X1 U56 ( .A(A[31]), .B(n19), .C(n23), .D(n78), .Z(LT) );
  HS65_LH_AOI32X3 U57 ( .A(n61), .B(n24), .C(n79), .D(B[30]), .E(n25), .Z(n78)
         );
  HS65_LH_OAI212X3 U58 ( .A(A[28]), .B(n17), .C(A[29]), .D(n18), .E(n80), .Z(
        n79) );
  HS65_LH_NAND3X2 U59 ( .A(n60), .B(n66), .C(n81), .Z(n80) );
  HS65_LH_OAI12X2 U60 ( .A(A[27]), .B(n16), .C(n82), .Z(n81) );
  HS65_LH_AOI32X3 U61 ( .A(n65), .B(n64), .C(n83), .D(B[26]), .E(n22), .Z(n82)
         );
  HS65_LH_OAI12X2 U62 ( .A(A[25]), .B(n15), .C(n84), .Z(n83) );
  HS65_LH_AOI32X3 U63 ( .A(n27), .B(n71), .C(n85), .D(B[24]), .E(n28), .Z(n84)
         );
  HS65_LH_OAI12X2 U64 ( .A(A[23]), .B(n14), .C(n86), .Z(n85) );
  HS65_LH_AOI32X3 U65 ( .A(n72), .B(n74), .C(n87), .D(B[22]), .E(n29), .Z(n86)
         );
  HS65_LH_OAI212X3 U66 ( .A(A[20]), .B(n12), .C(A[21]), .D(n13), .E(n88), .Z(
        n87) );
  HS65_LH_NAND3X2 U67 ( .A(n73), .B(n67), .C(n89), .Z(n88) );
  HS65_LH_OAI12X2 U68 ( .A(A[19]), .B(n11), .C(n90), .Z(n89) );
  HS65_LH_AOI32X3 U69 ( .A(n30), .B(n68), .C(n91), .D(B[18]), .E(n31), .Z(n90)
         );
  HS65_LH_OAI12X2 U70 ( .A(A[17]), .B(n10), .C(n92), .Z(n91) );
  HS65_LH_AOI32X3 U71 ( .A(n32), .B(n48), .C(n93), .D(B[16]), .E(n33), .Z(n92)
         );
  HS65_LH_OAI12X2 U72 ( .A(A[15]), .B(n9), .C(n94), .Z(n93) );
  HS65_LH_AOI32X3 U73 ( .A(n49), .B(n47), .C(n95), .D(B[14]), .E(n21), .Z(n94)
         );
  HS65_LH_OAI212X3 U74 ( .A(A[12]), .B(n7), .C(A[13]), .D(n8), .E(n96), .Z(n95) );
  HS65_LH_NAND3X2 U75 ( .A(n46), .B(n53), .C(n97), .Z(n96) );
  HS65_LH_OAI12X2 U76 ( .A(A[11]), .B(n6), .C(n98), .Z(n97) );
  HS65_LH_AOI32X3 U77 ( .A(n52), .B(n51), .C(n99), .D(B[10]), .E(n35), .Z(n98)
         );
  HS65_LH_OAI12X2 U78 ( .A(A[9]), .B(n5), .C(n100), .Z(n99) );
  HS65_LH_AOI32X3 U79 ( .A(n36), .B(n101), .C(n102), .D(B[8]), .E(n20), .Z(
        n100) );
  HS65_LH_OAI12X2 U80 ( .A(A[7]), .B(n4), .C(n103), .Z(n102) );
  HS65_LH_AOI32X3 U81 ( .A(n104), .B(n105), .C(n106), .D(B[6]), .E(n38), .Z(
        n103) );
  HS65_LH_OAI12X2 U82 ( .A(A[5]), .B(n3), .C(n107), .Z(n106) );
  HS65_LH_AOI32X3 U83 ( .A(n39), .B(n108), .C(n109), .D(B[4]), .E(n40), .Z(
        n107) );
  HS65_LH_OAI212X3 U84 ( .A(A[2]), .B(n1), .C(A[3]), .D(n2), .E(n110), .Z(n109) );
  HS65_LH_OAI212X3 U85 ( .A(B[1]), .B(n111), .C(n112), .D(n41), .E(n113), .Z(
        n110) );
  HS65_LH_AND2X4 U86 ( .A(n112), .B(n41), .Z(n111) );
  HS65_LH_NOR2AX3 U87 ( .A(B[0]), .B(A[0]), .Z(n112) );
  HS65_LH_NOR2X2 U88 ( .A(n20), .B(B[8]), .Z(n50) );
  HS65_LH_NAND2X2 U89 ( .A(A[9]), .B(n5), .Z(n51) );
  HS65_LH_NAND2AX4 U90 ( .A(B[10]), .B(A[10]), .Z(n52) );
  HS65_LH_NAND2X2 U91 ( .A(A[11]), .B(n6), .Z(n53) );
  HS65_LH_NAND2X2 U92 ( .A(A[12]), .B(n7), .Z(n46) );
  HS65_LH_NAND2X2 U93 ( .A(A[13]), .B(n8), .Z(n47) );
  HS65_LH_NAND2X2 U94 ( .A(A[15]), .B(n9), .Z(n48) );
  HS65_LH_NOR2X2 U95 ( .A(n33), .B(B[16]), .Z(n70) );
  HS65_LH_NAND2X2 U96 ( .A(A[17]), .B(n10), .Z(n68) );
  HS65_LH_NOR2X2 U97 ( .A(B[18]), .B(n31), .Z(n69) );
  HS65_LH_NAND2X2 U98 ( .A(A[19]), .B(n11), .Z(n67) );
  HS65_LH_NAND2X2 U99 ( .A(A[20]), .B(n12), .Z(n73) );
  HS65_LH_NAND2X2 U100 ( .A(A[21]), .B(n13), .Z(n74) );
  HS65_LH_NAND2AX4 U101 ( .A(B[22]), .B(A[22]), .Z(n72) );
  HS65_LH_NAND2X2 U102 ( .A(A[23]), .B(n14), .Z(n71) );
  HS65_LH_NOR2X2 U103 ( .A(n28), .B(B[24]), .Z(n63) );
  HS65_LH_NAND2X2 U104 ( .A(A[25]), .B(n15), .Z(n64) );
  HS65_LH_NAND2X2 U105 ( .A(A[27]), .B(n16), .Z(n66) );
  HS65_LH_NAND2X2 U106 ( .A(A[28]), .B(n17), .Z(n60) );
  HS65_LH_NOR2X2 U107 ( .A(n25), .B(B[30]), .Z(n59) );
  HS65_LH_NAND2X2 U108 ( .A(A[29]), .B(n18), .Z(n61) );
  HS65_LH_NAND4ABX3 U109 ( .A(n114), .B(n37), .C(n105), .D(n104), .Z(n77) );
  HS65_LH_NAND2AX4 U110 ( .A(B[6]), .B(A[6]), .Z(n104) );
  HS65_LH_NAND2X2 U111 ( .A(A[5]), .B(n3), .Z(n105) );
  HS65_LH_NAND2X2 U112 ( .A(A[7]), .B(n4), .Z(n101) );
  HS65_LH_NOR2X2 U113 ( .A(n40), .B(B[4]), .Z(n114) );
  HS65_LH_AND2X4 U114 ( .A(n113), .B(n108), .Z(n76) );
  HS65_LH_NAND2X2 U115 ( .A(A[3]), .B(n2), .Z(n108) );
  HS65_LH_NAND2X2 U116 ( .A(A[2]), .B(n1), .Z(n113) );
  HS65_LH_NAND2X2 U117 ( .A(A[31]), .B(n19), .Z(n75) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  HS65_LH_FA1X4 U1_23 ( .A0(A[23]), .B0(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S0(SUM[23]) );
  HS65_LH_FA1X4 U1_29 ( .A0(A[29]), .B0(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S0(SUM[29]) );
  HS65_LH_FA1X4 U1_26 ( .A0(A[26]), .B0(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S0(SUM[26]) );
  HS65_LH_FA1X4 U1_17 ( .A0(A[17]), .B0(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S0(SUM[17]) );
  HS65_LH_FA1X4 U1_5 ( .A0(A[5]), .B0(B[5]), .CI(carry[5]), .CO(carry[6]), 
        .S0(SUM[5]) );
  HS65_LH_FA1X4 U1_14 ( .A0(A[14]), .B0(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S0(SUM[14]) );
  HS65_LH_FA1X4 U1_8 ( .A0(A[8]), .B0(B[8]), .CI(carry[8]), .CO(carry[9]), 
        .S0(SUM[8]) );
  HS65_LH_FA1X4 U1_3 ( .A0(A[3]), .B0(B[3]), .CI(carry[3]), .CO(carry[4]), 
        .S0(SUM[3]) );
  HS65_LH_FA1X4 U1_1 ( .A0(A[1]), .B0(B[1]), .CI(n1), .CO(carry[2]), .S0(
        SUM[1]) );
  HS65_LH_FA1X4 U1_9 ( .A0(A[9]), .B0(B[9]), .CI(carry[9]), .CO(carry[10]), 
        .S0(SUM[9]) );
  HS65_LH_FA1X4 U1_7 ( .A0(A[7]), .B0(B[7]), .CI(carry[7]), .CO(carry[8]), 
        .S0(SUM[7]) );
  HS65_LH_FA1X4 U1_10 ( .A0(A[10]), .B0(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S0(SUM[10]) );
  HS65_LH_FA1X4 U1_6 ( .A0(A[6]), .B0(B[6]), .CI(carry[6]), .CO(carry[7]), 
        .S0(SUM[6]) );
  HS65_LH_FA1X4 U1_4 ( .A0(A[4]), .B0(B[4]), .CI(carry[4]), .CO(carry[5]), 
        .S0(SUM[4]) );
  HS65_LH_FA1X4 U1_30 ( .A0(A[30]), .B0(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S0(SUM[30]) );
  HS65_LH_FA1X4 U1_25 ( .A0(A[25]), .B0(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S0(SUM[25]) );
  HS65_LH_FA1X4 U1_19 ( .A0(A[19]), .B0(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S0(SUM[19]) );
  HS65_LH_FA1X4 U1_27 ( .A0(A[27]), .B0(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S0(SUM[27]) );
  HS65_LH_FA1X4 U1_24 ( .A0(A[24]), .B0(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S0(SUM[24]) );
  HS65_LH_FA1X4 U1_21 ( .A0(A[21]), .B0(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S0(SUM[21]) );
  HS65_LH_FA1X4 U1_18 ( .A0(A[18]), .B0(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S0(SUM[18]) );
  HS65_LH_FA1X4 U1_13 ( .A0(A[13]), .B0(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S0(SUM[13]) );
  HS65_LH_FA1X4 U1_12 ( .A0(A[12]), .B0(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S0(SUM[12]) );
  HS65_LH_FA1X4 U1_22 ( .A0(A[22]), .B0(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S0(SUM[22]) );
  HS65_LH_FA1X4 U1_15 ( .A0(A[15]), .B0(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S0(SUM[15]) );
  HS65_LH_FA1X4 U1_28 ( .A0(A[28]), .B0(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S0(SUM[28]) );
  HS65_LH_FA1X4 U1_16 ( .A0(A[16]), .B0(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S0(SUM[16]) );
  HS65_LHS_XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Z(SUM[31]) );
  HS65_LH_FA1X4 U1_2 ( .A0(A[2]), .B0(B[2]), .CI(carry[2]), .CO(carry[3]), 
        .S0(SUM[2]) );
  HS65_LH_FA1X4 U1_20 ( .A0(A[20]), .B0(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S0(SUM[20]) );
  HS65_LH_FA1X4 U1_11 ( .A0(A[11]), .B0(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S0(SUM[11]) );
  HS65_LH_AND2X4 U1 ( .A(A[0]), .B(B[0]), .Z(n1) );
  HS65_LHS_XOR2X6 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module alu_DW_mult_uns_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n7, n19, n31, n43, n55, n67, n79, n91, n103, n115, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n292, n293, n294, n295, n296, n297,
         n299, n300, n302, n303, n304, n305, n306, n307, n308, n309, n311,
         n312, n313, n314, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
         n360, n361, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105;
  assign n7 = a[2];
  assign n19 = a[5];
  assign n31 = a[8];
  assign n43 = a[11];
  assign n55 = a[14];
  assign n67 = a[17];
  assign n79 = a[20];
  assign n91 = a[23];
  assign n103 = a[26];
  assign n115 = a[29];

  HS65_LH_FA1X4 U228 ( .A0(n293), .B0(n292), .CI(n228), .CO(n227), .S0(
        product[62]) );
  HS65_LH_FA1X4 U229 ( .A0(n295), .B0(n294), .CI(n229), .CO(n228), .S0(
        product[61]) );
  HS65_LH_FA1X4 U230 ( .A0(n296), .B0(n299), .CI(n230), .CO(n229), .S0(
        product[60]) );
  HS65_LH_FA1X4 U231 ( .A0(n300), .B0(n302), .CI(n231), .CO(n230), .S0(
        product[59]) );
  HS65_LH_FA1X4 U232 ( .A0(n303), .B0(n305), .CI(n232), .CO(n231), .S0(
        product[58]) );
  HS65_LH_FA1X4 U233 ( .A0(n306), .B0(n311), .CI(n233), .CO(n232), .S0(
        product[57]) );
  HS65_LH_FA1X4 U234 ( .A0(n312), .B0(n316), .CI(n234), .CO(n233), .S0(
        product[56]) );
  HS65_LH_FA1X4 U235 ( .A0(n317), .B0(n322), .CI(n235), .CO(n234), .S0(
        product[55]) );
  HS65_LH_FA1X4 U236 ( .A0(n323), .B0(n330), .CI(n236), .CO(n235), .S0(
        product[54]) );
  HS65_LH_FA1X4 U237 ( .A0(n331), .B0(n337), .CI(n237), .CO(n236), .S0(
        product[53]) );
  HS65_LH_FA1X4 U238 ( .A0(n338), .B0(n344), .CI(n238), .CO(n237), .S0(
        product[52]) );
  HS65_LH_FA1X4 U239 ( .A0(n345), .B0(n354), .CI(n239), .CO(n238), .S0(
        product[51]) );
  HS65_LH_FA1X4 U240 ( .A0(n355), .B0(n363), .CI(n240), .CO(n239), .S0(
        product[50]) );
  HS65_LH_FA1X4 U241 ( .A0(n364), .B0(n373), .CI(n241), .CO(n240), .S0(
        product[49]) );
  HS65_LH_FA1X4 U242 ( .A0(n374), .B0(n385), .CI(n242), .CO(n241), .S0(
        product[48]) );
  HS65_LH_FA1X4 U243 ( .A0(n386), .B0(n396), .CI(n243), .CO(n242), .S0(
        product[47]) );
  HS65_LH_FA1X4 U244 ( .A0(n397), .B0(n407), .CI(n244), .CO(n243), .S0(
        product[46]) );
  HS65_LH_FA1X4 U245 ( .A0(n408), .B0(n421), .CI(n245), .CO(n244), .S0(
        product[45]) );
  HS65_LH_FA1X4 U246 ( .A0(n422), .B0(n434), .CI(n246), .CO(n245), .S0(
        product[44]) );
  HS65_LH_FA1X4 U247 ( .A0(n435), .B0(n448), .CI(n247), .CO(n246), .S0(
        product[43]) );
  HS65_LH_FA1X4 U248 ( .A0(n449), .B0(n464), .CI(n248), .CO(n247), .S0(
        product[42]) );
  HS65_LH_FA1X4 U249 ( .A0(n465), .B0(n479), .CI(n249), .CO(n248), .S0(
        product[41]) );
  HS65_LH_FA1X4 U250 ( .A0(n480), .B0(n494), .CI(n250), .CO(n249), .S0(
        product[40]) );
  HS65_LH_FA1X4 U251 ( .A0(n495), .B0(n512), .CI(n251), .CO(n250), .S0(
        product[39]) );
  HS65_LH_FA1X4 U252 ( .A0(n513), .B0(n529), .CI(n252), .CO(n251), .S0(
        product[38]) );
  HS65_LH_FA1X4 U253 ( .A0(n530), .B0(n546), .CI(n253), .CO(n252), .S0(
        product[37]) );
  HS65_LH_FA1X4 U254 ( .A0(n547), .B0(n564), .CI(n254), .CO(n253), .S0(
        product[36]) );
  HS65_LH_FA1X4 U255 ( .A0(n565), .B0(n582), .CI(n255), .CO(n254), .S0(
        product[35]) );
  HS65_LH_FA1X4 U256 ( .A0(n583), .B0(n600), .CI(n256), .CO(n255), .S0(
        product[34]) );
  HS65_LH_FA1X4 U257 ( .A0(n601), .B0(n1386), .CI(n257), .CO(n256), .S0(
        product[33]) );
  HS65_LH_FA1X4 U258 ( .A0(n1387), .B0(n619), .CI(n258), .CO(n257), .S0(
        product[32]) );
  HS65_LH_FA1X4 U259 ( .A0(n1388), .B0(n637), .CI(n259), .CO(n258), .S0(
        product[31]) );
  HS65_LH_FA1X4 U260 ( .A0(n1389), .B0(n655), .CI(n260), .CO(n259), .S0(
        product[30]) );
  HS65_LH_FA1X4 U261 ( .A0(n1390), .B0(n673), .CI(n261), .CO(n260), .S0(
        product[29]) );
  HS65_LH_FA1X4 U262 ( .A0(n1391), .B0(n691), .CI(n262), .CO(n261), .S0(
        product[28]) );
  HS65_LH_FA1X4 U263 ( .A0(n1392), .B0(n709), .CI(n263), .CO(n262), .S0(
        product[27]) );
  HS65_LH_FA1X4 U264 ( .A0(n1393), .B0(n727), .CI(n264), .CO(n263), .S0(
        product[26]) );
  HS65_LH_FA1X4 U265 ( .A0(n1394), .B0(n743), .CI(n265), .CO(n264), .S0(
        product[25]) );
  HS65_LH_FA1X4 U266 ( .A0(n1395), .B0(n759), .CI(n266), .CO(n265), .S0(
        product[24]) );
  HS65_LH_FA1X4 U267 ( .A0(n1396), .B0(n775), .CI(n267), .CO(n266), .S0(
        product[23]) );
  HS65_LH_FA1X4 U268 ( .A0(n1397), .B0(n789), .CI(n268), .CO(n267), .S0(
        product[22]) );
  HS65_LH_FA1X4 U269 ( .A0(n1398), .B0(n803), .CI(n269), .CO(n268), .S0(
        product[21]) );
  HS65_LH_FA1X4 U270 ( .A0(n1399), .B0(n817), .CI(n270), .CO(n269), .S0(
        product[20]) );
  HS65_LH_FA1X4 U271 ( .A0(n1400), .B0(n829), .CI(n271), .CO(n270), .S0(
        product[19]) );
  HS65_LH_FA1X4 U272 ( .A0(n1401), .B0(n841), .CI(n272), .CO(n271), .S0(
        product[18]) );
  HS65_LH_FA1X4 U273 ( .A0(n1402), .B0(n853), .CI(n273), .CO(n272), .S0(
        product[17]) );
  HS65_LH_FA1X4 U274 ( .A0(n1403), .B0(n863), .CI(n274), .CO(n273), .S0(
        product[16]) );
  HS65_LH_FA1X4 U275 ( .A0(n1404), .B0(n873), .CI(n275), .CO(n274), .S0(
        product[15]) );
  HS65_LH_FA1X4 U276 ( .A0(n1405), .B0(n883), .CI(n276), .CO(n275), .S0(
        product[14]) );
  HS65_LH_FA1X4 U277 ( .A0(n1406), .B0(n891), .CI(n277), .CO(n276), .S0(
        product[13]) );
  HS65_LH_FA1X4 U278 ( .A0(n1407), .B0(n899), .CI(n278), .CO(n277), .S0(
        product[12]) );
  HS65_LH_FA1X4 U279 ( .A0(n1408), .B0(n907), .CI(n279), .CO(n278), .S0(
        product[11]) );
  HS65_LH_FA1X4 U280 ( .A0(n1409), .B0(n913), .CI(n280), .CO(n279), .S0(
        product[10]) );
  HS65_LH_FA1X4 U281 ( .A0(n1410), .B0(n919), .CI(n281), .CO(n280), .S0(
        product[9]) );
  HS65_LH_FA1X4 U282 ( .A0(n1411), .B0(n925), .CI(n282), .CO(n281), .S0(
        product[8]) );
  HS65_LH_FA1X4 U283 ( .A0(n1412), .B0(n929), .CI(n283), .CO(n282), .S0(
        product[7]) );
  HS65_LH_FA1X4 U284 ( .A0(n1413), .B0(n933), .CI(n284), .CO(n283), .S0(
        product[6]) );
  HS65_LH_FA1X4 U285 ( .A0(n1414), .B0(n937), .CI(n285), .CO(n284), .S0(
        product[5]) );
  HS65_LH_FA1X4 U286 ( .A0(n1415), .B0(n939), .CI(n286), .CO(n285), .S0(
        product[4]) );
  HS65_LH_FA1X4 U287 ( .A0(n1416), .B0(n941), .CI(n287), .CO(n286), .S0(
        product[3]) );
  HS65_LH_HA1X4 U288 ( .A0(n1417), .B0(n288), .CO(n287), .S0(product[2]) );
  HS65_LH_HA1X4 U289 ( .A0(n1418), .B0(n289), .CO(n288), .S0(product[1]) );
  HS65_LH_HA1X4 U290 ( .A0(n2629), .B0(n1419), .CO(n289), .S0(product[0]) );
  HS65_LH_FA1X4 U293 ( .A0(n297), .B0(n2657), .CI(n1041), .CO(n293), .S0(n294)
         );
  HS65_LH_FA1X4 U294 ( .A0(n1042), .B0(n2658), .CI(n1071), .CO(n295), .S0(n296) );
  HS65_LH_FA1X4 U296 ( .A0(n2658), .B0(n1043), .CI(n1072), .CO(n299), .S0(n300) );
  HS65_LH_FA1X4 U298 ( .A0(n1073), .B0(n304), .CI(n307), .CO(n302), .S0(n303)
         );
  HS65_LH_FA1X4 U299 ( .A0(n309), .B0(n2654), .CI(n1044), .CO(n297), .S0(n304)
         );
  HS65_LH_FA1X4 U300 ( .A0(n1106), .B0(n1074), .CI(n308), .CO(n305), .S0(n306)
         );
  HS65_LH_FA1X4 U301 ( .A0(n1045), .B0(n2663), .CI(n313), .CO(n307), .S0(n308)
         );
  HS65_LH_FA1X4 U303 ( .A0(n314), .B0(n318), .CI(n1107), .CO(n311), .S0(n312)
         );
  HS65_LH_FA1X4 U304 ( .A0(n2663), .B0(n320), .CI(n1075), .CO(n313), .S0(n314)
         );
  HS65_LH_FA1X4 U306 ( .A0(n1108), .B0(n319), .CI(n324), .CO(n316), .S0(n317)
         );
  HS65_LH_FA1X4 U307 ( .A0(n326), .B0(n321), .CI(n1076), .CO(n318), .S0(n319)
         );
  HS65_LH_FA1X4 U308 ( .A0(n328), .B0(n2651), .CI(n1046), .CO(n320), .S0(n321)
         );
  HS65_LH_FA1X4 U309 ( .A0(n1141), .B0(n1109), .CI(n325), .CO(n322), .S0(n323)
         );
  HS65_LH_FA1X4 U310 ( .A0(n327), .B0(n334), .CI(n332), .CO(n324), .S0(n325)
         );
  HS65_LH_FA1X4 U311 ( .A0(n1047), .B0(n2659), .CI(n1077), .CO(n326), .S0(n327) );
  HS65_LH_FA1X4 U313 ( .A0(n333), .B0(n339), .CI(n1142), .CO(n330), .S0(n331)
         );
  HS65_LH_FA1X4 U314 ( .A0(n335), .B0(n341), .CI(n1110), .CO(n332), .S0(n333)
         );
  HS65_LH_FA1X4 U315 ( .A0(n2659), .B0(n1048), .CI(n1078), .CO(n334), .S0(n335) );
  HS65_LH_FA1X4 U317 ( .A0(n1143), .B0(n340), .CI(n346), .CO(n337), .S0(n338)
         );
  HS65_LH_FA1X4 U318 ( .A0(n348), .B0(n342), .CI(n1111), .CO(n339), .S0(n340)
         );
  HS65_LH_FA1X4 U319 ( .A0(n1079), .B0(n343), .CI(n350), .CO(n341), .S0(n342)
         );
  HS65_LH_FA1X4 U320 ( .A0(n352), .B0(n2648), .CI(n1049), .CO(n328), .S0(n343)
         );
  HS65_LH_FA1X4 U321 ( .A0(n1176), .B0(n1144), .CI(n347), .CO(n344), .S0(n345)
         );
  HS65_LH_FA1X4 U322 ( .A0(n349), .B0(n358), .CI(n356), .CO(n346), .S0(n347)
         );
  HS65_LH_FA1X4 U323 ( .A0(n351), .B0(n1080), .CI(n1112), .CO(n348), .S0(n349)
         );
  HS65_LH_FA1X4 U324 ( .A0(n1050), .B0(n2664), .CI(n360), .CO(n350), .S0(n351)
         );
  HS65_LH_FA1X4 U326 ( .A0(n357), .B0(n365), .CI(n1177), .CO(n354), .S0(n355)
         );
  HS65_LH_FA1X4 U327 ( .A0(n359), .B0(n367), .CI(n1145), .CO(n356), .S0(n357)
         );
  HS65_LH_FA1X4 U328 ( .A0(n361), .B0(n369), .CI(n1113), .CO(n358), .S0(n359)
         );
  HS65_LH_FA1X4 U329 ( .A0(n2664), .B0(n371), .CI(n1081), .CO(n360), .S0(n361)
         );
  HS65_LH_FA1X4 U331 ( .A0(n1178), .B0(n366), .CI(n375), .CO(n363), .S0(n364)
         );
  HS65_LH_FA1X4 U332 ( .A0(n377), .B0(n368), .CI(n1146), .CO(n365), .S0(n366)
         );
  HS65_LH_FA1X4 U333 ( .A0(n1114), .B0(n370), .CI(n379), .CO(n367), .S0(n368)
         );
  HS65_LH_FA1X4 U334 ( .A0(n381), .B0(n372), .CI(n1082), .CO(n369), .S0(n370)
         );
  HS65_LH_FA1X4 U335 ( .A0(n383), .B0(n2645), .CI(n1051), .CO(n371), .S0(n372)
         );
  HS65_LH_FA1X4 U336 ( .A0(n1211), .B0(n1179), .CI(n376), .CO(n373), .S0(n374)
         );
  HS65_LH_FA1X4 U337 ( .A0(n378), .B0(n389), .CI(n387), .CO(n375), .S0(n376)
         );
  HS65_LH_FA1X4 U338 ( .A0(n380), .B0(n1115), .CI(n1147), .CO(n377), .S0(n378)
         );
  HS65_LH_FA1X4 U339 ( .A0(n382), .B0(n393), .CI(n391), .CO(n379), .S0(n380)
         );
  HS65_LH_FA1X4 U340 ( .A0(n1052), .B0(n2660), .CI(n1083), .CO(n381), .S0(n382) );
  HS65_LH_FA1X4 U342 ( .A0(n388), .B0(n398), .CI(n1212), .CO(n385), .S0(n386)
         );
  HS65_LH_FA1X4 U343 ( .A0(n390), .B0(n400), .CI(n1180), .CO(n387), .S0(n388)
         );
  HS65_LH_FA1X4 U344 ( .A0(n392), .B0(n402), .CI(n1148), .CO(n389), .S0(n390)
         );
  HS65_LH_FA1X4 U345 ( .A0(n394), .B0(n404), .CI(n1116), .CO(n391), .S0(n392)
         );
  HS65_LH_FA1X4 U346 ( .A0(n2660), .B0(n1053), .CI(n1084), .CO(n393), .S0(n394) );
  HS65_LH_FA1X4 U348 ( .A0(n1213), .B0(n399), .CI(n409), .CO(n396), .S0(n397)
         );
  HS65_LH_FA1X4 U349 ( .A0(n411), .B0(n401), .CI(n1181), .CO(n398), .S0(n399)
         );
  HS65_LH_FA1X4 U350 ( .A0(n1149), .B0(n403), .CI(n413), .CO(n400), .S0(n401)
         );
  HS65_LH_FA1X4 U351 ( .A0(n415), .B0(n405), .CI(n1117), .CO(n402), .S0(n403)
         );
  HS65_LH_FA1X4 U352 ( .A0(n1085), .B0(n406), .CI(n417), .CO(n404), .S0(n405)
         );
  HS65_LH_FA1X4 U353 ( .A0(n419), .B0(n2642), .CI(n1054), .CO(n383), .S0(n406)
         );
  HS65_LH_FA1X4 U354 ( .A0(n1246), .B0(n1214), .CI(n410), .CO(n407), .S0(n408)
         );
  HS65_LH_FA1X4 U355 ( .A0(n412), .B0(n425), .CI(n423), .CO(n409), .S0(n410)
         );
  HS65_LH_FA1X4 U356 ( .A0(n414), .B0(n1150), .CI(n1182), .CO(n411), .S0(n412)
         );
  HS65_LH_FA1X4 U357 ( .A0(n416), .B0(n429), .CI(n427), .CO(n413), .S0(n414)
         );
  HS65_LH_FA1X4 U358 ( .A0(n418), .B0(n1086), .CI(n1118), .CO(n415), .S0(n416)
         );
  HS65_LH_FA1X4 U359 ( .A0(n1055), .B0(n2665), .CI(n431), .CO(n417), .S0(n418)
         );
  HS65_LH_FA1X4 U361 ( .A0(n424), .B0(n436), .CI(n1247), .CO(n421), .S0(n422)
         );
  HS65_LH_FA1X4 U362 ( .A0(n426), .B0(n438), .CI(n1215), .CO(n423), .S0(n424)
         );
  HS65_LH_FA1X4 U363 ( .A0(n428), .B0(n440), .CI(n1183), .CO(n425), .S0(n426)
         );
  HS65_LH_FA1X4 U364 ( .A0(n430), .B0(n442), .CI(n1151), .CO(n427), .S0(n428)
         );
  HS65_LH_FA1X4 U365 ( .A0(n432), .B0(n444), .CI(n1119), .CO(n429), .S0(n430)
         );
  HS65_LH_FA1X4 U366 ( .A0(n2665), .B0(n446), .CI(n1087), .CO(n431), .S0(n432)
         );
  HS65_LH_FA1X4 U368 ( .A0(n1248), .B0(n437), .CI(n450), .CO(n434), .S0(n435)
         );
  HS65_LH_FA1X4 U369 ( .A0(n452), .B0(n439), .CI(n1216), .CO(n436), .S0(n437)
         );
  HS65_LH_FA1X4 U370 ( .A0(n1184), .B0(n441), .CI(n454), .CO(n438), .S0(n439)
         );
  HS65_LH_FA1X4 U371 ( .A0(n456), .B0(n443), .CI(n1152), .CO(n440), .S0(n441)
         );
  HS65_LH_FA1X4 U372 ( .A0(n1120), .B0(n445), .CI(n458), .CO(n442), .S0(n443)
         );
  HS65_LH_FA1X4 U373 ( .A0(n460), .B0(n447), .CI(n1088), .CO(n444), .S0(n445)
         );
  HS65_LH_FA1X4 U374 ( .A0(n462), .B0(n2639), .CI(n1056), .CO(n446), .S0(n447)
         );
  HS65_LH_FA1X4 U375 ( .A0(n1281), .B0(n1249), .CI(n451), .CO(n448), .S0(n449)
         );
  HS65_LH_FA1X4 U376 ( .A0(n453), .B0(n468), .CI(n466), .CO(n450), .S0(n451)
         );
  HS65_LH_FA1X4 U377 ( .A0(n455), .B0(n1185), .CI(n1217), .CO(n452), .S0(n453)
         );
  HS65_LH_FA1X4 U378 ( .A0(n457), .B0(n472), .CI(n470), .CO(n454), .S0(n455)
         );
  HS65_LH_FA1X4 U379 ( .A0(n459), .B0(n1121), .CI(n1153), .CO(n456), .S0(n457)
         );
  HS65_LH_FA1X4 U380 ( .A0(n461), .B0(n476), .CI(n474), .CO(n458), .S0(n459)
         );
  HS65_LH_FA1X4 U381 ( .A0(n1057), .B0(n2661), .CI(n1089), .CO(n460), .S0(n461) );
  HS65_LH_FA1X4 U383 ( .A0(n467), .B0(n481), .CI(n1282), .CO(n464), .S0(n465)
         );
  HS65_LH_FA1X4 U384 ( .A0(n469), .B0(n483), .CI(n1250), .CO(n466), .S0(n467)
         );
  HS65_LH_FA1X4 U385 ( .A0(n471), .B0(n485), .CI(n1218), .CO(n468), .S0(n469)
         );
  HS65_LH_FA1X4 U386 ( .A0(n473), .B0(n487), .CI(n1186), .CO(n470), .S0(n471)
         );
  HS65_LH_FA1X4 U387 ( .A0(n475), .B0(n489), .CI(n1154), .CO(n472), .S0(n473)
         );
  HS65_LH_FA1X4 U388 ( .A0(n477), .B0(n491), .CI(n1122), .CO(n474), .S0(n475)
         );
  HS65_LH_FA1X4 U389 ( .A0(n2661), .B0(n1058), .CI(n1090), .CO(n476), .S0(n477) );
  HS65_LH_FA1X4 U391 ( .A0(n1283), .B0(n482), .CI(n496), .CO(n479), .S0(n480)
         );
  HS65_LH_FA1X4 U392 ( .A0(n498), .B0(n484), .CI(n1251), .CO(n481), .S0(n482)
         );
  HS65_LH_FA1X4 U393 ( .A0(n1219), .B0(n486), .CI(n500), .CO(n483), .S0(n484)
         );
  HS65_LH_FA1X4 U394 ( .A0(n502), .B0(n488), .CI(n1187), .CO(n485), .S0(n486)
         );
  HS65_LH_FA1X4 U395 ( .A0(n1155), .B0(n490), .CI(n504), .CO(n487), .S0(n488)
         );
  HS65_LH_FA1X4 U396 ( .A0(n506), .B0(n492), .CI(n1123), .CO(n489), .S0(n490)
         );
  HS65_LH_FA1X4 U397 ( .A0(n1091), .B0(n493), .CI(n508), .CO(n491), .S0(n492)
         );
  HS65_LH_FA1X4 U398 ( .A0(n510), .B0(n2636), .CI(n1059), .CO(n462), .S0(n493)
         );
  HS65_LH_FA1X4 U399 ( .A0(n1316), .B0(n1284), .CI(n497), .CO(n494), .S0(n495)
         );
  HS65_LH_FA1X4 U400 ( .A0(n499), .B0(n516), .CI(n514), .CO(n496), .S0(n497)
         );
  HS65_LH_FA1X4 U401 ( .A0(n501), .B0(n1220), .CI(n1252), .CO(n498), .S0(n499)
         );
  HS65_LH_FA1X4 U402 ( .A0(n503), .B0(n520), .CI(n518), .CO(n500), .S0(n501)
         );
  HS65_LH_FA1X4 U403 ( .A0(n505), .B0(n1156), .CI(n1188), .CO(n502), .S0(n503)
         );
  HS65_LH_FA1X4 U404 ( .A0(n507), .B0(n524), .CI(n522), .CO(n504), .S0(n505)
         );
  HS65_LH_FA1X4 U405 ( .A0(n509), .B0(n1092), .CI(n1124), .CO(n506), .S0(n507)
         );
  HS65_LH_FA1X4 U406 ( .A0(n1060), .B0(n2662), .CI(n526), .CO(n508), .S0(n509)
         );
  HS65_LH_FA1X4 U408 ( .A0(n515), .B0(n531), .CI(n1317), .CO(n512), .S0(n513)
         );
  HS65_LH_FA1X4 U409 ( .A0(n517), .B0(n533), .CI(n1285), .CO(n514), .S0(n515)
         );
  HS65_LH_FA1X4 U410 ( .A0(n519), .B0(n535), .CI(n1253), .CO(n516), .S0(n517)
         );
  HS65_LH_FA1X4 U411 ( .A0(n521), .B0(n537), .CI(n1221), .CO(n518), .S0(n519)
         );
  HS65_LH_FA1X4 U412 ( .A0(n523), .B0(n539), .CI(n1189), .CO(n520), .S0(n521)
         );
  HS65_LH_FA1X4 U413 ( .A0(n525), .B0(n541), .CI(n1157), .CO(n522), .S0(n523)
         );
  HS65_LH_FA1X4 U414 ( .A0(n527), .B0(n543), .CI(n1125), .CO(n524), .S0(n525)
         );
  HS65_LH_FA1X4 U415 ( .A0(n2662), .B0(n1061), .CI(n1093), .CO(n526), .S0(n527) );
  HS65_LH_FA1X4 U417 ( .A0(n1318), .B0(n532), .CI(n548), .CO(n529), .S0(n530)
         );
  HS65_LH_FA1X4 U418 ( .A0(n550), .B0(n534), .CI(n1286), .CO(n531), .S0(n532)
         );
  HS65_LH_FA1X4 U419 ( .A0(n1254), .B0(n536), .CI(n552), .CO(n533), .S0(n534)
         );
  HS65_LH_FA1X4 U420 ( .A0(n554), .B0(n538), .CI(n1222), .CO(n535), .S0(n536)
         );
  HS65_LH_FA1X4 U421 ( .A0(n1190), .B0(n540), .CI(n556), .CO(n537), .S0(n538)
         );
  HS65_LH_FA1X4 U422 ( .A0(n1158), .B0(n542), .CI(n558), .CO(n539), .S0(n540)
         );
  HS65_LH_FA1X4 U423 ( .A0(n1126), .B0(n544), .CI(n560), .CO(n541), .S0(n542)
         );
  HS65_LH_FA1X4 U424 ( .A0(n562), .B0(n545), .CI(n1094), .CO(n543), .S0(n544)
         );
  HS65_LH_FA1X4 U425 ( .A0(n2633), .B0(n2630), .CI(n1062), .CO(n510), .S0(n545) );
  HS65_LH_FA1X4 U426 ( .A0(n1351), .B0(n1319), .CI(n549), .CO(n546), .S0(n547)
         );
  HS65_LH_FA1X4 U427 ( .A0(n551), .B0(n1287), .CI(n566), .CO(n548), .S0(n549)
         );
  HS65_LH_FA1X4 U428 ( .A0(n553), .B0(n1255), .CI(n568), .CO(n550), .S0(n551)
         );
  HS65_LH_FA1X4 U429 ( .A0(n555), .B0(n572), .CI(n570), .CO(n552), .S0(n553)
         );
  HS65_LH_FA1X4 U430 ( .A0(n557), .B0(n1191), .CI(n1223), .CO(n554), .S0(n555)
         );
  HS65_LH_FA1X4 U431 ( .A0(n559), .B0(n576), .CI(n574), .CO(n556), .S0(n557)
         );
  HS65_LH_FA1X4 U432 ( .A0(n561), .B0(n1127), .CI(n1159), .CO(n558), .S0(n559)
         );
  HS65_LH_FA1X4 U433 ( .A0(n563), .B0(n1095), .CI(n578), .CO(n560), .S0(n561)
         );
  HS65_LH_FA1X4 U434 ( .A0(n1063), .B0(n2628), .CI(n580), .CO(n562), .S0(n563)
         );
  HS65_LH_FA1X4 U435 ( .A0(n567), .B0(n1320), .CI(n1352), .CO(n564), .S0(n565)
         );
  HS65_LH_FA1X4 U436 ( .A0(n569), .B0(n1288), .CI(n584), .CO(n566), .S0(n567)
         );
  HS65_LH_FA1X4 U437 ( .A0(n571), .B0(n1256), .CI(n586), .CO(n568), .S0(n569)
         );
  HS65_LH_FA1X4 U438 ( .A0(n573), .B0(n590), .CI(n588), .CO(n570), .S0(n571)
         );
  HS65_LH_FA1X4 U439 ( .A0(n575), .B0(n1192), .CI(n1224), .CO(n572), .S0(n573)
         );
  HS65_LH_FA1X4 U440 ( .A0(n577), .B0(n594), .CI(n592), .CO(n574), .S0(n575)
         );
  HS65_LH_FA1X4 U441 ( .A0(n579), .B0(n1128), .CI(n1160), .CO(n576), .S0(n577)
         );
  HS65_LH_FA1X4 U442 ( .A0(n581), .B0(n1096), .CI(n596), .CO(n578), .S0(n579)
         );
  HS65_LH_FA1X4 U443 ( .A0(n1064), .B0(n2628), .CI(n598), .CO(n580), .S0(n581)
         );
  HS65_LH_FA1X4 U444 ( .A0(n585), .B0(n602), .CI(n1353), .CO(n582), .S0(n583)
         );
  HS65_LH_FA1X4 U445 ( .A0(n587), .B0(n604), .CI(n1321), .CO(n584), .S0(n585)
         );
  HS65_LH_FA1X4 U446 ( .A0(n589), .B0(n606), .CI(n1289), .CO(n586), .S0(n587)
         );
  HS65_LH_FA1X4 U447 ( .A0(n591), .B0(n608), .CI(n1257), .CO(n588), .S0(n589)
         );
  HS65_LH_FA1X4 U448 ( .A0(n593), .B0(n610), .CI(n1225), .CO(n590), .S0(n591)
         );
  HS65_LH_FA1X4 U449 ( .A0(n595), .B0(n612), .CI(n1193), .CO(n592), .S0(n593)
         );
  HS65_LH_FA1X4 U450 ( .A0(n597), .B0(n614), .CI(n1161), .CO(n594), .S0(n595)
         );
  HS65_LH_FA1X4 U451 ( .A0(n599), .B0(n616), .CI(n1129), .CO(n596), .S0(n597)
         );
  HS65_LH_FA1X4 U452 ( .A0(n1065), .B0(n2628), .CI(n1097), .CO(n598), .S0(n599) );
  HS65_LH_FA1X4 U453 ( .A0(n1354), .B0(n603), .CI(n618), .CO(n600), .S0(n601)
         );
  HS65_LH_FA1X4 U454 ( .A0(n1322), .B0(n605), .CI(n620), .CO(n602), .S0(n603)
         );
  HS65_LH_FA1X4 U455 ( .A0(n1290), .B0(n607), .CI(n622), .CO(n604), .S0(n605)
         );
  HS65_LH_FA1X4 U456 ( .A0(n1258), .B0(n609), .CI(n624), .CO(n606), .S0(n607)
         );
  HS65_LH_FA1X4 U457 ( .A0(n1226), .B0(n611), .CI(n626), .CO(n608), .S0(n609)
         );
  HS65_LH_FA1X4 U458 ( .A0(n1194), .B0(n613), .CI(n628), .CO(n610), .S0(n611)
         );
  HS65_LH_FA1X4 U459 ( .A0(n1162), .B0(n615), .CI(n630), .CO(n612), .S0(n613)
         );
  HS65_LH_FA1X4 U460 ( .A0(n1130), .B0(n617), .CI(n632), .CO(n614), .S0(n615)
         );
  HS65_LH_FA1X4 U461 ( .A0(n1098), .B0(n1066), .CI(n634), .CO(n616), .S0(n617)
         );
  HS65_LH_FA1X4 U462 ( .A0(n1355), .B0(n621), .CI(n636), .CO(n618), .S0(n619)
         );
  HS65_LH_FA1X4 U463 ( .A0(n1323), .B0(n623), .CI(n638), .CO(n620), .S0(n621)
         );
  HS65_LH_FA1X4 U464 ( .A0(n1291), .B0(n625), .CI(n640), .CO(n622), .S0(n623)
         );
  HS65_LH_FA1X4 U465 ( .A0(n1259), .B0(n627), .CI(n642), .CO(n624), .S0(n625)
         );
  HS65_LH_FA1X4 U466 ( .A0(n1227), .B0(n629), .CI(n644), .CO(n626), .S0(n627)
         );
  HS65_LH_FA1X4 U467 ( .A0(n1195), .B0(n631), .CI(n646), .CO(n628), .S0(n629)
         );
  HS65_LH_FA1X4 U468 ( .A0(n1163), .B0(n633), .CI(n648), .CO(n630), .S0(n631)
         );
  HS65_LH_FA1X4 U469 ( .A0(n1131), .B0(n635), .CI(n650), .CO(n632), .S0(n633)
         );
  HS65_LH_FA1X4 U470 ( .A0(n1099), .B0(n1067), .CI(n652), .CO(n634), .S0(n635)
         );
  HS65_LH_FA1X4 U471 ( .A0(n1356), .B0(n639), .CI(n654), .CO(n636), .S0(n637)
         );
  HS65_LH_FA1X4 U472 ( .A0(n1324), .B0(n641), .CI(n656), .CO(n638), .S0(n639)
         );
  HS65_LH_FA1X4 U473 ( .A0(n1292), .B0(n643), .CI(n658), .CO(n640), .S0(n641)
         );
  HS65_LH_FA1X4 U474 ( .A0(n1260), .B0(n645), .CI(n660), .CO(n642), .S0(n643)
         );
  HS65_LH_FA1X4 U475 ( .A0(n1228), .B0(n647), .CI(n662), .CO(n644), .S0(n645)
         );
  HS65_LH_FA1X4 U476 ( .A0(n1196), .B0(n649), .CI(n664), .CO(n646), .S0(n647)
         );
  HS65_LH_FA1X4 U477 ( .A0(n1164), .B0(n651), .CI(n666), .CO(n648), .S0(n649)
         );
  HS65_LH_FA1X4 U478 ( .A0(n1132), .B0(n653), .CI(n668), .CO(n650), .S0(n651)
         );
  HS65_LH_FA1X4 U479 ( .A0(n1100), .B0(n1068), .CI(n670), .CO(n652), .S0(n653)
         );
  HS65_LH_FA1X4 U480 ( .A0(n1357), .B0(n657), .CI(n672), .CO(n654), .S0(n655)
         );
  HS65_LH_FA1X4 U481 ( .A0(n1325), .B0(n659), .CI(n674), .CO(n656), .S0(n657)
         );
  HS65_LH_FA1X4 U482 ( .A0(n1293), .B0(n661), .CI(n676), .CO(n658), .S0(n659)
         );
  HS65_LH_FA1X4 U483 ( .A0(n1261), .B0(n663), .CI(n678), .CO(n660), .S0(n661)
         );
  HS65_LH_FA1X4 U484 ( .A0(n1229), .B0(n665), .CI(n680), .CO(n662), .S0(n663)
         );
  HS65_LH_FA1X4 U485 ( .A0(n1197), .B0(n667), .CI(n682), .CO(n664), .S0(n665)
         );
  HS65_LH_FA1X4 U486 ( .A0(n1165), .B0(n669), .CI(n684), .CO(n666), .S0(n667)
         );
  HS65_LH_FA1X4 U487 ( .A0(n1133), .B0(n671), .CI(n686), .CO(n668), .S0(n669)
         );
  HS65_LH_FA1X4 U488 ( .A0(n1101), .B0(n1069), .CI(n688), .CO(n670), .S0(n671)
         );
  HS65_LH_FA1X4 U489 ( .A0(n1358), .B0(n675), .CI(n690), .CO(n672), .S0(n673)
         );
  HS65_LH_FA1X4 U490 ( .A0(n1326), .B0(n677), .CI(n692), .CO(n674), .S0(n675)
         );
  HS65_LH_FA1X4 U491 ( .A0(n1294), .B0(n679), .CI(n694), .CO(n676), .S0(n677)
         );
  HS65_LH_FA1X4 U492 ( .A0(n1262), .B0(n681), .CI(n696), .CO(n678), .S0(n679)
         );
  HS65_LH_FA1X4 U493 ( .A0(n1230), .B0(n683), .CI(n698), .CO(n680), .S0(n681)
         );
  HS65_LH_FA1X4 U494 ( .A0(n1198), .B0(n685), .CI(n700), .CO(n682), .S0(n683)
         );
  HS65_LH_FA1X4 U495 ( .A0(n1166), .B0(n687), .CI(n702), .CO(n684), .S0(n685)
         );
  HS65_LH_FA1X4 U496 ( .A0(n1134), .B0(n689), .CI(n704), .CO(n686), .S0(n687)
         );
  HS65_LH_HA1X4 U497 ( .A0(n1102), .B0(n706), .CO(n688), .S0(n689) );
  HS65_LH_FA1X4 U498 ( .A0(n1359), .B0(n693), .CI(n708), .CO(n690), .S0(n691)
         );
  HS65_LH_FA1X4 U499 ( .A0(n1327), .B0(n695), .CI(n710), .CO(n692), .S0(n693)
         );
  HS65_LH_FA1X4 U500 ( .A0(n1295), .B0(n697), .CI(n712), .CO(n694), .S0(n695)
         );
  HS65_LH_FA1X4 U501 ( .A0(n1263), .B0(n699), .CI(n714), .CO(n696), .S0(n697)
         );
  HS65_LH_FA1X4 U502 ( .A0(n1231), .B0(n701), .CI(n716), .CO(n698), .S0(n699)
         );
  HS65_LH_FA1X4 U503 ( .A0(n1199), .B0(n703), .CI(n718), .CO(n700), .S0(n701)
         );
  HS65_LH_FA1X4 U504 ( .A0(n1167), .B0(n705), .CI(n720), .CO(n702), .S0(n703)
         );
  HS65_LH_FA1X4 U505 ( .A0(n1135), .B0(n707), .CI(n722), .CO(n704), .S0(n705)
         );
  HS65_LH_HA1X4 U506 ( .A0(n1103), .B0(n724), .CO(n706), .S0(n707) );
  HS65_LH_FA1X4 U507 ( .A0(n1360), .B0(n711), .CI(n726), .CO(n708), .S0(n709)
         );
  HS65_LH_FA1X4 U508 ( .A0(n1328), .B0(n713), .CI(n728), .CO(n710), .S0(n711)
         );
  HS65_LH_FA1X4 U509 ( .A0(n1296), .B0(n715), .CI(n730), .CO(n712), .S0(n713)
         );
  HS65_LH_FA1X4 U510 ( .A0(n1264), .B0(n717), .CI(n732), .CO(n714), .S0(n715)
         );
  HS65_LH_FA1X4 U511 ( .A0(n1232), .B0(n719), .CI(n734), .CO(n716), .S0(n717)
         );
  HS65_LH_FA1X4 U512 ( .A0(n1200), .B0(n721), .CI(n736), .CO(n718), .S0(n719)
         );
  HS65_LH_FA1X4 U513 ( .A0(n1168), .B0(n723), .CI(n738), .CO(n720), .S0(n721)
         );
  HS65_LH_FA1X4 U514 ( .A0(n1136), .B0(n725), .CI(n740), .CO(n722), .S0(n723)
         );
  HS65_LH_HA1X4 U515 ( .A0(n2656), .B0(n1104), .CO(n724), .S0(n725) );
  HS65_LH_FA1X4 U516 ( .A0(n1361), .B0(n729), .CI(n742), .CO(n726), .S0(n727)
         );
  HS65_LH_FA1X4 U517 ( .A0(n1329), .B0(n731), .CI(n744), .CO(n728), .S0(n729)
         );
  HS65_LH_FA1X4 U518 ( .A0(n1297), .B0(n733), .CI(n746), .CO(n730), .S0(n731)
         );
  HS65_LH_FA1X4 U519 ( .A0(n1265), .B0(n735), .CI(n748), .CO(n732), .S0(n733)
         );
  HS65_LH_FA1X4 U520 ( .A0(n1233), .B0(n737), .CI(n750), .CO(n734), .S0(n735)
         );
  HS65_LH_FA1X4 U521 ( .A0(n1201), .B0(n739), .CI(n752), .CO(n736), .S0(n737)
         );
  HS65_LH_FA1X4 U522 ( .A0(n1169), .B0(n741), .CI(n754), .CO(n738), .S0(n739)
         );
  HS65_LH_HA1X4 U523 ( .A0(n1137), .B0(n756), .CO(n740), .S0(n741) );
  HS65_LH_FA1X4 U524 ( .A0(n1362), .B0(n745), .CI(n758), .CO(n742), .S0(n743)
         );
  HS65_LH_FA1X4 U525 ( .A0(n1330), .B0(n747), .CI(n760), .CO(n744), .S0(n745)
         );
  HS65_LH_FA1X4 U526 ( .A0(n1298), .B0(n749), .CI(n762), .CO(n746), .S0(n747)
         );
  HS65_LH_FA1X4 U527 ( .A0(n1266), .B0(n751), .CI(n764), .CO(n748), .S0(n749)
         );
  HS65_LH_FA1X4 U528 ( .A0(n1234), .B0(n753), .CI(n766), .CO(n750), .S0(n751)
         );
  HS65_LH_FA1X4 U529 ( .A0(n1202), .B0(n755), .CI(n768), .CO(n752), .S0(n753)
         );
  HS65_LH_FA1X4 U530 ( .A0(n1170), .B0(n757), .CI(n770), .CO(n754), .S0(n755)
         );
  HS65_LH_HA1X4 U531 ( .A0(n1138), .B0(n772), .CO(n756), .S0(n757) );
  HS65_LH_FA1X4 U532 ( .A0(n1363), .B0(n761), .CI(n774), .CO(n758), .S0(n759)
         );
  HS65_LH_FA1X4 U533 ( .A0(n1331), .B0(n763), .CI(n776), .CO(n760), .S0(n761)
         );
  HS65_LH_FA1X4 U534 ( .A0(n1299), .B0(n765), .CI(n778), .CO(n762), .S0(n763)
         );
  HS65_LH_FA1X4 U535 ( .A0(n1267), .B0(n767), .CI(n780), .CO(n764), .S0(n765)
         );
  HS65_LH_FA1X4 U536 ( .A0(n1235), .B0(n769), .CI(n782), .CO(n766), .S0(n767)
         );
  HS65_LH_FA1X4 U537 ( .A0(n1203), .B0(n771), .CI(n784), .CO(n768), .S0(n769)
         );
  HS65_LH_FA1X4 U538 ( .A0(n1171), .B0(n773), .CI(n786), .CO(n770), .S0(n771)
         );
  HS65_LH_HA1X4 U539 ( .A0(n2653), .B0(n1139), .CO(n772), .S0(n773) );
  HS65_LH_FA1X4 U540 ( .A0(n1364), .B0(n777), .CI(n788), .CO(n774), .S0(n775)
         );
  HS65_LH_FA1X4 U541 ( .A0(n1332), .B0(n779), .CI(n790), .CO(n776), .S0(n777)
         );
  HS65_LH_FA1X4 U542 ( .A0(n1300), .B0(n781), .CI(n792), .CO(n778), .S0(n779)
         );
  HS65_LH_FA1X4 U543 ( .A0(n1268), .B0(n783), .CI(n794), .CO(n780), .S0(n781)
         );
  HS65_LH_FA1X4 U544 ( .A0(n1236), .B0(n785), .CI(n796), .CO(n782), .S0(n783)
         );
  HS65_LH_FA1X4 U545 ( .A0(n1204), .B0(n787), .CI(n798), .CO(n784), .S0(n785)
         );
  HS65_LH_HA1X4 U546 ( .A0(n1172), .B0(n800), .CO(n786), .S0(n787) );
  HS65_LH_FA1X4 U547 ( .A0(n1365), .B0(n791), .CI(n802), .CO(n788), .S0(n789)
         );
  HS65_LH_FA1X4 U548 ( .A0(n1333), .B0(n793), .CI(n804), .CO(n790), .S0(n791)
         );
  HS65_LH_FA1X4 U549 ( .A0(n1301), .B0(n795), .CI(n806), .CO(n792), .S0(n793)
         );
  HS65_LH_FA1X4 U550 ( .A0(n1269), .B0(n797), .CI(n808), .CO(n794), .S0(n795)
         );
  HS65_LH_FA1X4 U551 ( .A0(n1237), .B0(n799), .CI(n810), .CO(n796), .S0(n797)
         );
  HS65_LH_FA1X4 U552 ( .A0(n1205), .B0(n801), .CI(n812), .CO(n798), .S0(n799)
         );
  HS65_LH_HA1X4 U553 ( .A0(n1173), .B0(n814), .CO(n800), .S0(n801) );
  HS65_LH_FA1X4 U554 ( .A0(n1366), .B0(n805), .CI(n816), .CO(n802), .S0(n803)
         );
  HS65_LH_FA1X4 U555 ( .A0(n1334), .B0(n807), .CI(n818), .CO(n804), .S0(n805)
         );
  HS65_LH_FA1X4 U556 ( .A0(n1302), .B0(n809), .CI(n820), .CO(n806), .S0(n807)
         );
  HS65_LH_FA1X4 U557 ( .A0(n1270), .B0(n811), .CI(n822), .CO(n808), .S0(n809)
         );
  HS65_LH_FA1X4 U558 ( .A0(n1238), .B0(n813), .CI(n824), .CO(n810), .S0(n811)
         );
  HS65_LH_FA1X4 U559 ( .A0(n1206), .B0(n815), .CI(n826), .CO(n812), .S0(n813)
         );
  HS65_LH_HA1X4 U560 ( .A0(n2650), .B0(n1174), .CO(n814), .S0(n815) );
  HS65_LH_FA1X4 U561 ( .A0(n1367), .B0(n819), .CI(n828), .CO(n816), .S0(n817)
         );
  HS65_LH_FA1X4 U562 ( .A0(n1335), .B0(n821), .CI(n830), .CO(n818), .S0(n819)
         );
  HS65_LH_FA1X4 U563 ( .A0(n1303), .B0(n823), .CI(n832), .CO(n820), .S0(n821)
         );
  HS65_LH_FA1X4 U564 ( .A0(n1271), .B0(n825), .CI(n834), .CO(n822), .S0(n823)
         );
  HS65_LH_FA1X4 U565 ( .A0(n1239), .B0(n827), .CI(n836), .CO(n824), .S0(n825)
         );
  HS65_LH_HA1X4 U566 ( .A0(n1207), .B0(n838), .CO(n826), .S0(n827) );
  HS65_LH_FA1X4 U567 ( .A0(n1368), .B0(n831), .CI(n840), .CO(n828), .S0(n829)
         );
  HS65_LH_FA1X4 U568 ( .A0(n1336), .B0(n833), .CI(n842), .CO(n830), .S0(n831)
         );
  HS65_LH_FA1X4 U569 ( .A0(n1304), .B0(n835), .CI(n844), .CO(n832), .S0(n833)
         );
  HS65_LH_FA1X4 U570 ( .A0(n1272), .B0(n837), .CI(n846), .CO(n834), .S0(n835)
         );
  HS65_LH_FA1X4 U571 ( .A0(n1240), .B0(n839), .CI(n848), .CO(n836), .S0(n837)
         );
  HS65_LH_HA1X4 U572 ( .A0(n1208), .B0(n850), .CO(n838), .S0(n839) );
  HS65_LH_FA1X4 U573 ( .A0(n1369), .B0(n843), .CI(n852), .CO(n840), .S0(n841)
         );
  HS65_LH_FA1X4 U574 ( .A0(n1337), .B0(n845), .CI(n854), .CO(n842), .S0(n843)
         );
  HS65_LH_FA1X4 U575 ( .A0(n1305), .B0(n847), .CI(n856), .CO(n844), .S0(n845)
         );
  HS65_LH_FA1X4 U576 ( .A0(n1273), .B0(n849), .CI(n858), .CO(n846), .S0(n847)
         );
  HS65_LH_FA1X4 U577 ( .A0(n1241), .B0(n851), .CI(n860), .CO(n848), .S0(n849)
         );
  HS65_LH_HA1X4 U578 ( .A0(n2647), .B0(n1209), .CO(n850), .S0(n851) );
  HS65_LH_FA1X4 U579 ( .A0(n1370), .B0(n855), .CI(n862), .CO(n852), .S0(n853)
         );
  HS65_LH_FA1X4 U580 ( .A0(n1338), .B0(n857), .CI(n864), .CO(n854), .S0(n855)
         );
  HS65_LH_FA1X4 U581 ( .A0(n1306), .B0(n859), .CI(n866), .CO(n856), .S0(n857)
         );
  HS65_LH_FA1X4 U582 ( .A0(n1274), .B0(n861), .CI(n868), .CO(n858), .S0(n859)
         );
  HS65_LH_HA1X4 U583 ( .A0(n1242), .B0(n870), .CO(n860), .S0(n861) );
  HS65_LH_FA1X4 U584 ( .A0(n1371), .B0(n865), .CI(n872), .CO(n862), .S0(n863)
         );
  HS65_LH_FA1X4 U585 ( .A0(n1339), .B0(n867), .CI(n874), .CO(n864), .S0(n865)
         );
  HS65_LH_FA1X4 U586 ( .A0(n1307), .B0(n869), .CI(n876), .CO(n866), .S0(n867)
         );
  HS65_LH_FA1X4 U587 ( .A0(n1275), .B0(n871), .CI(n878), .CO(n868), .S0(n869)
         );
  HS65_LH_HA1X4 U588 ( .A0(n1243), .B0(n880), .CO(n870), .S0(n871) );
  HS65_LH_FA1X4 U589 ( .A0(n1372), .B0(n875), .CI(n882), .CO(n872), .S0(n873)
         );
  HS65_LH_FA1X4 U590 ( .A0(n1340), .B0(n877), .CI(n884), .CO(n874), .S0(n875)
         );
  HS65_LH_FA1X4 U591 ( .A0(n1308), .B0(n879), .CI(n886), .CO(n876), .S0(n877)
         );
  HS65_LH_FA1X4 U592 ( .A0(n1276), .B0(n881), .CI(n888), .CO(n878), .S0(n879)
         );
  HS65_LH_HA1X4 U593 ( .A0(n2644), .B0(n1244), .CO(n880), .S0(n881) );
  HS65_LH_FA1X4 U594 ( .A0(n1373), .B0(n885), .CI(n890), .CO(n882), .S0(n883)
         );
  HS65_LH_FA1X4 U595 ( .A0(n1341), .B0(n887), .CI(n892), .CO(n884), .S0(n885)
         );
  HS65_LH_FA1X4 U596 ( .A0(n1309), .B0(n889), .CI(n894), .CO(n886), .S0(n887)
         );
  HS65_LH_HA1X4 U597 ( .A0(n1277), .B0(n896), .CO(n888), .S0(n889) );
  HS65_LH_FA1X4 U598 ( .A0(n1374), .B0(n893), .CI(n898), .CO(n890), .S0(n891)
         );
  HS65_LH_FA1X4 U599 ( .A0(n1342), .B0(n895), .CI(n900), .CO(n892), .S0(n893)
         );
  HS65_LH_FA1X4 U600 ( .A0(n1310), .B0(n897), .CI(n902), .CO(n894), .S0(n895)
         );
  HS65_LH_HA1X4 U601 ( .A0(n1278), .B0(n904), .CO(n896), .S0(n897) );
  HS65_LH_FA1X4 U602 ( .A0(n1375), .B0(n901), .CI(n906), .CO(n898), .S0(n899)
         );
  HS65_LH_FA1X4 U603 ( .A0(n1343), .B0(n903), .CI(n908), .CO(n900), .S0(n901)
         );
  HS65_LH_FA1X4 U604 ( .A0(n1311), .B0(n905), .CI(n910), .CO(n902), .S0(n903)
         );
  HS65_LH_HA1X4 U605 ( .A0(n2641), .B0(n1279), .CO(n904), .S0(n905) );
  HS65_LH_FA1X4 U606 ( .A0(n1376), .B0(n909), .CI(n912), .CO(n906), .S0(n907)
         );
  HS65_LH_FA1X4 U607 ( .A0(n1344), .B0(n911), .CI(n914), .CO(n908), .S0(n909)
         );
  HS65_LH_HA1X4 U608 ( .A0(n1312), .B0(n916), .CO(n910), .S0(n911) );
  HS65_LH_FA1X4 U609 ( .A0(n1377), .B0(n915), .CI(n918), .CO(n912), .S0(n913)
         );
  HS65_LH_FA1X4 U610 ( .A0(n1345), .B0(n917), .CI(n920), .CO(n914), .S0(n915)
         );
  HS65_LH_HA1X4 U611 ( .A0(n1313), .B0(n922), .CO(n916), .S0(n917) );
  HS65_LH_FA1X4 U612 ( .A0(n1378), .B0(n921), .CI(n924), .CO(n918), .S0(n919)
         );
  HS65_LH_FA1X4 U613 ( .A0(n1346), .B0(n923), .CI(n926), .CO(n920), .S0(n921)
         );
  HS65_LH_HA1X4 U614 ( .A0(n2638), .B0(n1314), .CO(n922), .S0(n923) );
  HS65_LH_FA1X4 U615 ( .A0(n1379), .B0(n927), .CI(n928), .CO(n924), .S0(n925)
         );
  HS65_LH_HA1X4 U616 ( .A0(n1347), .B0(n930), .CO(n926), .S0(n927) );
  HS65_LH_FA1X4 U617 ( .A0(n1380), .B0(n931), .CI(n932), .CO(n928), .S0(n929)
         );
  HS65_LH_HA1X4 U618 ( .A0(n1348), .B0(n934), .CO(n930), .S0(n931) );
  HS65_LH_FA1X4 U619 ( .A0(n1381), .B0(n935), .CI(n936), .CO(n932), .S0(n933)
         );
  HS65_LH_HA1X4 U620 ( .A0(n2635), .B0(n1349), .CO(n934), .S0(n935) );
  HS65_LH_HA1X4 U621 ( .A0(n1382), .B0(n938), .CO(n936), .S0(n937) );
  HS65_LH_HA1X4 U622 ( .A0(n1383), .B0(n940), .CO(n938), .S0(n939) );
  HS65_LH_HA1X4 U623 ( .A0(n2632), .B0(n1384), .CO(n940), .S0(n941) );
  HS65_LH_HA1X4 U1907 ( .A0(n2626), .B0(n975), .CO(n1006), .S0(n1007) );
  HS65_LH_FA1X4 U1908 ( .A0(n2624), .B0(n2626), .CI(n976), .CO(n975), .S0(
        n1008) );
  HS65_LH_FA1X4 U1909 ( .A0(n2622), .B0(n2624), .CI(n977), .CO(n976), .S0(
        n1009) );
  HS65_LH_FA1X4 U1910 ( .A0(n2620), .B0(n2622), .CI(n978), .CO(n977), .S0(
        n1010) );
  HS65_LH_FA1X4 U1911 ( .A0(n2618), .B0(n2620), .CI(n979), .CO(n978), .S0(
        n1011) );
  HS65_LH_FA1X4 U1912 ( .A0(n2616), .B0(n2618), .CI(n980), .CO(n979), .S0(
        n1012) );
  HS65_LH_FA1X4 U1913 ( .A0(n2614), .B0(n2616), .CI(n981), .CO(n980), .S0(
        n1013) );
  HS65_LH_FA1X4 U1914 ( .A0(n2612), .B0(n2614), .CI(n982), .CO(n981), .S0(
        n1014) );
  HS65_LH_FA1X4 U1915 ( .A0(n2610), .B0(n2612), .CI(n983), .CO(n982), .S0(
        n1015) );
  HS65_LH_FA1X4 U1916 ( .A0(n2608), .B0(n2610), .CI(n984), .CO(n983), .S0(
        n1016) );
  HS65_LH_FA1X4 U1917 ( .A0(n2606), .B0(n2608), .CI(n985), .CO(n984), .S0(
        n1017) );
  HS65_LH_FA1X4 U1918 ( .A0(n2604), .B0(n2606), .CI(n986), .CO(n985), .S0(
        n1018) );
  HS65_LH_FA1X4 U1919 ( .A0(n2602), .B0(n2604), .CI(n987), .CO(n986), .S0(
        n1019) );
  HS65_LH_FA1X4 U1920 ( .A0(n2600), .B0(n2602), .CI(n988), .CO(n987), .S0(
        n1020) );
  HS65_LH_FA1X4 U1921 ( .A0(n2598), .B0(n2600), .CI(n989), .CO(n988), .S0(
        n1021) );
  HS65_LH_FA1X4 U1922 ( .A0(n2596), .B0(n2598), .CI(n990), .CO(n989), .S0(
        n1022) );
  HS65_LH_FA1X4 U1923 ( .A0(n2594), .B0(n2596), .CI(n991), .CO(n990), .S0(
        n1023) );
  HS65_LH_FA1X4 U1924 ( .A0(n2592), .B0(n2594), .CI(n992), .CO(n991), .S0(
        n1024) );
  HS65_LH_FA1X4 U1925 ( .A0(n2590), .B0(n2592), .CI(n993), .CO(n992), .S0(
        n1025) );
  HS65_LH_FA1X4 U1926 ( .A0(n2588), .B0(n2590), .CI(n994), .CO(n993), .S0(
        n1026) );
  HS65_LH_FA1X4 U1927 ( .A0(n2586), .B0(n2588), .CI(n995), .CO(n994), .S0(
        n1027) );
  HS65_LH_FA1X4 U1928 ( .A0(n2584), .B0(n2586), .CI(n996), .CO(n995), .S0(
        n1028) );
  HS65_LH_FA1X4 U1929 ( .A0(n2582), .B0(n2584), .CI(n997), .CO(n996), .S0(
        n1029) );
  HS65_LH_FA1X4 U1930 ( .A0(n2580), .B0(n2582), .CI(n998), .CO(n997), .S0(
        n1030) );
  HS65_LH_FA1X4 U1931 ( .A0(n2578), .B0(n2580), .CI(n999), .CO(n998), .S0(
        n1031) );
  HS65_LH_FA1X4 U1932 ( .A0(n2576), .B0(n2578), .CI(n1000), .CO(n999), .S0(
        n1032) );
  HS65_LH_FA1X4 U1933 ( .A0(n2574), .B0(n2576), .CI(n1001), .CO(n1000), .S0(
        n1033) );
  HS65_LH_FA1X4 U1934 ( .A0(n2572), .B0(n2574), .CI(n1002), .CO(n1001), .S0(
        n1034) );
  HS65_LH_FA1X4 U1935 ( .A0(n2570), .B0(n2572), .CI(n1003), .CO(n1002), .S0(
        n1035) );
  HS65_LH_FA1X4 U1936 ( .A0(n2568), .B0(n2570), .CI(n1004), .CO(n1003), .S0(
        n1036) );
  HS65_LH_FA1X4 U1937 ( .A0(n2566), .B0(n2568), .CI(n1005), .CO(n1004), .S0(
        n1037) );
  HS65_LH_IVX9 U1941 ( .A(n7), .Z(n2630) );
  HS65_LH_IVX9 U1942 ( .A(n1007), .Z(n2667) );
  HS65_LH_IVX9 U1943 ( .A(n2630), .Z(n2628) );
  HS65_LH_IVX9 U1944 ( .A(n2630), .Z(n2629) );
  HS65_LH_BFX9 U1945 ( .A(n2668), .Z(n2422) );
  HS65_LH_BFX9 U1946 ( .A(n2445), .Z(n2446) );
  HS65_LH_BFX9 U1947 ( .A(n2457), .Z(n2454) );
  HS65_LH_BFX9 U1948 ( .A(n2457), .Z(n2455) );
  HS65_LH_BFX9 U1949 ( .A(n2453), .Z(n2450) );
  HS65_LH_BFX9 U1950 ( .A(n2466), .Z(n2463) );
  HS65_LH_IVX9 U1951 ( .A(n2636), .Z(n2635) );
  HS65_LH_IVX9 U1952 ( .A(n2633), .Z(n2632) );
  HS65_LH_IVX9 U1953 ( .A(n2449), .Z(n2448) );
  HS65_LH_BFX9 U1954 ( .A(n2668), .Z(n2421) );
  HS65_LH_BFX9 U1955 ( .A(n2458), .Z(n2459) );
  HS65_LH_BFX9 U1956 ( .A(n2484), .Z(n2485) );
  HS65_LH_BFX9 U1957 ( .A(n2497), .Z(n2498) );
  HS65_LH_BFX9 U1958 ( .A(n2510), .Z(n2511) );
  HS65_LH_BFX9 U1959 ( .A(n2471), .Z(n2472) );
  HS65_LH_BFX9 U1960 ( .A(n2453), .Z(n2451) );
  HS65_LH_BFX9 U1961 ( .A(n2479), .Z(n2477) );
  HS65_LH_BFX9 U1962 ( .A(n2470), .Z(n2467) );
  HS65_LH_BFX9 U1963 ( .A(n2496), .Z(n2493) );
  HS65_LH_BFX9 U1964 ( .A(n2509), .Z(n2506) );
  HS65_LH_BFX9 U1965 ( .A(n2522), .Z(n2519) );
  HS65_LH_BFX9 U1966 ( .A(n2470), .Z(n2468) );
  HS65_LH_BFX9 U1967 ( .A(n2496), .Z(n2494) );
  HS65_LH_BFX9 U1968 ( .A(n2509), .Z(n2507) );
  HS65_LH_BFX9 U1969 ( .A(n2522), .Z(n2520) );
  HS65_LH_BFX9 U1970 ( .A(n2483), .Z(n2480) );
  HS65_LH_BFX9 U1971 ( .A(n2479), .Z(n2476) );
  HS65_LH_BFX9 U1972 ( .A(n2492), .Z(n2489) );
  HS65_LH_BFX9 U1973 ( .A(n2505), .Z(n2502) );
  HS65_LH_BFX9 U1974 ( .A(n2518), .Z(n2515) );
  HS65_LH_BFX9 U1975 ( .A(n2483), .Z(n2481) );
  HS65_LH_IVX9 U1976 ( .A(n2642), .Z(n2641) );
  HS65_LH_IVX9 U1977 ( .A(n2639), .Z(n2638) );
  HS65_LH_IVX9 U1978 ( .A(n2648), .Z(n2647) );
  HS65_LH_IVX9 U1979 ( .A(n2645), .Z(n2644) );
  HS65_LH_IVX9 U1980 ( .A(n2462), .Z(n2461) );
  HS65_LH_IVX9 U1981 ( .A(n2475), .Z(n2474) );
  HS65_LH_IVX9 U1982 ( .A(n2488), .Z(n2487) );
  HS65_LH_IVX9 U1983 ( .A(n2501), .Z(n2500) );
  HS65_LH_IVX9 U1984 ( .A(n2514), .Z(n2513) );
  HS65_LH_BFX9 U1985 ( .A(n2536), .Z(n2537) );
  HS65_LH_BFX9 U1986 ( .A(n2549), .Z(n2550) );
  HS65_LH_BFX9 U1987 ( .A(n2523), .Z(n2524) );
  HS65_LH_BFX9 U1988 ( .A(n2535), .Z(n2533) );
  HS65_LH_BFX9 U1989 ( .A(n2466), .Z(n2464) );
  HS65_LH_BFX9 U1990 ( .A(n2492), .Z(n2490) );
  HS65_LH_BFX9 U1991 ( .A(n2505), .Z(n2503) );
  HS65_LH_BFX9 U1992 ( .A(n2518), .Z(n2516) );
  HS65_LH_BFX9 U1993 ( .A(n2561), .Z(n2558) );
  HS65_LH_BFX9 U1994 ( .A(n2548), .Z(n2545) );
  HS65_LH_BFX9 U1995 ( .A(n2548), .Z(n2546) );
  HS65_LH_BFX9 U1996 ( .A(n2561), .Z(n2559) );
  HS65_LH_BFX9 U1997 ( .A(n2535), .Z(n2532) );
  HS65_LH_BFX9 U1998 ( .A(n2531), .Z(n2528) );
  HS65_LH_BFX9 U1999 ( .A(n2544), .Z(n2541) );
  HS65_LH_BFX9 U2000 ( .A(n2557), .Z(n2554) );
  HS65_LH_IVX9 U2001 ( .A(n2654), .Z(n2653) );
  HS65_LH_IVX9 U2002 ( .A(n2657), .Z(n2656) );
  HS65_LH_IVX9 U2003 ( .A(n2651), .Z(n2650) );
  HS65_LH_IVX9 U2004 ( .A(n2527), .Z(n2526) );
  HS65_LH_IVX9 U2005 ( .A(n2540), .Z(n2539) );
  HS65_LH_IVX9 U2006 ( .A(n2553), .Z(n2552) );
  HS65_LH_IVX9 U2007 ( .A(n510), .Z(n2662) );
  HS65_LH_IVX9 U2008 ( .A(n462), .Z(n2661) );
  HS65_LH_BFX9 U2009 ( .A(n2666), .Z(n2418) );
  HS65_LH_BFX9 U2010 ( .A(n2668), .Z(n2420) );
  HS65_LH_BFX9 U2011 ( .A(n2666), .Z(n2419) );
  HS65_LH_BFX9 U2012 ( .A(n2433), .Z(n2430) );
  HS65_LH_BFX9 U2013 ( .A(n2471), .Z(n2473) );
  HS65_LH_BFX9 U2014 ( .A(n2531), .Z(n2529) );
  HS65_LH_BFX9 U2015 ( .A(n2544), .Z(n2542) );
  HS65_LH_BFX9 U2016 ( .A(n2557), .Z(n2555) );
  HS65_LH_BFX9 U2017 ( .A(n2445), .Z(n2447) );
  HS65_LH_BFX9 U2018 ( .A(n2458), .Z(n2460) );
  HS65_LH_BFX9 U2019 ( .A(n2484), .Z(n2486) );
  HS65_LH_BFX9 U2020 ( .A(n2433), .Z(n2432) );
  HS65_LH_IVX9 U2021 ( .A(n419), .Z(n2665) );
  HS65_LH_IVX9 U2022 ( .A(n352), .Z(n2664) );
  HS65_LH_IVX9 U2023 ( .A(n383), .Z(n2660) );
  HS65_LH_IVX9 U2024 ( .A(n328), .Z(n2659) );
  HS65_LH_BFX9 U2025 ( .A(n2523), .Z(n2525) );
  HS65_LH_BFX9 U2026 ( .A(n2497), .Z(n2499) );
  HS65_LH_BFX9 U2027 ( .A(n2510), .Z(n2512) );
  HS65_LH_BFX9 U2028 ( .A(n2457), .Z(n2456) );
  HS65_LH_BFX9 U2029 ( .A(n2470), .Z(n2469) );
  HS65_LH_BFX9 U2030 ( .A(n2453), .Z(n2452) );
  HS65_LH_BFX9 U2031 ( .A(n2466), .Z(n2465) );
  HS65_LH_BFX9 U2032 ( .A(n2479), .Z(n2478) );
  HS65_LH_IVX9 U2033 ( .A(n309), .Z(n2663) );
  HS65_LH_IVX9 U2034 ( .A(n297), .Z(n2658) );
  HS65_LH_BFX9 U2035 ( .A(n2433), .Z(n2431) );
  HS65_LH_BFX9 U2036 ( .A(n2536), .Z(n2538) );
  HS65_LH_BFX9 U2037 ( .A(n2549), .Z(n2551) );
  HS65_LH_BFX9 U2038 ( .A(n2496), .Z(n2495) );
  HS65_LH_BFX9 U2039 ( .A(n2509), .Z(n2508) );
  HS65_LH_BFX9 U2040 ( .A(n2483), .Z(n2482) );
  HS65_LH_BFX9 U2041 ( .A(n2492), .Z(n2491) );
  HS65_LH_BFX9 U2042 ( .A(n2505), .Z(n2504) );
  HS65_LH_BFX9 U2043 ( .A(n2666), .Z(n2417) );
  HS65_LH_BFX9 U2044 ( .A(n2522), .Z(n2521) );
  HS65_LH_BFX9 U2045 ( .A(n2531), .Z(n2530) );
  HS65_LH_BFX9 U2046 ( .A(n2518), .Z(n2517) );
  HS65_LH_BFX9 U2047 ( .A(n2548), .Z(n2547) );
  HS65_LH_BFX9 U2048 ( .A(n2561), .Z(n2560) );
  HS65_LH_BFX9 U2049 ( .A(n2535), .Z(n2534) );
  HS65_LH_BFX9 U2050 ( .A(n2544), .Z(n2543) );
  HS65_LH_BFX9 U2051 ( .A(n2557), .Z(n2556) );
  HS65_LH_IVX9 U2052 ( .A(n2713), .Z(n2668) );
  HS65_LH_BFX9 U2053 ( .A(n2723), .Z(n2457) );
  HS65_LH_BFX9 U2054 ( .A(n2721), .Z(n2453) );
  HS65_LH_BFX9 U2055 ( .A(n2764), .Z(n2466) );
  HS65_LH_IVX9 U2056 ( .A(n19), .Z(n2633) );
  HS65_LH_IVX9 U2057 ( .A(n2719), .Z(n2449) );
  HS65_LH_IVX9 U2058 ( .A(n2762), .Z(n2462) );
  HS65_LH_HA1X4 U2059 ( .A0(n2566), .B0(n2563), .CO(n1005), .S0(n1038) );
  HS65_LH_BFX9 U2060 ( .A(n2718), .Z(n2445) );
  HS65_LH_BFX9 U2061 ( .A(b[2]), .Z(n2568) );
  HS65_LH_BFX9 U2062 ( .A(n2562), .Z(n2563) );
  HS65_LH_BFX9 U2063 ( .A(n2436), .Z(n2434) );
  HS65_LH_BFX9 U2064 ( .A(n2444), .Z(n2441) );
  HS65_LH_BFX9 U2065 ( .A(n2444), .Z(n2442) );
  HS65_LH_IVX9 U2066 ( .A(n2633), .Z(n2631) );
  HS65_LH_BFX9 U2067 ( .A(n2444), .Z(n2443) );
  HS65_LH_BFX9 U2068 ( .A(n2766), .Z(n2470) );
  HS65_LH_BFX9 U2069 ( .A(n2809), .Z(n2483) );
  HS65_LH_IVX9 U2070 ( .A(n2891), .Z(n2501) );
  HS65_LH_IVX9 U2071 ( .A(n2934), .Z(n2514) );
  HS65_LH_BFX9 U2072 ( .A(n2852), .Z(n2496) );
  HS65_LH_BFX9 U2073 ( .A(n2895), .Z(n2509) );
  HS65_LH_BFX9 U2074 ( .A(n2938), .Z(n2522) );
  HS65_LH_BFX9 U2075 ( .A(n2850), .Z(n2492) );
  HS65_LH_BFX9 U2076 ( .A(n2893), .Z(n2505) );
  HS65_LH_BFX9 U2077 ( .A(n2936), .Z(n2518) );
  HS65_LH_BFX9 U2078 ( .A(n2807), .Z(n2479) );
  HS65_LH_IVX9 U2079 ( .A(n55), .Z(n2642) );
  HS65_LH_IVX9 U2080 ( .A(n43), .Z(n2639) );
  HS65_LH_IVX9 U2081 ( .A(n79), .Z(n2648) );
  HS65_LH_IVX9 U2082 ( .A(n67), .Z(n2645) );
  HS65_LH_IVX9 U2083 ( .A(n2848), .Z(n2488) );
  HS65_LH_IVX9 U2084 ( .A(n2977), .Z(n2527) );
  HS65_LH_IVX9 U2085 ( .A(n2805), .Z(n2475) );
  HS65_LH_BFX9 U2086 ( .A(n2761), .Z(n2458) );
  HS65_LH_BFX9 U2087 ( .A(n2804), .Z(n2471) );
  HS65_LH_BFX9 U2088 ( .A(n2847), .Z(n2484) );
  HS65_LH_BFX9 U2089 ( .A(n2890), .Z(n2497) );
  HS65_LH_BFX9 U2090 ( .A(n2933), .Z(n2510) );
  HS65_LH_BFX9 U2091 ( .A(b[3]), .Z(n2570) );
  HS65_LH_BFX9 U2092 ( .A(b[4]), .Z(n2572) );
  HS65_LH_BFX9 U2093 ( .A(n2562), .Z(n2564) );
  HS65_LH_BFX9 U2094 ( .A(b[2]), .Z(n2569) );
  HS65_LH_BFX9 U2095 ( .A(b[3]), .Z(n2571) );
  HS65_LH_BFX9 U2096 ( .A(n2440), .Z(n2437) );
  HS65_LH_BFX9 U2097 ( .A(b[4]), .Z(n2573) );
  HS65_LH_IVX9 U2098 ( .A(n2636), .Z(n2634) );
  HS65_LH_IVX9 U2099 ( .A(n31), .Z(n2636) );
  HS65_LH_IVX9 U2100 ( .A(n2642), .Z(n2640) );
  HS65_LH_IVX9 U2101 ( .A(n2639), .Z(n2637) );
  HS65_LH_IVX9 U2102 ( .A(n2648), .Z(n2646) );
  HS65_LH_IVX9 U2103 ( .A(n2645), .Z(n2643) );
  HS65_LH_BFX9 U2104 ( .A(n2562), .Z(n2565) );
  HS65_LH_BFX9 U2105 ( .A(n2440), .Z(n2439) );
  HS65_LH_BFX9 U2106 ( .A(n3067), .Z(n2561) );
  HS65_LH_BFX9 U2107 ( .A(n3022), .Z(n2544) );
  HS65_LH_BFX9 U2108 ( .A(n2981), .Z(n2535) );
  HS65_LH_BFX9 U2109 ( .A(n3024), .Z(n2548) );
  HS65_LH_BFX9 U2110 ( .A(n2979), .Z(n2531) );
  HS65_LH_BFX9 U2111 ( .A(n3065), .Z(n2557) );
  HS65_LH_IVX9 U2112 ( .A(n115), .Z(n2657) );
  HS65_LH_IVX9 U2113 ( .A(n3020), .Z(n2540) );
  HS65_LH_IVX9 U2114 ( .A(n3063), .Z(n2553) );
  HS65_LH_BFX9 U2115 ( .A(n2976), .Z(n2523) );
  HS65_LH_BFX9 U2116 ( .A(n3019), .Z(n2536) );
  HS65_LH_BFX9 U2117 ( .A(n3062), .Z(n2549) );
  HS65_LH_IVX9 U2118 ( .A(n2654), .Z(n2652) );
  HS65_LH_IVX9 U2119 ( .A(n103), .Z(n2654) );
  HS65_LH_IVX9 U2120 ( .A(n2651), .Z(n2649) );
  HS65_LH_IVX9 U2121 ( .A(n91), .Z(n2651) );
  HS65_LH_BFX9 U2122 ( .A(b[11]), .Z(n2586) );
  HS65_LH_BFX9 U2123 ( .A(b[11]), .Z(n2587) );
  HS65_LH_BFX9 U2124 ( .A(n2440), .Z(n2438) );
  HS65_LH_BFX9 U2125 ( .A(n2436), .Z(n2435) );
  HS65_LH_IVX9 U2126 ( .A(n2657), .Z(n2655) );
  HS65_LH_BFX9 U2127 ( .A(n2429), .Z(n2428) );
  HS65_LH_BFX9 U2128 ( .A(n2672), .Z(n2433) );
  HS65_LH_IVX9 U2129 ( .A(n2673), .Z(n2666) );
  HS65_LH_BFX9 U2130 ( .A(b[20]), .Z(n2604) );
  HS65_LH_BFX9 U2131 ( .A(n2425), .Z(n2423) );
  HS65_LH_BFX9 U2132 ( .A(n2429), .Z(n2426) );
  HS65_LH_BFX9 U2133 ( .A(b[27]), .Z(n2618) );
  HS65_LH_BFX9 U2134 ( .A(b[28]), .Z(n2620) );
  HS65_LH_BFX9 U2135 ( .A(n2425), .Z(n2424) );
  HS65_LH_BFX9 U2136 ( .A(b[20]), .Z(n2605) );
  HS65_LH_BFX9 U2137 ( .A(b[31]), .Z(n2626) );
  HS65_LH_BFX9 U2138 ( .A(b[27]), .Z(n2619) );
  HS65_LH_BFX9 U2139 ( .A(b[28]), .Z(n2621) );
  HS65_LH_BFX9 U2140 ( .A(b[31]), .Z(n2627) );
  HS65_LH_BFX9 U2141 ( .A(n2429), .Z(n2427) );
  HS65_LH_BFX9 U2142 ( .A(n2681), .Z(n2444) );
  HS65_LH_BFX9 U2143 ( .A(n2677), .Z(n2436) );
  HS65_LH_BFX9 U2144 ( .A(b[0]), .Z(n2562) );
  HS65_LH_BFX9 U2145 ( .A(n2679), .Z(n2440) );
  HS65_LH_BFX9 U2146 ( .A(b[1]), .Z(n2566) );
  HS65_LH_BFX9 U2147 ( .A(b[5]), .Z(n2574) );
  HS65_LH_BFX9 U2148 ( .A(b[7]), .Z(n2578) );
  HS65_LH_BFX9 U2149 ( .A(b[6]), .Z(n2576) );
  HS65_LH_BFX9 U2150 ( .A(b[8]), .Z(n2580) );
  HS65_LH_BFX9 U2151 ( .A(b[5]), .Z(n2575) );
  HS65_LH_BFX9 U2152 ( .A(b[1]), .Z(n2567) );
  HS65_LH_BFX9 U2153 ( .A(b[6]), .Z(n2577) );
  HS65_LH_BFX9 U2154 ( .A(n2671), .Z(n2429) );
  HS65_LH_BFX9 U2155 ( .A(b[12]), .Z(n2588) );
  HS65_LH_BFX9 U2156 ( .A(b[13]), .Z(n2590) );
  HS65_LH_BFX9 U2157 ( .A(b[9]), .Z(n2582) );
  HS65_LH_BFX9 U2158 ( .A(b[14]), .Z(n2592) );
  HS65_LH_BFX9 U2159 ( .A(b[10]), .Z(n2584) );
  HS65_LH_BFX9 U2160 ( .A(b[12]), .Z(n2589) );
  HS65_LH_BFX9 U2161 ( .A(b[7]), .Z(n2579) );
  HS65_LH_BFX9 U2162 ( .A(b[9]), .Z(n2583) );
  HS65_LH_BFX9 U2163 ( .A(b[8]), .Z(n2581) );
  HS65_LH_BFX9 U2164 ( .A(b[10]), .Z(n2585) );
  HS65_LH_BFX9 U2165 ( .A(n2670), .Z(n2425) );
  HS65_LH_BFX9 U2166 ( .A(b[19]), .Z(n2602) );
  HS65_LH_BFX9 U2167 ( .A(b[18]), .Z(n2600) );
  HS65_LH_BFX9 U2168 ( .A(b[15]), .Z(n2594) );
  HS65_LH_BFX9 U2169 ( .A(b[17]), .Z(n2598) );
  HS65_LH_BFX9 U2170 ( .A(b[21]), .Z(n2606) );
  HS65_LH_BFX9 U2171 ( .A(b[16]), .Z(n2596) );
  HS65_LH_BFX9 U2172 ( .A(b[19]), .Z(n2603) );
  HS65_LH_BFX9 U2173 ( .A(b[13]), .Z(n2591) );
  HS65_LH_BFX9 U2174 ( .A(b[18]), .Z(n2601) );
  HS65_LH_BFX9 U2175 ( .A(b[15]), .Z(n2595) );
  HS65_LH_BFX9 U2176 ( .A(b[17]), .Z(n2599) );
  HS65_LH_BFX9 U2177 ( .A(b[14]), .Z(n2593) );
  HS65_LH_BFX9 U2178 ( .A(b[16]), .Z(n2597) );
  HS65_LH_BFX9 U2179 ( .A(b[23]), .Z(n2610) );
  HS65_LH_BFX9 U2180 ( .A(b[25]), .Z(n2614) );
  HS65_LH_BFX9 U2181 ( .A(b[24]), .Z(n2612) );
  HS65_LH_BFX9 U2182 ( .A(b[26]), .Z(n2616) );
  HS65_LH_BFX9 U2183 ( .A(b[22]), .Z(n2608) );
  HS65_LH_BFX9 U2184 ( .A(b[23]), .Z(n2611) );
  HS65_LH_BFX9 U2185 ( .A(b[25]), .Z(n2615) );
  HS65_LH_BFX9 U2186 ( .A(b[24]), .Z(n2613) );
  HS65_LH_BFX9 U2187 ( .A(b[21]), .Z(n2607) );
  HS65_LH_BFX9 U2188 ( .A(b[22]), .Z(n2609) );
  HS65_LH_BFX9 U2189 ( .A(b[29]), .Z(n2622) );
  HS65_LH_BFX9 U2190 ( .A(b[30]), .Z(n2624) );
  HS65_LH_BFX9 U2191 ( .A(b[26]), .Z(n2617) );
  HS65_LH_BFX9 U2192 ( .A(b[29]), .Z(n2623) );
  HS65_LH_BFX9 U2193 ( .A(b[30]), .Z(n2625) );
  HS65_LHS_XOR3X2 U2194 ( .A(n292), .B(n227), .C(n2669), .Z(product[63]) );
  HS65_LH_AO22X4 U2195 ( .A(n2627), .B(n2423), .C(n2419), .D(n1006), .Z(n2669)
         );
  HS65_LH_MX41X4 U2196 ( .D0(n1025), .S0(n2419), .D1(n2593), .S1(n2427), .D2(
        n2591), .S2(n2431), .D3(n2589), .S3(n2423), .Z(n419) );
  HS65_LH_MX41X4 U2197 ( .D0(n1019), .S0(n2419), .D1(n2601), .S1(n2423), .D2(
        n2603), .S2(n2430), .D3(n2605), .S3(n2426), .Z(n352) );
  HS65_LH_MX41X4 U2198 ( .D0(n1013), .S0(n2419), .D1(n2613), .S1(n2423), .D2(
        n2615), .S2(n2430), .D3(n2617), .S3(n2426), .Z(n309) );
  HS65_LH_OA12X4 U2199 ( .A(n2673), .B(n2667), .C(n2674), .Z(n292) );
  HS65_LH_OAI22X1 U2200 ( .A(n2625), .B(n2675), .C(n2423), .D(n2675), .Z(n2674) );
  HS65_LH_AND2X4 U2201 ( .A(n2626), .B(n2430), .Z(n2675) );
  HS65_LHS_XOR2X3 U2202 ( .A(n2628), .B(n2676), .Z(n1419) );
  HS65_LH_AO22X4 U2203 ( .A(n2565), .B(n2434), .C(n2422), .D(n2564), .Z(n2676)
         );
  HS65_LHS_XOR2X3 U2204 ( .A(n2628), .B(n2678), .Z(n1418) );
  HS65_LH_AO222X4 U2205 ( .A(n2564), .B(n2437), .C(n2434), .D(n2566), .E(n2422), .F(n1038), .Z(n2678) );
  HS65_LHS_XOR2X3 U2206 ( .A(n2628), .B(n2680), .Z(n1417) );
  HS65_LH_MX41X4 U2207 ( .D0(n1037), .S0(n2422), .D1(n2442), .S1(n2564), .D2(
        n2439), .S2(n2566), .D3(n2569), .S3(n2434), .Z(n2680) );
  HS65_LHS_XOR2X3 U2208 ( .A(n2628), .B(n2682), .Z(n1416) );
  HS65_LH_MX41X4 U2209 ( .D0(n1036), .S0(n2421), .D1(n2443), .S1(n2567), .D2(
        n2569), .S2(n2437), .D3(n2571), .S3(n2434), .Z(n2682) );
  HS65_LHS_XOR2X3 U2210 ( .A(n2629), .B(n2683), .Z(n1415) );
  HS65_LH_MX41X4 U2211 ( .D0(n1035), .S0(n2422), .D1(n2443), .S1(n2569), .D2(
        n2571), .S2(n2437), .D3(n2573), .S3(n2434), .Z(n2683) );
  HS65_LHS_XOR2X3 U2212 ( .A(n2628), .B(n2684), .Z(n1414) );
  HS65_LH_MX41X4 U2213 ( .D0(n1034), .S0(n2422), .D1(n2571), .S1(n2441), .D2(
        n2573), .S2(n2437), .D3(n2575), .S3(n2434), .Z(n2684) );
  HS65_LHS_XOR2X3 U2214 ( .A(n2628), .B(n2685), .Z(n1413) );
  HS65_LH_MX41X4 U2215 ( .D0(n1033), .S0(n2421), .D1(n2573), .S1(n2441), .D2(
        n2575), .S2(n2437), .D3(n2577), .S3(n2434), .Z(n2685) );
  HS65_LHS_XOR2X3 U2216 ( .A(n2628), .B(n2686), .Z(n1412) );
  HS65_LH_MX41X4 U2217 ( .D0(n1032), .S0(n2421), .D1(n2575), .S1(n2441), .D2(
        n2577), .S2(n2437), .D3(n2579), .S3(n2434), .Z(n2686) );
  HS65_LHS_XOR2X3 U2218 ( .A(n2628), .B(n2687), .Z(n1411) );
  HS65_LH_MX41X4 U2219 ( .D0(n1031), .S0(n2421), .D1(n2577), .S1(n2441), .D2(
        n2579), .S2(n2437), .D3(n2581), .S3(n2434), .Z(n2687) );
  HS65_LHS_XOR2X3 U2220 ( .A(n2628), .B(n2688), .Z(n1410) );
  HS65_LH_MX41X4 U2221 ( .D0(n1030), .S0(n2421), .D1(n2579), .S1(n2441), .D2(
        n2581), .S2(n2437), .D3(n2583), .S3(n2434), .Z(n2688) );
  HS65_LHS_XOR2X3 U2222 ( .A(n2628), .B(n2689), .Z(n1409) );
  HS65_LH_MX41X4 U2223 ( .D0(n1029), .S0(n2421), .D1(n2581), .S1(n2441), .D2(
        n2583), .S2(n2437), .D3(n2585), .S3(n2434), .Z(n2689) );
  HS65_LHS_XOR2X3 U2224 ( .A(n2628), .B(n2690), .Z(n1408) );
  HS65_LH_MX41X4 U2225 ( .D0(n1028), .S0(n2421), .D1(n2583), .S1(n2441), .D2(
        n2585), .S2(n2437), .D3(n2587), .S3(n2434), .Z(n2690) );
  HS65_LHS_XOR2X3 U2226 ( .A(n2628), .B(n2691), .Z(n1407) );
  HS65_LH_MX41X4 U2227 ( .D0(n1027), .S0(n2421), .D1(n2585), .S1(n2441), .D2(
        n2587), .S2(n2437), .D3(n2435), .S3(n2589), .Z(n2691) );
  HS65_LHS_XOR2X3 U2228 ( .A(n2628), .B(n2692), .Z(n1406) );
  HS65_LH_MX41X4 U2229 ( .D0(n1026), .S0(n2421), .D1(n2587), .S1(n2441), .D2(
        n2438), .S2(n2588), .D3(n2435), .S3(n2591), .Z(n2692) );
  HS65_LHS_XOR2X3 U2230 ( .A(n2628), .B(n2693), .Z(n1405) );
  HS65_LH_MX41X4 U2231 ( .D0(n2422), .S0(n1025), .D1(n2442), .S1(n2589), .D2(
        n2438), .S2(n2590), .D3(n2435), .S3(n2593), .Z(n2693) );
  HS65_LHS_XOR2X3 U2232 ( .A(n2628), .B(n2694), .Z(n1404) );
  HS65_LH_MX41X4 U2233 ( .D0(n1024), .S0(n2421), .D1(n2442), .S1(n2591), .D2(
        n2438), .S2(n2592), .D3(n2595), .S3(n2434), .Z(n2694) );
  HS65_LHS_XOR2X3 U2234 ( .A(n2629), .B(n2695), .Z(n1403) );
  HS65_LH_MX41X4 U2235 ( .D0(n1023), .S0(n2421), .D1(n2442), .S1(n2593), .D2(
        n2595), .S2(n2437), .D3(n2597), .S3(n2434), .Z(n2695) );
  HS65_LHS_XOR2X3 U2236 ( .A(n2629), .B(n2696), .Z(n1402) );
  HS65_LH_MX41X4 U2237 ( .D0(n1022), .S0(n2420), .D1(n2595), .S1(n2441), .D2(
        n2597), .S2(n2437), .D3(n2599), .S3(n2434), .Z(n2696) );
  HS65_LHS_XOR2X3 U2238 ( .A(n2629), .B(n2697), .Z(n1401) );
  HS65_LH_MX41X4 U2239 ( .D0(n1021), .S0(n2420), .D1(n2597), .S1(n2441), .D2(
        n2599), .S2(n2437), .D3(n2435), .S3(n2601), .Z(n2697) );
  HS65_LHS_XOR2X3 U2240 ( .A(n2629), .B(n2698), .Z(n1400) );
  HS65_LH_MX41X4 U2241 ( .D0(n1020), .S0(n2420), .D1(n2599), .S1(n2441), .D2(
        n2438), .S2(n2600), .D3(n2435), .S3(n2603), .Z(n2698) );
  HS65_LHS_XOR2X3 U2242 ( .A(n2629), .B(n2699), .Z(n1399) );
  HS65_LH_MX41X4 U2243 ( .D0(n2422), .S0(n1019), .D1(n2442), .S1(n2601), .D2(
        n2438), .S2(n2602), .D3(n2435), .S3(n2605), .Z(n2699) );
  HS65_LHS_XOR2X3 U2244 ( .A(n2629), .B(n2700), .Z(n1398) );
  HS65_LH_MX41X4 U2245 ( .D0(n1018), .S0(n2420), .D1(n2442), .S1(n2603), .D2(
        n2438), .S2(n2604), .D3(n2607), .S3(n2435), .Z(n2700) );
  HS65_LHS_XOR2X3 U2246 ( .A(n2629), .B(n2701), .Z(n1397) );
  HS65_LH_MX41X4 U2247 ( .D0(n1017), .S0(n2420), .D1(n2442), .S1(n2605), .D2(
        n2607), .S2(n2438), .D3(n2609), .S3(n2434), .Z(n2701) );
  HS65_LHS_XOR2X3 U2248 ( .A(n2629), .B(n2702), .Z(n1396) );
  HS65_LH_MX41X4 U2249 ( .D0(n1016), .S0(n2420), .D1(n2607), .S1(n2442), .D2(
        n2609), .S2(n2438), .D3(n2611), .S3(n2435), .Z(n2702) );
  HS65_LHS_XOR2X3 U2250 ( .A(n2629), .B(n2703), .Z(n1395) );
  HS65_LH_MX41X4 U2251 ( .D0(n1015), .S0(n2421), .D1(n2609), .S1(n2442), .D2(
        n2611), .S2(n2438), .D3(n2435), .S3(n2613), .Z(n2703) );
  HS65_LHS_XOR2X3 U2252 ( .A(n2629), .B(n2704), .Z(n1394) );
  HS65_LH_MX41X4 U2253 ( .D0(n1014), .S0(n2420), .D1(n2611), .S1(n2442), .D2(
        n2439), .S2(n2612), .D3(n2435), .S3(n2615), .Z(n2704) );
  HS65_LHS_XOR2X3 U2254 ( .A(n2629), .B(n2705), .Z(n1393) );
  HS65_LH_MX41X4 U2255 ( .D0(n2422), .S0(n1013), .D1(n2443), .S1(n2613), .D2(
        n2438), .S2(n2614), .D3(n2435), .S3(n2617), .Z(n2705) );
  HS65_LHS_XOR2X3 U2256 ( .A(n2629), .B(n2706), .Z(n1392) );
  HS65_LH_MX41X4 U2257 ( .D0(n1012), .S0(n2420), .D1(n2443), .S1(n2615), .D2(
        n2439), .S2(n2616), .D3(n2619), .S3(n2435), .Z(n2706) );
  HS65_LHS_XOR2X3 U2258 ( .A(n2629), .B(n2707), .Z(n1391) );
  HS65_LH_MX41X4 U2259 ( .D0(n1011), .S0(n2420), .D1(n2443), .S1(n2617), .D2(
        n2619), .S2(n2438), .D3(n2621), .S3(n2435), .Z(n2707) );
  HS65_LHS_XOR2X3 U2260 ( .A(n2629), .B(n2708), .Z(n1390) );
  HS65_LH_MX41X4 U2261 ( .D0(n1010), .S0(n2420), .D1(n2619), .S1(n2442), .D2(
        n2621), .S2(n2438), .D3(n2623), .S3(n2435), .Z(n2708) );
  HS65_LHS_XOR2X3 U2262 ( .A(n2629), .B(n2709), .Z(n1389) );
  HS65_LH_MX41X4 U2263 ( .D0(n1009), .S0(n2420), .D1(n2621), .S1(n2442), .D2(
        n2623), .S2(n2438), .D3(n2625), .S3(n2435), .Z(n2709) );
  HS65_LHS_XOR2X3 U2264 ( .A(n2629), .B(n2710), .Z(n1388) );
  HS65_LH_MX41X4 U2265 ( .D0(n1008), .S0(n2420), .D1(n2623), .S1(n2442), .D2(
        n2625), .S2(n2438), .D3(n2435), .S3(n2627), .Z(n2710) );
  HS65_LH_NOR2AX3 U2266 ( .A(a[0]), .B(n2711), .Z(n2677) );
  HS65_LHS_XOR2X3 U2267 ( .A(n2629), .B(n2712), .Z(n1387) );
  HS65_LH_OAI12X2 U2268 ( .A(n2667), .B(n2713), .C(n2714), .Z(n2712) );
  HS65_LH_OAI22X1 U2269 ( .A(n2625), .B(n2715), .C(n2441), .D(n2715), .Z(n2714) );
  HS65_LH_AND2X4 U2270 ( .A(n2438), .B(n2626), .Z(n2715) );
  HS65_LH_NOR2AX3 U2271 ( .A(a[1]), .B(a[0]), .Z(n2679) );
  HS65_LHS_XOR2X3 U2272 ( .A(n2630), .B(n2716), .Z(n1386) );
  HS65_LH_AOI22X1 U2273 ( .A(n2422), .B(n1006), .C(n2443), .D(n2627), .Z(n2716) );
  HS65_LH_NOR3AX2 U2274 ( .A(n2711), .B(a[0]), .C(a[1]), .Z(n2681) );
  HS65_LH_NAND2X2 U2275 ( .A(a[0]), .B(n2711), .Z(n2713) );
  HS65_LHS_XOR2X3 U2276 ( .A(n2629), .B(a[1]), .Z(n2711) );
  HS65_LHS_XOR2X3 U2277 ( .A(n2631), .B(n2717), .Z(n1384) );
  HS65_LH_AO22X4 U2278 ( .A(n2565), .B(n2446), .C(n2564), .D(n2719), .Z(n2717)
         );
  HS65_LHS_XOR2X3 U2279 ( .A(n2631), .B(n2720), .Z(n1383) );
  HS65_LH_AO222X4 U2280 ( .A(n2567), .B(n2446), .C(n2563), .D(n2450), .E(n1038), .F(n2448), .Z(n2720) );
  HS65_LHS_XOR2X3 U2281 ( .A(n2631), .B(n2722), .Z(n1382) );
  HS65_LH_MX41X4 U2282 ( .D0(n2448), .S0(n1037), .D1(n2455), .S1(n2564), .D2(
        n2450), .S2(n2566), .D3(n2446), .S3(n2569), .Z(n2722) );
  HS65_LHS_XOR2X3 U2283 ( .A(n2631), .B(n2724), .Z(n1381) );
  HS65_LH_MX41X4 U2284 ( .D0(n2448), .S0(n1036), .D1(n2454), .S1(n2567), .D2(
        n2450), .S2(n2568), .D3(n2446), .S3(n2571), .Z(n2724) );
  HS65_LHS_XOR2X3 U2285 ( .A(n2631), .B(n2725), .Z(n1380) );
  HS65_LH_MX41X4 U2286 ( .D0(n2448), .S0(n1035), .D1(n2454), .S1(n2569), .D2(
        n2450), .S2(n2570), .D3(n2446), .S3(n2573), .Z(n2725) );
  HS65_LHS_XOR2X3 U2287 ( .A(n2631), .B(n2726), .Z(n1379) );
  HS65_LH_MX41X4 U2288 ( .D0(n2448), .S0(n1034), .D1(n2454), .S1(n2571), .D2(
        n2450), .S2(n2572), .D3(n2446), .S3(n2575), .Z(n2726) );
  HS65_LHS_XOR2X3 U2289 ( .A(n2631), .B(n2727), .Z(n1378) );
  HS65_LH_MX41X4 U2290 ( .D0(n2448), .S0(n1033), .D1(n2454), .S1(n2573), .D2(
        n2450), .S2(n2574), .D3(n2446), .S3(n2577), .Z(n2727) );
  HS65_LHS_XOR2X3 U2291 ( .A(n2631), .B(n2728), .Z(n1377) );
  HS65_LH_MX41X4 U2292 ( .D0(n2448), .S0(n1032), .D1(n2454), .S1(n2575), .D2(
        n2450), .S2(n2576), .D3(n2446), .S3(n2579), .Z(n2728) );
  HS65_LHS_XOR2X3 U2293 ( .A(n2631), .B(n2729), .Z(n1376) );
  HS65_LH_MX41X4 U2294 ( .D0(n2448), .S0(n1031), .D1(n2454), .S1(n2577), .D2(
        n2450), .S2(n2578), .D3(n2446), .S3(n2581), .Z(n2729) );
  HS65_LHS_XOR2X3 U2295 ( .A(n2631), .B(n2730), .Z(n1375) );
  HS65_LH_MX41X4 U2296 ( .D0(n2448), .S0(n1030), .D1(n2454), .S1(n2579), .D2(
        n2451), .S2(n2580), .D3(n2446), .S3(n2583), .Z(n2730) );
  HS65_LHS_XOR2X3 U2297 ( .A(n2631), .B(n2731), .Z(n1374) );
  HS65_LH_MX41X4 U2298 ( .D0(n2448), .S0(n1029), .D1(n2454), .S1(n2581), .D2(
        n2450), .S2(n2582), .D3(n2446), .S3(n2585), .Z(n2731) );
  HS65_LHS_XOR2X3 U2299 ( .A(n2631), .B(n2732), .Z(n1373) );
  HS65_LH_MX41X4 U2300 ( .D0(n2448), .S0(n1028), .D1(n2454), .S1(n2583), .D2(
        n2450), .S2(n2584), .D3(n2446), .S3(n2587), .Z(n2732) );
  HS65_LHS_XOR2X3 U2301 ( .A(n2631), .B(n2733), .Z(n1372) );
  HS65_LH_MX41X4 U2302 ( .D0(n2448), .S0(n1027), .D1(n2454), .S1(n2585), .D2(
        n2450), .S2(n2586), .D3(n2446), .S3(n2589), .Z(n2733) );
  HS65_LHS_XOR2X3 U2303 ( .A(n2631), .B(n2734), .Z(n1371) );
  HS65_LH_MX41X4 U2304 ( .D0(n2448), .S0(n1026), .D1(n2454), .S1(n2587), .D2(
        n2451), .S2(n2588), .D3(n2446), .S3(n2591), .Z(n2734) );
  HS65_LHS_XOR2X3 U2305 ( .A(n2631), .B(n2735), .Z(n1370) );
  HS65_LH_MX41X4 U2306 ( .D0(n2448), .S0(n1025), .D1(n2454), .S1(n2589), .D2(
        n2451), .S2(n2590), .D3(n2446), .S3(n2592), .Z(n2735) );
  HS65_LHS_XOR2X3 U2307 ( .A(n2631), .B(n2736), .Z(n1369) );
  HS65_LH_MX41X4 U2308 ( .D0(n2448), .S0(n1024), .D1(n2455), .S1(n2591), .D2(
        n2451), .S2(n2592), .D3(n2446), .S3(n2595), .Z(n2736) );
  HS65_LHS_XOR2X3 U2309 ( .A(n2631), .B(n2737), .Z(n1368) );
  HS65_LH_MX41X4 U2310 ( .D0(n2448), .S0(n1023), .D1(n2455), .S1(n2593), .D2(
        n2451), .S2(n2594), .D3(n2446), .S3(n2597), .Z(n2737) );
  HS65_LHS_XOR2X3 U2311 ( .A(n2631), .B(n2738), .Z(n1367) );
  HS65_LH_MX41X4 U2312 ( .D0(n2448), .S0(n1022), .D1(n2455), .S1(n2595), .D2(
        n2451), .S2(n2596), .D3(n2447), .S3(n2599), .Z(n2738) );
  HS65_LHS_XOR2X3 U2313 ( .A(n2631), .B(n2739), .Z(n1366) );
  HS65_LH_MX41X4 U2314 ( .D0(n2448), .S0(n1021), .D1(n2455), .S1(n2597), .D2(
        n2451), .S2(n2598), .D3(n2447), .S3(n2600), .Z(n2739) );
  HS65_LHS_XOR2X3 U2315 ( .A(n19), .B(n2740), .Z(n1365) );
  HS65_LH_MX41X4 U2316 ( .D0(n2448), .S0(n1020), .D1(n2455), .S1(n2599), .D2(
        n2451), .S2(n2600), .D3(n2447), .S3(n2602), .Z(n2740) );
  HS65_LHS_XOR2X3 U2317 ( .A(n19), .B(n2741), .Z(n1364) );
  HS65_LH_MX41X4 U2318 ( .D0(n2448), .S0(n1019), .D1(n2455), .S1(n2601), .D2(
        n2451), .S2(n2602), .D3(n2447), .S3(n2604), .Z(n2741) );
  HS65_LHS_XOR2X3 U2319 ( .A(n19), .B(n2742), .Z(n1363) );
  HS65_LH_MX41X4 U2320 ( .D0(n2719), .S0(n1018), .D1(n2455), .S1(n2603), .D2(
        n2451), .S2(n2604), .D3(n2447), .S3(n2607), .Z(n2742) );
  HS65_LHS_XOR2X3 U2321 ( .A(n19), .B(n2743), .Z(n1362) );
  HS65_LH_MX41X4 U2322 ( .D0(n2719), .S0(n1017), .D1(n2455), .S1(n2605), .D2(
        n2451), .S2(n2606), .D3(n2447), .S3(n2609), .Z(n2743) );
  HS65_LHS_XOR2X3 U2323 ( .A(n2632), .B(n2744), .Z(n1361) );
  HS65_LH_MX41X4 U2324 ( .D0(n2719), .S0(n1016), .D1(n2455), .S1(n2607), .D2(
        n2451), .S2(n2608), .D3(n2447), .S3(n2611), .Z(n2744) );
  HS65_LHS_XOR2X3 U2325 ( .A(n2632), .B(n2745), .Z(n1360) );
  HS65_LH_MX41X4 U2326 ( .D0(n2719), .S0(n1015), .D1(n2455), .S1(n2609), .D2(
        n2451), .S2(n2610), .D3(n2447), .S3(n2612), .Z(n2745) );
  HS65_LHS_XOR2X3 U2327 ( .A(n2632), .B(n2746), .Z(n1359) );
  HS65_LH_MX41X4 U2328 ( .D0(n2719), .S0(n1014), .D1(n2455), .S1(n2611), .D2(
        n2451), .S2(n2612), .D3(n2447), .S3(n2614), .Z(n2746) );
  HS65_LHS_XOR2X3 U2329 ( .A(n2632), .B(n2747), .Z(n1358) );
  HS65_LH_MX41X4 U2330 ( .D0(n2719), .S0(n1013), .D1(n2455), .S1(n2613), .D2(
        n2452), .S2(n2614), .D3(n2447), .S3(n2616), .Z(n2747) );
  HS65_LHS_XOR2X3 U2331 ( .A(n2632), .B(n2748), .Z(n1357) );
  HS65_LH_MX41X4 U2332 ( .D0(n2719), .S0(n1012), .D1(n2456), .S1(n2615), .D2(
        n2452), .S2(n2616), .D3(n2447), .S3(n2619), .Z(n2748) );
  HS65_LHS_XOR2X3 U2333 ( .A(n2632), .B(n2749), .Z(n1356) );
  HS65_LH_MX41X4 U2334 ( .D0(n2719), .S0(n1011), .D1(n2456), .S1(n2617), .D2(
        n2452), .S2(n2618), .D3(n2447), .S3(n2621), .Z(n2749) );
  HS65_LHS_XOR2X3 U2335 ( .A(n2632), .B(n2750), .Z(n1355) );
  HS65_LH_MX41X4 U2336 ( .D0(n2719), .S0(n1010), .D1(n2456), .S1(n2619), .D2(
        n2452), .S2(n2620), .D3(n2447), .S3(n2623), .Z(n2750) );
  HS65_LHS_XOR2X3 U2337 ( .A(n2632), .B(n2751), .Z(n1354) );
  HS65_LH_MX41X4 U2338 ( .D0(n2719), .S0(n1009), .D1(n2456), .S1(n2621), .D2(
        n2452), .S2(n2622), .D3(n2447), .S3(n2624), .Z(n2751) );
  HS65_LHS_XOR2X3 U2339 ( .A(n2632), .B(n2752), .Z(n1353) );
  HS65_LH_MX41X4 U2340 ( .D0(n2719), .S0(n1008), .D1(n2456), .S1(n2623), .D2(
        n2450), .S2(n2624), .D3(n2447), .S3(n2627), .Z(n2752) );
  HS65_LH_AND2X4 U2341 ( .A(n2753), .B(n2754), .Z(n2718) );
  HS65_LHS_XOR2X3 U2342 ( .A(n2632), .B(n2755), .Z(n1352) );
  HS65_LH_OAI12X2 U2343 ( .A(n2667), .B(n2449), .C(n2756), .Z(n2755) );
  HS65_LH_OAI22X1 U2344 ( .A(n2625), .B(n2757), .C(n2454), .D(n2757), .Z(n2756) );
  HS65_LH_AND2X4 U2345 ( .A(n2450), .B(n2626), .Z(n2757) );
  HS65_LH_NOR2X2 U2346 ( .A(n2753), .B(n2758), .Z(n2721) );
  HS65_LHS_XOR2X3 U2347 ( .A(n2633), .B(n2759), .Z(n1351) );
  HS65_LH_AOI22X1 U2348 ( .A(n2719), .B(n1006), .C(n2456), .D(n2627), .Z(n2759) );
  HS65_LH_NOR3AX2 U2349 ( .A(n2758), .B(n2754), .C(n2753), .Z(n2723) );
  HS65_LHS_XNOR2X3 U2350 ( .A(a[4]), .B(a[3]), .Z(n2758) );
  HS65_LH_NOR2AX3 U2351 ( .A(n2753), .B(n2754), .Z(n2719) );
  HS65_LHS_XNOR2X3 U2352 ( .A(n2632), .B(a[4]), .Z(n2754) );
  HS65_LHS_XOR2X3 U2353 ( .A(n2628), .B(a[3]), .Z(n2753) );
  HS65_LHS_XOR2X3 U2354 ( .A(n2634), .B(n2760), .Z(n1349) );
  HS65_LH_AO22X4 U2355 ( .A(n2565), .B(n2459), .C(n2564), .D(n2762), .Z(n2760)
         );
  HS65_LHS_XOR2X3 U2356 ( .A(n2634), .B(n2763), .Z(n1348) );
  HS65_LH_AO222X4 U2357 ( .A(n2567), .B(n2459), .C(n2563), .D(n2463), .E(n1038), .F(n2461), .Z(n2763) );
  HS65_LHS_XOR2X3 U2358 ( .A(n2634), .B(n2765), .Z(n1347) );
  HS65_LH_MX41X4 U2359 ( .D0(n2461), .S0(n1037), .D1(n2468), .S1(n2564), .D2(
        n2463), .S2(n2566), .D3(n2459), .S3(n2569), .Z(n2765) );
  HS65_LHS_XOR2X3 U2360 ( .A(n2634), .B(n2767), .Z(n1346) );
  HS65_LH_MX41X4 U2361 ( .D0(n2461), .S0(n1036), .D1(n2467), .S1(n2566), .D2(
        n2463), .S2(n2568), .D3(n2459), .S3(n2571), .Z(n2767) );
  HS65_LHS_XOR2X3 U2362 ( .A(n2634), .B(n2768), .Z(n1345) );
  HS65_LH_MX41X4 U2363 ( .D0(n2461), .S0(n1035), .D1(n2467), .S1(n2569), .D2(
        n2463), .S2(n2570), .D3(n2459), .S3(n2573), .Z(n2768) );
  HS65_LHS_XOR2X3 U2364 ( .A(n2634), .B(n2769), .Z(n1344) );
  HS65_LH_MX41X4 U2365 ( .D0(n2461), .S0(n1034), .D1(n2467), .S1(n2571), .D2(
        n2463), .S2(n2572), .D3(n2459), .S3(n2575), .Z(n2769) );
  HS65_LHS_XOR2X3 U2366 ( .A(n2634), .B(n2770), .Z(n1343) );
  HS65_LH_MX41X4 U2367 ( .D0(n2461), .S0(n1033), .D1(n2467), .S1(n2573), .D2(
        n2463), .S2(n2574), .D3(n2459), .S3(n2577), .Z(n2770) );
  HS65_LHS_XOR2X3 U2368 ( .A(n2634), .B(n2771), .Z(n1342) );
  HS65_LH_MX41X4 U2369 ( .D0(n2461), .S0(n1032), .D1(n2467), .S1(n2575), .D2(
        n2463), .S2(n2576), .D3(n2459), .S3(n2579), .Z(n2771) );
  HS65_LHS_XOR2X3 U2370 ( .A(n2634), .B(n2772), .Z(n1341) );
  HS65_LH_MX41X4 U2371 ( .D0(n2461), .S0(n1031), .D1(n2467), .S1(n2577), .D2(
        n2463), .S2(n2578), .D3(n2459), .S3(n2581), .Z(n2772) );
  HS65_LHS_XOR2X3 U2372 ( .A(n2634), .B(n2773), .Z(n1340) );
  HS65_LH_MX41X4 U2373 ( .D0(n2461), .S0(n1030), .D1(n2467), .S1(n2579), .D2(
        n2464), .S2(n2580), .D3(n2459), .S3(n2583), .Z(n2773) );
  HS65_LHS_XOR2X3 U2374 ( .A(n2634), .B(n2774), .Z(n1339) );
  HS65_LH_MX41X4 U2375 ( .D0(n2461), .S0(n1029), .D1(n2467), .S1(n2581), .D2(
        n2463), .S2(n2582), .D3(n2459), .S3(n2585), .Z(n2774) );
  HS65_LHS_XOR2X3 U2376 ( .A(n2634), .B(n2775), .Z(n1338) );
  HS65_LH_MX41X4 U2377 ( .D0(n2461), .S0(n1028), .D1(n2467), .S1(n2583), .D2(
        n2463), .S2(n2584), .D3(n2459), .S3(n2587), .Z(n2775) );
  HS65_LHS_XOR2X3 U2378 ( .A(n2634), .B(n2776), .Z(n1337) );
  HS65_LH_MX41X4 U2379 ( .D0(n2461), .S0(n1027), .D1(n2467), .S1(n2585), .D2(
        n2463), .S2(n2586), .D3(n2459), .S3(n2589), .Z(n2776) );
  HS65_LHS_XOR2X3 U2380 ( .A(n2634), .B(n2777), .Z(n1336) );
  HS65_LH_MX41X4 U2381 ( .D0(n2461), .S0(n1026), .D1(n2467), .S1(n2587), .D2(
        n2464), .S2(n2588), .D3(n2459), .S3(n2591), .Z(n2777) );
  HS65_LHS_XOR2X3 U2382 ( .A(n2634), .B(n2778), .Z(n1335) );
  HS65_LH_MX41X4 U2383 ( .D0(n2461), .S0(n1025), .D1(n2467), .S1(n2589), .D2(
        n2464), .S2(n2590), .D3(n2459), .S3(n2593), .Z(n2778) );
  HS65_LHS_XOR2X3 U2384 ( .A(n2634), .B(n2779), .Z(n1334) );
  HS65_LH_MX41X4 U2385 ( .D0(n2461), .S0(n1024), .D1(n2468), .S1(n2591), .D2(
        n2464), .S2(n2592), .D3(n2459), .S3(n2595), .Z(n2779) );
  HS65_LHS_XOR2X3 U2386 ( .A(n2634), .B(n2780), .Z(n1333) );
  HS65_LH_MX41X4 U2387 ( .D0(n2461), .S0(n1023), .D1(n2468), .S1(n2593), .D2(
        n2464), .S2(n2594), .D3(n2459), .S3(n2597), .Z(n2780) );
  HS65_LHS_XOR2X3 U2388 ( .A(n2634), .B(n2781), .Z(n1332) );
  HS65_LH_MX41X4 U2389 ( .D0(n2461), .S0(n1022), .D1(n2468), .S1(n2595), .D2(
        n2464), .S2(n2596), .D3(n2460), .S3(n2599), .Z(n2781) );
  HS65_LHS_XOR2X3 U2390 ( .A(n2634), .B(n2782), .Z(n1331) );
  HS65_LH_MX41X4 U2391 ( .D0(n2461), .S0(n1021), .D1(n2468), .S1(n2597), .D2(
        n2464), .S2(n2598), .D3(n2460), .S3(n2601), .Z(n2782) );
  HS65_LHS_XOR2X3 U2392 ( .A(n31), .B(n2783), .Z(n1330) );
  HS65_LH_MX41X4 U2393 ( .D0(n2461), .S0(n1020), .D1(n2468), .S1(n2599), .D2(
        n2464), .S2(n2600), .D3(n2460), .S3(n2603), .Z(n2783) );
  HS65_LHS_XOR2X3 U2394 ( .A(n31), .B(n2784), .Z(n1329) );
  HS65_LH_MX41X4 U2395 ( .D0(n2461), .S0(n1019), .D1(n2468), .S1(n2601), .D2(
        n2464), .S2(n2602), .D3(n2460), .S3(n2605), .Z(n2784) );
  HS65_LHS_XOR2X3 U2396 ( .A(n31), .B(n2785), .Z(n1328) );
  HS65_LH_MX41X4 U2397 ( .D0(n2762), .S0(n1018), .D1(n2468), .S1(n2603), .D2(
        n2464), .S2(n2604), .D3(n2460), .S3(n2607), .Z(n2785) );
  HS65_LHS_XOR2X3 U2398 ( .A(n31), .B(n2786), .Z(n1327) );
  HS65_LH_MX41X4 U2399 ( .D0(n2762), .S0(n1017), .D1(n2468), .S1(n2605), .D2(
        n2464), .S2(n2606), .D3(n2460), .S3(n2609), .Z(n2786) );
  HS65_LHS_XOR2X3 U2400 ( .A(n2635), .B(n2787), .Z(n1326) );
  HS65_LH_MX41X4 U2401 ( .D0(n2762), .S0(n1016), .D1(n2468), .S1(n2607), .D2(
        n2464), .S2(n2608), .D3(n2460), .S3(n2611), .Z(n2787) );
  HS65_LHS_XOR2X3 U2402 ( .A(n2635), .B(n2788), .Z(n1325) );
  HS65_LH_MX41X4 U2403 ( .D0(n2762), .S0(n1015), .D1(n2468), .S1(n2609), .D2(
        n2464), .S2(n2610), .D3(n2460), .S3(n2613), .Z(n2788) );
  HS65_LHS_XOR2X3 U2404 ( .A(n2635), .B(n2789), .Z(n1324) );
  HS65_LH_MX41X4 U2405 ( .D0(n2762), .S0(n1014), .D1(n2468), .S1(n2611), .D2(
        n2464), .S2(n2612), .D3(n2460), .S3(n2615), .Z(n2789) );
  HS65_LHS_XOR2X3 U2406 ( .A(n2635), .B(n2790), .Z(n1323) );
  HS65_LH_MX41X4 U2407 ( .D0(n2762), .S0(n1013), .D1(n2468), .S1(n2613), .D2(
        n2465), .S2(n2614), .D3(n2460), .S3(n2617), .Z(n2790) );
  HS65_LHS_XOR2X3 U2408 ( .A(n2635), .B(n2791), .Z(n1322) );
  HS65_LH_MX41X4 U2409 ( .D0(n2762), .S0(n1012), .D1(n2469), .S1(n2615), .D2(
        n2465), .S2(n2616), .D3(n2460), .S3(n2619), .Z(n2791) );
  HS65_LHS_XOR2X3 U2410 ( .A(n2635), .B(n2792), .Z(n1321) );
  HS65_LH_MX41X4 U2411 ( .D0(n2762), .S0(n1011), .D1(n2469), .S1(n2617), .D2(
        n2465), .S2(n2618), .D3(n2460), .S3(n2621), .Z(n2792) );
  HS65_LHS_XOR2X3 U2412 ( .A(n2635), .B(n2793), .Z(n1320) );
  HS65_LH_MX41X4 U2413 ( .D0(n2762), .S0(n1010), .D1(n2469), .S1(n2619), .D2(
        n2465), .S2(n2620), .D3(n2460), .S3(n2623), .Z(n2793) );
  HS65_LHS_XOR2X3 U2414 ( .A(n2635), .B(n2794), .Z(n1319) );
  HS65_LH_MX41X4 U2415 ( .D0(n2762), .S0(n1009), .D1(n2469), .S1(n2621), .D2(
        n2465), .S2(n2622), .D3(n2460), .S3(n2624), .Z(n2794) );
  HS65_LHS_XOR2X3 U2416 ( .A(n2635), .B(n2795), .Z(n1318) );
  HS65_LH_MX41X4 U2417 ( .D0(n2762), .S0(n1008), .D1(n2469), .S1(n2623), .D2(
        n2463), .S2(n2624), .D3(n2460), .S3(n2627), .Z(n2795) );
  HS65_LH_AND2X4 U2418 ( .A(n2796), .B(n2797), .Z(n2761) );
  HS65_LHS_XOR2X3 U2419 ( .A(n2635), .B(n2798), .Z(n1317) );
  HS65_LH_OAI12X2 U2420 ( .A(n2667), .B(n2462), .C(n2799), .Z(n2798) );
  HS65_LH_OAI22X1 U2421 ( .A(n2625), .B(n2800), .C(n2467), .D(n2800), .Z(n2799) );
  HS65_LH_AND2X4 U2422 ( .A(n2463), .B(n2626), .Z(n2800) );
  HS65_LH_NOR2X2 U2423 ( .A(n2796), .B(n2801), .Z(n2764) );
  HS65_LHS_XOR2X3 U2424 ( .A(n2636), .B(n2802), .Z(n1316) );
  HS65_LH_AOI22X1 U2425 ( .A(n2762), .B(n1006), .C(n2469), .D(n2627), .Z(n2802) );
  HS65_LH_NOR3AX2 U2426 ( .A(n2801), .B(n2797), .C(n2796), .Z(n2766) );
  HS65_LHS_XNOR2X3 U2427 ( .A(a[7]), .B(a[6]), .Z(n2801) );
  HS65_LH_NOR2AX3 U2428 ( .A(n2796), .B(n2797), .Z(n2762) );
  HS65_LHS_XNOR2X3 U2429 ( .A(n2635), .B(a[7]), .Z(n2797) );
  HS65_LHS_XOR2X3 U2430 ( .A(n2631), .B(a[6]), .Z(n2796) );
  HS65_LHS_XOR2X3 U2431 ( .A(n2637), .B(n2803), .Z(n1314) );
  HS65_LH_AO22X4 U2432 ( .A(n2565), .B(n2472), .C(n2564), .D(n2805), .Z(n2803)
         );
  HS65_LHS_XOR2X3 U2433 ( .A(n2637), .B(n2806), .Z(n1313) );
  HS65_LH_AO222X4 U2434 ( .A(n2567), .B(n2472), .C(n2563), .D(n2476), .E(n1038), .F(n2474), .Z(n2806) );
  HS65_LHS_XOR2X3 U2435 ( .A(n2637), .B(n2808), .Z(n1312) );
  HS65_LH_MX41X4 U2436 ( .D0(n2474), .S0(n1037), .D1(n2472), .S1(n2569), .D2(
        n2477), .S2(n2566), .D3(n2481), .S3(n2564), .Z(n2808) );
  HS65_LHS_XOR2X3 U2437 ( .A(n2637), .B(n2810), .Z(n1311) );
  HS65_LH_MX41X4 U2438 ( .D0(n2474), .S0(n1036), .D1(n2472), .S1(n2571), .D2(
        n2476), .S2(n2568), .D3(n2480), .S3(n2566), .Z(n2810) );
  HS65_LHS_XOR2X3 U2439 ( .A(n2637), .B(n2811), .Z(n1310) );
  HS65_LH_MX41X4 U2440 ( .D0(n2474), .S0(n1035), .D1(n2472), .S1(n2573), .D2(
        n2476), .S2(n2570), .D3(n2480), .S3(n2569), .Z(n2811) );
  HS65_LHS_XOR2X3 U2441 ( .A(n2637), .B(n2812), .Z(n1309) );
  HS65_LH_MX41X4 U2442 ( .D0(n2474), .S0(n1034), .D1(n2472), .S1(n2575), .D2(
        n2476), .S2(n2572), .D3(n2480), .S3(n2571), .Z(n2812) );
  HS65_LHS_XOR2X3 U2443 ( .A(n2637), .B(n2813), .Z(n1308) );
  HS65_LH_MX41X4 U2444 ( .D0(n2474), .S0(n1033), .D1(n2472), .S1(n2577), .D2(
        n2476), .S2(n2574), .D3(n2480), .S3(n2573), .Z(n2813) );
  HS65_LHS_XOR2X3 U2445 ( .A(n2637), .B(n2814), .Z(n1307) );
  HS65_LH_MX41X4 U2446 ( .D0(n2474), .S0(n1032), .D1(n2472), .S1(n2579), .D2(
        n2476), .S2(n2576), .D3(n2480), .S3(n2575), .Z(n2814) );
  HS65_LHS_XOR2X3 U2447 ( .A(n2637), .B(n2815), .Z(n1306) );
  HS65_LH_MX41X4 U2448 ( .D0(n2474), .S0(n1031), .D1(n2472), .S1(n2581), .D2(
        n2476), .S2(n2578), .D3(n2480), .S3(n2577), .Z(n2815) );
  HS65_LHS_XOR2X3 U2449 ( .A(n2637), .B(n2816), .Z(n1305) );
  HS65_LH_MX41X4 U2450 ( .D0(n2474), .S0(n1030), .D1(n2472), .S1(n2583), .D2(
        n2477), .S2(n2580), .D3(n2480), .S3(n2579), .Z(n2816) );
  HS65_LHS_XOR2X3 U2451 ( .A(n2637), .B(n2817), .Z(n1304) );
  HS65_LH_MX41X4 U2452 ( .D0(n2474), .S0(n1029), .D1(n2472), .S1(n2585), .D2(
        n2476), .S2(n2582), .D3(n2480), .S3(n2581), .Z(n2817) );
  HS65_LHS_XOR2X3 U2453 ( .A(n2637), .B(n2818), .Z(n1303) );
  HS65_LH_MX41X4 U2454 ( .D0(n2474), .S0(n1028), .D1(n2472), .S1(n2587), .D2(
        n2477), .S2(n2584), .D3(n2480), .S3(n2583), .Z(n2818) );
  HS65_LHS_XOR2X3 U2455 ( .A(n2637), .B(n2819), .Z(n1302) );
  HS65_LH_MX41X4 U2456 ( .D0(n2474), .S0(n1027), .D1(n2472), .S1(n2589), .D2(
        n2477), .S2(n2586), .D3(n2480), .S3(n2585), .Z(n2819) );
  HS65_LHS_XOR2X3 U2457 ( .A(n2637), .B(n2820), .Z(n1301) );
  HS65_LH_MX41X4 U2458 ( .D0(n2474), .S0(n1026), .D1(n2472), .S1(n2591), .D2(
        n2477), .S2(n2588), .D3(n2480), .S3(n2587), .Z(n2820) );
  HS65_LHS_XOR2X3 U2459 ( .A(n2637), .B(n2821), .Z(n1300) );
  HS65_LH_MX41X4 U2460 ( .D0(n2474), .S0(n1025), .D1(n2472), .S1(n2593), .D2(
        n2477), .S2(n2590), .D3(n2480), .S3(n2589), .Z(n2821) );
  HS65_LHS_XOR2X3 U2461 ( .A(n2637), .B(n2822), .Z(n1299) );
  HS65_LH_MX41X4 U2462 ( .D0(n2474), .S0(n1024), .D1(n2476), .S1(n2593), .D2(
        n2473), .S2(n2594), .D3(n2481), .S3(n2591), .Z(n2822) );
  HS65_LHS_XOR2X3 U2463 ( .A(n2637), .B(n2823), .Z(n1298) );
  HS65_LH_MX41X4 U2464 ( .D0(n2474), .S0(n1023), .D1(n2476), .S1(n2595), .D2(
        n2473), .S2(n2596), .D3(n2481), .S3(n2593), .Z(n2823) );
  HS65_LHS_XOR2X3 U2465 ( .A(n2637), .B(n2824), .Z(n1297) );
  HS65_LH_MX41X4 U2466 ( .D0(n2474), .S0(n1022), .D1(n2473), .S1(n2599), .D2(
        n2477), .S2(n2596), .D3(n2481), .S3(n2595), .Z(n2824) );
  HS65_LHS_XOR2X3 U2467 ( .A(n2637), .B(n2825), .Z(n1296) );
  HS65_LH_MX41X4 U2468 ( .D0(n2474), .S0(n1021), .D1(n2473), .S1(n2601), .D2(
        n2477), .S2(n2598), .D3(n2481), .S3(n2597), .Z(n2825) );
  HS65_LHS_XOR2X3 U2469 ( .A(n43), .B(n2826), .Z(n1295) );
  HS65_LH_MX41X4 U2470 ( .D0(n2474), .S0(n1020), .D1(n2472), .S1(n2603), .D2(
        n2477), .S2(n2600), .D3(n2481), .S3(n2599), .Z(n2826) );
  HS65_LHS_XOR2X3 U2471 ( .A(n43), .B(n2827), .Z(n1294) );
  HS65_LH_MX41X4 U2472 ( .D0(n2474), .S0(n1019), .D1(n2473), .S1(n2605), .D2(
        n2477), .S2(n2602), .D3(n2481), .S3(n2601), .Z(n2827) );
  HS65_LHS_XOR2X3 U2473 ( .A(n43), .B(n2828), .Z(n1293) );
  HS65_LH_MX41X4 U2474 ( .D0(n2805), .S0(n1018), .D1(n2473), .S1(n2607), .D2(
        n2477), .S2(n2604), .D3(n2481), .S3(n2603), .Z(n2828) );
  HS65_LHS_XOR2X3 U2475 ( .A(n43), .B(n2829), .Z(n1292) );
  HS65_LH_MX41X4 U2476 ( .D0(n2805), .S0(n1017), .D1(n2473), .S1(n2609), .D2(
        n2477), .S2(n2606), .D3(n2481), .S3(n2605), .Z(n2829) );
  HS65_LHS_XOR2X3 U2477 ( .A(n2638), .B(n2830), .Z(n1291) );
  HS65_LH_MX41X4 U2478 ( .D0(n2805), .S0(n1016), .D1(n2473), .S1(n2611), .D2(
        n2477), .S2(n2608), .D3(n2481), .S3(n2607), .Z(n2830) );
  HS65_LHS_XOR2X3 U2479 ( .A(n2638), .B(n2831), .Z(n1290) );
  HS65_LH_MX41X4 U2480 ( .D0(n2805), .S0(n1015), .D1(n2473), .S1(n2613), .D2(
        n2477), .S2(n2610), .D3(n2481), .S3(n2609), .Z(n2831) );
  HS65_LHS_XOR2X3 U2481 ( .A(n2638), .B(n2832), .Z(n1289) );
  HS65_LH_MX41X4 U2482 ( .D0(n2805), .S0(n1014), .D1(n2473), .S1(n2615), .D2(
        n2478), .S2(n2612), .D3(n2481), .S3(n2611), .Z(n2832) );
  HS65_LHS_XOR2X3 U2483 ( .A(n2638), .B(n2833), .Z(n1288) );
  HS65_LH_MX41X4 U2484 ( .D0(n2805), .S0(n1013), .D1(n2473), .S1(n2617), .D2(
        n2478), .S2(n2614), .D3(n2481), .S3(n2613), .Z(n2833) );
  HS65_LHS_XOR2X3 U2485 ( .A(n2638), .B(n2834), .Z(n1287) );
  HS65_LH_MX41X4 U2486 ( .D0(n2805), .S0(n1012), .D1(n2473), .S1(n2619), .D2(
        n2478), .S2(n2616), .D3(n2482), .S3(n2615), .Z(n2834) );
  HS65_LHS_XOR2X3 U2487 ( .A(n2638), .B(n2835), .Z(n1286) );
  HS65_LH_MX41X4 U2488 ( .D0(n2805), .S0(n1011), .D1(n2473), .S1(n2621), .D2(
        n2478), .S2(n2618), .D3(n2482), .S3(n2617), .Z(n2835) );
  HS65_LHS_XOR2X3 U2489 ( .A(n2638), .B(n2836), .Z(n1285) );
  HS65_LH_MX41X4 U2490 ( .D0(n2805), .S0(n1010), .D1(n2473), .S1(n2623), .D2(
        n2478), .S2(n2620), .D3(n2482), .S3(n2619), .Z(n2836) );
  HS65_LHS_XOR2X3 U2491 ( .A(n2638), .B(n2837), .Z(n1284) );
  HS65_LH_MX41X4 U2492 ( .D0(n2805), .S0(n1009), .D1(n2473), .S1(n2624), .D2(
        n2476), .S2(n2622), .D3(n2482), .S3(n2621), .Z(n2837) );
  HS65_LHS_XOR2X3 U2493 ( .A(n2638), .B(n2838), .Z(n1283) );
  HS65_LH_MX41X4 U2494 ( .D0(n2805), .S0(n1008), .D1(n2476), .S1(n2624), .D2(
        n2473), .S2(n2626), .D3(n2482), .S3(n2623), .Z(n2838) );
  HS65_LH_AND2X4 U2495 ( .A(n2839), .B(n2840), .Z(n2804) );
  HS65_LHS_XOR2X3 U2496 ( .A(n2638), .B(n2841), .Z(n1282) );
  HS65_LH_OAI12X2 U2497 ( .A(n2667), .B(n2475), .C(n2842), .Z(n2841) );
  HS65_LH_OAI22X1 U2498 ( .A(n2625), .B(n2843), .C(n2480), .D(n2843), .Z(n2842) );
  HS65_LH_AND2X4 U2499 ( .A(n2476), .B(n2626), .Z(n2843) );
  HS65_LH_NOR2X2 U2500 ( .A(n2839), .B(n2844), .Z(n2807) );
  HS65_LHS_XOR2X3 U2501 ( .A(n2639), .B(n2845), .Z(n1281) );
  HS65_LH_AOI22X1 U2502 ( .A(n2805), .B(n1006), .C(n2482), .D(n2627), .Z(n2845) );
  HS65_LH_NOR3AX2 U2503 ( .A(n2844), .B(n2840), .C(n2839), .Z(n2809) );
  HS65_LHS_XNOR2X3 U2504 ( .A(a[9]), .B(a[10]), .Z(n2844) );
  HS65_LH_NOR2AX3 U2505 ( .A(n2839), .B(n2840), .Z(n2805) );
  HS65_LHS_XNOR2X3 U2506 ( .A(n2638), .B(a[10]), .Z(n2840) );
  HS65_LHS_XOR2X3 U2507 ( .A(n2634), .B(a[9]), .Z(n2839) );
  HS65_LHS_XOR2X3 U2508 ( .A(n2640), .B(n2846), .Z(n1279) );
  HS65_LH_AO22X4 U2509 ( .A(n2565), .B(n2485), .C(n2564), .D(n2848), .Z(n2846)
         );
  HS65_LHS_XOR2X3 U2510 ( .A(n2640), .B(n2849), .Z(n1278) );
  HS65_LH_AO222X4 U2511 ( .A(n2567), .B(n2485), .C(n2563), .D(n2489), .E(n1038), .F(n2487), .Z(n2849) );
  HS65_LHS_XOR2X3 U2512 ( .A(n2640), .B(n2851), .Z(n1277) );
  HS65_LH_MX41X4 U2513 ( .D0(n2487), .S0(n1037), .D1(n2494), .S1(n2563), .D2(
        n2489), .S2(n2566), .D3(n2485), .S3(n2569), .Z(n2851) );
  HS65_LHS_XOR2X3 U2514 ( .A(n2640), .B(n2853), .Z(n1276) );
  HS65_LH_MX41X4 U2515 ( .D0(n2487), .S0(n1036), .D1(n2493), .S1(n2566), .D2(
        n2489), .S2(n2568), .D3(n2485), .S3(n2571), .Z(n2853) );
  HS65_LHS_XOR2X3 U2516 ( .A(n2640), .B(n2854), .Z(n1275) );
  HS65_LH_MX41X4 U2517 ( .D0(n2487), .S0(n1035), .D1(n2493), .S1(n2569), .D2(
        n2489), .S2(n2570), .D3(n2485), .S3(n2573), .Z(n2854) );
  HS65_LHS_XOR2X3 U2518 ( .A(n2640), .B(n2855), .Z(n1274) );
  HS65_LH_MX41X4 U2519 ( .D0(n2487), .S0(n1034), .D1(n2493), .S1(n2571), .D2(
        n2489), .S2(n2572), .D3(n2485), .S3(n2575), .Z(n2855) );
  HS65_LHS_XOR2X3 U2520 ( .A(n2640), .B(n2856), .Z(n1273) );
  HS65_LH_MX41X4 U2521 ( .D0(n2487), .S0(n1033), .D1(n2493), .S1(n2573), .D2(
        n2489), .S2(n2574), .D3(n2485), .S3(n2577), .Z(n2856) );
  HS65_LHS_XOR2X3 U2522 ( .A(n2640), .B(n2857), .Z(n1272) );
  HS65_LH_MX41X4 U2523 ( .D0(n2487), .S0(n1032), .D1(n2493), .S1(n2575), .D2(
        n2489), .S2(n2576), .D3(n2485), .S3(n2579), .Z(n2857) );
  HS65_LHS_XOR2X3 U2524 ( .A(n2640), .B(n2858), .Z(n1271) );
  HS65_LH_MX41X4 U2525 ( .D0(n2487), .S0(n1031), .D1(n2493), .S1(n2577), .D2(
        n2489), .S2(n2578), .D3(n2485), .S3(n2581), .Z(n2858) );
  HS65_LHS_XOR2X3 U2526 ( .A(n2640), .B(n2859), .Z(n1270) );
  HS65_LH_MX41X4 U2527 ( .D0(n2487), .S0(n1030), .D1(n2493), .S1(n2579), .D2(
        n2490), .S2(n2580), .D3(n2485), .S3(n2583), .Z(n2859) );
  HS65_LHS_XOR2X3 U2528 ( .A(n2640), .B(n2860), .Z(n1269) );
  HS65_LH_MX41X4 U2529 ( .D0(n2487), .S0(n1029), .D1(n2493), .S1(n2581), .D2(
        n2489), .S2(n2582), .D3(n2485), .S3(n2585), .Z(n2860) );
  HS65_LHS_XOR2X3 U2530 ( .A(n2640), .B(n2861), .Z(n1268) );
  HS65_LH_MX41X4 U2531 ( .D0(n2487), .S0(n1028), .D1(n2493), .S1(n2583), .D2(
        n2489), .S2(n2584), .D3(n2485), .S3(n2587), .Z(n2861) );
  HS65_LHS_XOR2X3 U2532 ( .A(n2640), .B(n2862), .Z(n1267) );
  HS65_LH_MX41X4 U2533 ( .D0(n2487), .S0(n1027), .D1(n2493), .S1(n2585), .D2(
        n2489), .S2(n2586), .D3(n2485), .S3(n2589), .Z(n2862) );
  HS65_LHS_XOR2X3 U2534 ( .A(n2640), .B(n2863), .Z(n1266) );
  HS65_LH_MX41X4 U2535 ( .D0(n2487), .S0(n1026), .D1(n2493), .S1(n2587), .D2(
        n2490), .S2(n2588), .D3(n2485), .S3(n2591), .Z(n2863) );
  HS65_LHS_XOR2X3 U2536 ( .A(n2640), .B(n2864), .Z(n1265) );
  HS65_LH_MX41X4 U2537 ( .D0(n2487), .S0(n1025), .D1(n2493), .S1(n2589), .D2(
        n2490), .S2(n2590), .D3(n2485), .S3(n2593), .Z(n2864) );
  HS65_LHS_XOR2X3 U2538 ( .A(n2640), .B(n2865), .Z(n1264) );
  HS65_LH_MX41X4 U2539 ( .D0(n2487), .S0(n1024), .D1(n2494), .S1(n2591), .D2(
        n2490), .S2(n2592), .D3(n2485), .S3(n2595), .Z(n2865) );
  HS65_LHS_XOR2X3 U2540 ( .A(n2640), .B(n2866), .Z(n1263) );
  HS65_LH_MX41X4 U2541 ( .D0(n2487), .S0(n1023), .D1(n2494), .S1(n2593), .D2(
        n2490), .S2(n2594), .D3(n2485), .S3(n2597), .Z(n2866) );
  HS65_LHS_XOR2X3 U2542 ( .A(n2640), .B(n2867), .Z(n1262) );
  HS65_LH_MX41X4 U2543 ( .D0(n2487), .S0(n1022), .D1(n2494), .S1(n2595), .D2(
        n2490), .S2(n2596), .D3(n2486), .S3(n2599), .Z(n2867) );
  HS65_LHS_XOR2X3 U2544 ( .A(n2640), .B(n2868), .Z(n1261) );
  HS65_LH_MX41X4 U2545 ( .D0(n2487), .S0(n1021), .D1(n2494), .S1(n2597), .D2(
        n2490), .S2(n2598), .D3(n2486), .S3(n2601), .Z(n2868) );
  HS65_LHS_XOR2X3 U2546 ( .A(n55), .B(n2869), .Z(n1260) );
  HS65_LH_MX41X4 U2547 ( .D0(n2487), .S0(n1020), .D1(n2494), .S1(n2599), .D2(
        n2490), .S2(n2600), .D3(n2486), .S3(n2603), .Z(n2869) );
  HS65_LHS_XOR2X3 U2548 ( .A(n55), .B(n2870), .Z(n1259) );
  HS65_LH_MX41X4 U2549 ( .D0(n2487), .S0(n1019), .D1(n2494), .S1(n2601), .D2(
        n2490), .S2(n2602), .D3(n2486), .S3(n2605), .Z(n2870) );
  HS65_LHS_XOR2X3 U2550 ( .A(n55), .B(n2871), .Z(n1258) );
  HS65_LH_MX41X4 U2551 ( .D0(n2848), .S0(n1018), .D1(n2494), .S1(n2603), .D2(
        n2490), .S2(n2604), .D3(n2486), .S3(n2607), .Z(n2871) );
  HS65_LHS_XOR2X3 U2552 ( .A(n55), .B(n2872), .Z(n1257) );
  HS65_LH_MX41X4 U2553 ( .D0(n2848), .S0(n1017), .D1(n2494), .S1(n2605), .D2(
        n2490), .S2(n2606), .D3(n2486), .S3(n2609), .Z(n2872) );
  HS65_LHS_XOR2X3 U2554 ( .A(n2641), .B(n2873), .Z(n1256) );
  HS65_LH_MX41X4 U2555 ( .D0(n2848), .S0(n1016), .D1(n2494), .S1(n2607), .D2(
        n2490), .S2(n2608), .D3(n2486), .S3(n2611), .Z(n2873) );
  HS65_LHS_XOR2X3 U2556 ( .A(n2641), .B(n2874), .Z(n1255) );
  HS65_LH_MX41X4 U2557 ( .D0(n2848), .S0(n1015), .D1(n2494), .S1(n2609), .D2(
        n2490), .S2(n2610), .D3(n2486), .S3(n2613), .Z(n2874) );
  HS65_LHS_XOR2X3 U2558 ( .A(n2641), .B(n2875), .Z(n1254) );
  HS65_LH_MX41X4 U2559 ( .D0(n2848), .S0(n1014), .D1(n2494), .S1(n2611), .D2(
        n2490), .S2(n2612), .D3(n2486), .S3(n2615), .Z(n2875) );
  HS65_LHS_XOR2X3 U2560 ( .A(n2641), .B(n2876), .Z(n1253) );
  HS65_LH_MX41X4 U2561 ( .D0(n2848), .S0(n1013), .D1(n2494), .S1(n2613), .D2(
        n2491), .S2(n2614), .D3(n2486), .S3(n2617), .Z(n2876) );
  HS65_LHS_XOR2X3 U2562 ( .A(n2641), .B(n2877), .Z(n1252) );
  HS65_LH_MX41X4 U2563 ( .D0(n2848), .S0(n1012), .D1(n2495), .S1(n2615), .D2(
        n2491), .S2(n2616), .D3(n2486), .S3(n2619), .Z(n2877) );
  HS65_LHS_XOR2X3 U2564 ( .A(n2641), .B(n2878), .Z(n1251) );
  HS65_LH_MX41X4 U2565 ( .D0(n2848), .S0(n1011), .D1(n2495), .S1(n2617), .D2(
        n2491), .S2(n2618), .D3(n2486), .S3(n2621), .Z(n2878) );
  HS65_LHS_XOR2X3 U2566 ( .A(n2641), .B(n2879), .Z(n1250) );
  HS65_LH_MX41X4 U2567 ( .D0(n2848), .S0(n1010), .D1(n2495), .S1(n2619), .D2(
        n2491), .S2(n2620), .D3(n2486), .S3(n2623), .Z(n2879) );
  HS65_LHS_XOR2X3 U2568 ( .A(n2641), .B(n2880), .Z(n1249) );
  HS65_LH_MX41X4 U2569 ( .D0(n2848), .S0(n1009), .D1(n2495), .S1(n2621), .D2(
        n2491), .S2(n2622), .D3(n2486), .S3(n2624), .Z(n2880) );
  HS65_LHS_XOR2X3 U2570 ( .A(n2641), .B(n2881), .Z(n1248) );
  HS65_LH_MX41X4 U2571 ( .D0(n2848), .S0(n1008), .D1(n2495), .S1(n2623), .D2(
        n2489), .S2(n2624), .D3(n2486), .S3(n2627), .Z(n2881) );
  HS65_LH_AND2X4 U2572 ( .A(n2882), .B(n2883), .Z(n2847) );
  HS65_LHS_XOR2X3 U2573 ( .A(n2641), .B(n2884), .Z(n1247) );
  HS65_LH_OAI12X2 U2574 ( .A(n2667), .B(n2488), .C(n2885), .Z(n2884) );
  HS65_LH_OAI22X1 U2575 ( .A(n2625), .B(n2886), .C(n2493), .D(n2886), .Z(n2885) );
  HS65_LH_AND2X4 U2576 ( .A(n2489), .B(n2626), .Z(n2886) );
  HS65_LH_NOR2X2 U2577 ( .A(n2882), .B(n2887), .Z(n2850) );
  HS65_LHS_XOR2X3 U2578 ( .A(n2642), .B(n2888), .Z(n1246) );
  HS65_LH_AOI22X1 U2579 ( .A(n2848), .B(n1006), .C(n2495), .D(n2627), .Z(n2888) );
  HS65_LH_NOR3AX2 U2580 ( .A(n2887), .B(n2883), .C(n2882), .Z(n2852) );
  HS65_LHS_XNOR2X3 U2581 ( .A(a[13]), .B(a[12]), .Z(n2887) );
  HS65_LH_NOR2AX3 U2582 ( .A(n2882), .B(n2883), .Z(n2848) );
  HS65_LHS_XNOR2X3 U2583 ( .A(n2641), .B(a[13]), .Z(n2883) );
  HS65_LHS_XOR2X3 U2584 ( .A(n2637), .B(a[12]), .Z(n2882) );
  HS65_LHS_XOR2X3 U2585 ( .A(n2643), .B(n2889), .Z(n1244) );
  HS65_LH_AO22X4 U2586 ( .A(n2564), .B(n2498), .C(n2564), .D(n2891), .Z(n2889)
         );
  HS65_LHS_XOR2X3 U2587 ( .A(n2643), .B(n2892), .Z(n1243) );
  HS65_LH_AO222X4 U2588 ( .A(n2567), .B(n2498), .C(n2563), .D(n2502), .E(n1038), .F(n2500), .Z(n2892) );
  HS65_LHS_XOR2X3 U2589 ( .A(n2643), .B(n2894), .Z(n1242) );
  HS65_LH_MX41X4 U2590 ( .D0(n2500), .S0(n1037), .D1(n2507), .S1(n2563), .D2(
        n2502), .S2(n2566), .D3(n2498), .S3(n2569), .Z(n2894) );
  HS65_LHS_XOR2X3 U2591 ( .A(n2643), .B(n2896), .Z(n1241) );
  HS65_LH_MX41X4 U2592 ( .D0(n2500), .S0(n1036), .D1(n2506), .S1(n2566), .D2(
        n2502), .S2(n2568), .D3(n2498), .S3(n2571), .Z(n2896) );
  HS65_LHS_XOR2X3 U2593 ( .A(n2643), .B(n2897), .Z(n1240) );
  HS65_LH_MX41X4 U2594 ( .D0(n2500), .S0(n1035), .D1(n2506), .S1(n2568), .D2(
        n2502), .S2(n2570), .D3(n2498), .S3(n2573), .Z(n2897) );
  HS65_LHS_XOR2X3 U2595 ( .A(n2643), .B(n2898), .Z(n1239) );
  HS65_LH_MX41X4 U2596 ( .D0(n2500), .S0(n1034), .D1(n2506), .S1(n2570), .D2(
        n2502), .S2(n2572), .D3(n2498), .S3(n2575), .Z(n2898) );
  HS65_LHS_XOR2X3 U2597 ( .A(n2643), .B(n2899), .Z(n1238) );
  HS65_LH_MX41X4 U2598 ( .D0(n2500), .S0(n1033), .D1(n2506), .S1(n2572), .D2(
        n2502), .S2(n2574), .D3(n2498), .S3(n2577), .Z(n2899) );
  HS65_LHS_XOR2X3 U2599 ( .A(n2643), .B(n2900), .Z(n1237) );
  HS65_LH_MX41X4 U2600 ( .D0(n2500), .S0(n1032), .D1(n2506), .S1(n2574), .D2(
        n2502), .S2(n2576), .D3(n2498), .S3(n2579), .Z(n2900) );
  HS65_LHS_XOR2X3 U2601 ( .A(n2643), .B(n2901), .Z(n1236) );
  HS65_LH_MX41X4 U2602 ( .D0(n2500), .S0(n1031), .D1(n2506), .S1(n2576), .D2(
        n2502), .S2(n2578), .D3(n2498), .S3(n2581), .Z(n2901) );
  HS65_LHS_XOR2X3 U2603 ( .A(n2643), .B(n2902), .Z(n1235) );
  HS65_LH_MX41X4 U2604 ( .D0(n2500), .S0(n1030), .D1(n2506), .S1(n2578), .D2(
        n2503), .S2(n2580), .D3(n2498), .S3(n2583), .Z(n2902) );
  HS65_LHS_XOR2X3 U2605 ( .A(n2643), .B(n2903), .Z(n1234) );
  HS65_LH_MX41X4 U2606 ( .D0(n2500), .S0(n1029), .D1(n2506), .S1(n2580), .D2(
        n2502), .S2(n2582), .D3(n2498), .S3(n2585), .Z(n2903) );
  HS65_LHS_XOR2X3 U2607 ( .A(n2643), .B(n2904), .Z(n1233) );
  HS65_LH_MX41X4 U2608 ( .D0(n2500), .S0(n1028), .D1(n2506), .S1(n2582), .D2(
        n2502), .S2(n2584), .D3(n2498), .S3(n2587), .Z(n2904) );
  HS65_LHS_XOR2X3 U2609 ( .A(n2643), .B(n2905), .Z(n1232) );
  HS65_LH_MX41X4 U2610 ( .D0(n2500), .S0(n1027), .D1(n2506), .S1(n2584), .D2(
        n2502), .S2(n2586), .D3(n2498), .S3(n2589), .Z(n2905) );
  HS65_LHS_XOR2X3 U2611 ( .A(n2643), .B(n2906), .Z(n1231) );
  HS65_LH_MX41X4 U2612 ( .D0(n2500), .S0(n1026), .D1(n2506), .S1(n2586), .D2(
        n2503), .S2(n2588), .D3(n2498), .S3(n2591), .Z(n2906) );
  HS65_LHS_XOR2X3 U2613 ( .A(n2643), .B(n2907), .Z(n1230) );
  HS65_LH_MX41X4 U2614 ( .D0(n2500), .S0(n1025), .D1(n2506), .S1(n2589), .D2(
        n2503), .S2(n2590), .D3(n2498), .S3(n2593), .Z(n2907) );
  HS65_LHS_XOR2X3 U2615 ( .A(n2643), .B(n2908), .Z(n1229) );
  HS65_LH_MX41X4 U2616 ( .D0(n2500), .S0(n1024), .D1(n2507), .S1(n2591), .D2(
        n2503), .S2(n2592), .D3(n2498), .S3(n2595), .Z(n2908) );
  HS65_LHS_XOR2X3 U2617 ( .A(n2643), .B(n2909), .Z(n1228) );
  HS65_LH_MX41X4 U2618 ( .D0(n2500), .S0(n1023), .D1(n2507), .S1(n2593), .D2(
        n2503), .S2(n2594), .D3(n2498), .S3(n2597), .Z(n2909) );
  HS65_LHS_XOR2X3 U2619 ( .A(n2643), .B(n2910), .Z(n1227) );
  HS65_LH_MX41X4 U2620 ( .D0(n2500), .S0(n1022), .D1(n2507), .S1(n2594), .D2(
        n2503), .S2(n2596), .D3(n2499), .S3(n2599), .Z(n2910) );
  HS65_LHS_XOR2X3 U2621 ( .A(n2643), .B(n2911), .Z(n1226) );
  HS65_LH_MX41X4 U2622 ( .D0(n2500), .S0(n1021), .D1(n2507), .S1(n2597), .D2(
        n2503), .S2(n2598), .D3(n2499), .S3(n2601), .Z(n2911) );
  HS65_LHS_XOR2X3 U2623 ( .A(n67), .B(n2912), .Z(n1225) );
  HS65_LH_MX41X4 U2624 ( .D0(n2500), .S0(n1020), .D1(n2507), .S1(n2598), .D2(
        n2503), .S2(n2600), .D3(n2499), .S3(n2603), .Z(n2912) );
  HS65_LHS_XOR2X3 U2625 ( .A(n67), .B(n2913), .Z(n1224) );
  HS65_LH_MX41X4 U2626 ( .D0(n2500), .S0(n1019), .D1(n2507), .S1(n2601), .D2(
        n2503), .S2(n2602), .D3(n2499), .S3(n2605), .Z(n2913) );
  HS65_LHS_XOR2X3 U2627 ( .A(n67), .B(n2914), .Z(n1223) );
  HS65_LH_MX41X4 U2628 ( .D0(n2891), .S0(n1018), .D1(n2507), .S1(n2603), .D2(
        n2503), .S2(n2604), .D3(n2499), .S3(n2607), .Z(n2914) );
  HS65_LHS_XOR2X3 U2629 ( .A(n67), .B(n2915), .Z(n1222) );
  HS65_LH_MX41X4 U2630 ( .D0(n2891), .S0(n1017), .D1(n2507), .S1(n2605), .D2(
        n2503), .S2(n2606), .D3(n2499), .S3(n2609), .Z(n2915) );
  HS65_LHS_XOR2X3 U2631 ( .A(n2644), .B(n2916), .Z(n1221) );
  HS65_LH_MX41X4 U2632 ( .D0(n2891), .S0(n1016), .D1(n2507), .S1(n2606), .D2(
        n2503), .S2(n2608), .D3(n2499), .S3(n2611), .Z(n2916) );
  HS65_LHS_XOR2X3 U2633 ( .A(n2644), .B(n2917), .Z(n1220) );
  HS65_LH_MX41X4 U2634 ( .D0(n2891), .S0(n1015), .D1(n2507), .S1(n2608), .D2(
        n2503), .S2(n2610), .D3(n2499), .S3(n2613), .Z(n2917) );
  HS65_LHS_XOR2X3 U2635 ( .A(n2644), .B(n2918), .Z(n1219) );
  HS65_LH_MX41X4 U2636 ( .D0(n2891), .S0(n1014), .D1(n2507), .S1(n2610), .D2(
        n2503), .S2(n2612), .D3(n2499), .S3(n2615), .Z(n2918) );
  HS65_LHS_XOR2X3 U2637 ( .A(n2644), .B(n2919), .Z(n1218) );
  HS65_LH_MX41X4 U2638 ( .D0(n2891), .S0(n1013), .D1(n2507), .S1(n2613), .D2(
        n2504), .S2(n2614), .D3(n2499), .S3(n2617), .Z(n2919) );
  HS65_LHS_XOR2X3 U2639 ( .A(n2644), .B(n2920), .Z(n1217) );
  HS65_LH_MX41X4 U2640 ( .D0(n2891), .S0(n1012), .D1(n2508), .S1(n2615), .D2(
        n2504), .S2(n2616), .D3(n2499), .S3(n2619), .Z(n2920) );
  HS65_LHS_XOR2X3 U2641 ( .A(n2644), .B(n2921), .Z(n1216) );
  HS65_LH_MX41X4 U2642 ( .D0(n2891), .S0(n1011), .D1(n2508), .S1(n2617), .D2(
        n2504), .S2(n2618), .D3(n2499), .S3(n2621), .Z(n2921) );
  HS65_LHS_XOR2X3 U2643 ( .A(n2644), .B(n2922), .Z(n1215) );
  HS65_LH_MX41X4 U2644 ( .D0(n2891), .S0(n1010), .D1(n2508), .S1(n2618), .D2(
        n2504), .S2(n2620), .D3(n2499), .S3(n2623), .Z(n2922) );
  HS65_LHS_XOR2X3 U2645 ( .A(n2644), .B(n2923), .Z(n1214) );
  HS65_LH_MX41X4 U2646 ( .D0(n2891), .S0(n1009), .D1(n2508), .S1(n2620), .D2(
        n2504), .S2(n2622), .D3(n2499), .S3(n2624), .Z(n2923) );
  HS65_LHS_XOR2X3 U2647 ( .A(n2644), .B(n2924), .Z(n1213) );
  HS65_LH_MX41X4 U2648 ( .D0(n2891), .S0(n1008), .D1(n2508), .S1(n2622), .D2(
        n2502), .S2(n2624), .D3(n2499), .S3(n2626), .Z(n2924) );
  HS65_LH_AND2X4 U2649 ( .A(n2925), .B(n2926), .Z(n2890) );
  HS65_LHS_XOR2X3 U2650 ( .A(n2644), .B(n2927), .Z(n1212) );
  HS65_LH_OAI12X2 U2651 ( .A(n2667), .B(n2501), .C(n2928), .Z(n2927) );
  HS65_LH_OAI22X1 U2652 ( .A(n2625), .B(n2929), .C(n2506), .D(n2929), .Z(n2928) );
  HS65_LH_AND2X4 U2653 ( .A(n2502), .B(n2626), .Z(n2929) );
  HS65_LH_NOR2X2 U2654 ( .A(n2925), .B(n2930), .Z(n2893) );
  HS65_LHS_XOR2X3 U2655 ( .A(n2645), .B(n2931), .Z(n1211) );
  HS65_LH_AOI22X1 U2656 ( .A(n2891), .B(n1006), .C(n2508), .D(n2627), .Z(n2931) );
  HS65_LH_NOR3AX2 U2657 ( .A(n2930), .B(n2926), .C(n2925), .Z(n2895) );
  HS65_LHS_XNOR2X3 U2658 ( .A(a[16]), .B(a[15]), .Z(n2930) );
  HS65_LH_NOR2AX3 U2659 ( .A(n2925), .B(n2926), .Z(n2891) );
  HS65_LHS_XNOR2X3 U2660 ( .A(n2644), .B(a[16]), .Z(n2926) );
  HS65_LHS_XOR2X3 U2661 ( .A(n2640), .B(a[15]), .Z(n2925) );
  HS65_LHS_XOR2X3 U2662 ( .A(n2646), .B(n2932), .Z(n1209) );
  HS65_LH_AO22X4 U2663 ( .A(n2565), .B(n2511), .C(n2564), .D(n2934), .Z(n2932)
         );
  HS65_LHS_XOR2X3 U2664 ( .A(n2646), .B(n2935), .Z(n1208) );
  HS65_LH_AO222X4 U2665 ( .A(n2567), .B(n2511), .C(n2563), .D(n2515), .E(n1038), .F(n2513), .Z(n2935) );
  HS65_LHS_XOR2X3 U2666 ( .A(n2646), .B(n2937), .Z(n1207) );
  HS65_LH_MX41X4 U2667 ( .D0(n2513), .S0(n1037), .D1(n2520), .S1(n2564), .D2(
        n2515), .S2(n2566), .D3(n2511), .S3(n2568), .Z(n2937) );
  HS65_LHS_XOR2X3 U2668 ( .A(n2646), .B(n2939), .Z(n1206) );
  HS65_LH_MX41X4 U2669 ( .D0(n2513), .S0(n1036), .D1(n2519), .S1(n2566), .D2(
        n2515), .S2(n2568), .D3(n2511), .S3(n2570), .Z(n2939) );
  HS65_LHS_XOR2X3 U2670 ( .A(n2646), .B(n2940), .Z(n1205) );
  HS65_LH_MX41X4 U2671 ( .D0(n2513), .S0(n1035), .D1(n2519), .S1(n2568), .D2(
        n2515), .S2(n2570), .D3(n2511), .S3(n2572), .Z(n2940) );
  HS65_LHS_XOR2X3 U2672 ( .A(n2646), .B(n2941), .Z(n1204) );
  HS65_LH_MX41X4 U2673 ( .D0(n2513), .S0(n1034), .D1(n2519), .S1(n2570), .D2(
        n2515), .S2(n2572), .D3(n2511), .S3(n2574), .Z(n2941) );
  HS65_LHS_XOR2X3 U2674 ( .A(n2646), .B(n2942), .Z(n1203) );
  HS65_LH_MX41X4 U2675 ( .D0(n2513), .S0(n1033), .D1(n2519), .S1(n2572), .D2(
        n2515), .S2(n2574), .D3(n2511), .S3(n2576), .Z(n2942) );
  HS65_LHS_XOR2X3 U2676 ( .A(n2646), .B(n2943), .Z(n1202) );
  HS65_LH_MX41X4 U2677 ( .D0(n2513), .S0(n1032), .D1(n2519), .S1(n2574), .D2(
        n2515), .S2(n2576), .D3(n2511), .S3(n2578), .Z(n2943) );
  HS65_LHS_XOR2X3 U2678 ( .A(n2646), .B(n2944), .Z(n1201) );
  HS65_LH_MX41X4 U2679 ( .D0(n2513), .S0(n1031), .D1(n2519), .S1(n2576), .D2(
        n2515), .S2(n2578), .D3(n2511), .S3(n2580), .Z(n2944) );
  HS65_LHS_XOR2X3 U2680 ( .A(n2646), .B(n2945), .Z(n1200) );
  HS65_LH_MX41X4 U2681 ( .D0(n2513), .S0(n1030), .D1(n2519), .S1(n2578), .D2(
        n2516), .S2(n2580), .D3(n2511), .S3(n2582), .Z(n2945) );
  HS65_LHS_XOR2X3 U2682 ( .A(n2646), .B(n2946), .Z(n1199) );
  HS65_LH_MX41X4 U2683 ( .D0(n2513), .S0(n1029), .D1(n2519), .S1(n2580), .D2(
        n2515), .S2(n2582), .D3(n2511), .S3(n2584), .Z(n2946) );
  HS65_LHS_XOR2X3 U2684 ( .A(n2646), .B(n2947), .Z(n1198) );
  HS65_LH_MX41X4 U2685 ( .D0(n2513), .S0(n1028), .D1(n2519), .S1(n2582), .D2(
        n2515), .S2(n2584), .D3(n2511), .S3(n2586), .Z(n2947) );
  HS65_LHS_XOR2X3 U2686 ( .A(n2646), .B(n2948), .Z(n1197) );
  HS65_LH_MX41X4 U2687 ( .D0(n2513), .S0(n1027), .D1(n2519), .S1(n2584), .D2(
        n2515), .S2(n2586), .D3(n2511), .S3(n2589), .Z(n2948) );
  HS65_LHS_XOR2X3 U2688 ( .A(n2646), .B(n2949), .Z(n1196) );
  HS65_LH_MX41X4 U2689 ( .D0(n2513), .S0(n1026), .D1(n2519), .S1(n2586), .D2(
        n2516), .S2(n2588), .D3(n2511), .S3(n2591), .Z(n2949) );
  HS65_LHS_XOR2X3 U2690 ( .A(n2646), .B(n2950), .Z(n1195) );
  HS65_LH_MX41X4 U2691 ( .D0(n2513), .S0(n1025), .D1(n2519), .S1(n2588), .D2(
        n2516), .S2(n2590), .D3(n2511), .S3(n2592), .Z(n2950) );
  HS65_LHS_XOR2X3 U2692 ( .A(n2646), .B(n2951), .Z(n1194) );
  HS65_LH_MX41X4 U2693 ( .D0(n2513), .S0(n1024), .D1(n2520), .S1(n2590), .D2(
        n2516), .S2(n2592), .D3(n2511), .S3(n2594), .Z(n2951) );
  HS65_LHS_XOR2X3 U2694 ( .A(n2646), .B(n2952), .Z(n1193) );
  HS65_LH_MX41X4 U2695 ( .D0(n2513), .S0(n1023), .D1(n2520), .S1(n2592), .D2(
        n2516), .S2(n2594), .D3(n2511), .S3(n2596), .Z(n2952) );
  HS65_LHS_XOR2X3 U2696 ( .A(n2646), .B(n2953), .Z(n1192) );
  HS65_LH_MX41X4 U2697 ( .D0(n2513), .S0(n1022), .D1(n2520), .S1(n2594), .D2(
        n2516), .S2(n2596), .D3(n2512), .S3(n2598), .Z(n2953) );
  HS65_LHS_XOR2X3 U2698 ( .A(n2646), .B(n2954), .Z(n1191) );
  HS65_LH_MX41X4 U2699 ( .D0(n2513), .S0(n1021), .D1(n2520), .S1(n2596), .D2(
        n2516), .S2(n2598), .D3(n2512), .S3(n2601), .Z(n2954) );
  HS65_LHS_XOR2X3 U2700 ( .A(n79), .B(n2955), .Z(n1190) );
  HS65_LH_MX41X4 U2701 ( .D0(n2513), .S0(n1020), .D1(n2520), .S1(n2598), .D2(
        n2516), .S2(n2600), .D3(n2512), .S3(n2603), .Z(n2955) );
  HS65_LHS_XOR2X3 U2702 ( .A(n79), .B(n2956), .Z(n1189) );
  HS65_LH_MX41X4 U2703 ( .D0(n2513), .S0(n1019), .D1(n2520), .S1(n2600), .D2(
        n2516), .S2(n2602), .D3(n2512), .S3(n2605), .Z(n2956) );
  HS65_LHS_XOR2X3 U2704 ( .A(n79), .B(n2957), .Z(n1188) );
  HS65_LH_MX41X4 U2705 ( .D0(n2934), .S0(n1018), .D1(n2520), .S1(n2602), .D2(
        n2516), .S2(n2604), .D3(n2512), .S3(n2606), .Z(n2957) );
  HS65_LHS_XOR2X3 U2706 ( .A(n79), .B(n2958), .Z(n1187) );
  HS65_LH_MX41X4 U2707 ( .D0(n2934), .S0(n1017), .D1(n2520), .S1(n2604), .D2(
        n2516), .S2(n2606), .D3(n2512), .S3(n2608), .Z(n2958) );
  HS65_LHS_XOR2X3 U2708 ( .A(n2647), .B(n2959), .Z(n1186) );
  HS65_LH_MX41X4 U2709 ( .D0(n2934), .S0(n1016), .D1(n2520), .S1(n2606), .D2(
        n2516), .S2(n2608), .D3(n2512), .S3(n2610), .Z(n2959) );
  HS65_LHS_XOR2X3 U2710 ( .A(n2647), .B(n2960), .Z(n1185) );
  HS65_LH_MX41X4 U2711 ( .D0(n2934), .S0(n1015), .D1(n2520), .S1(n2608), .D2(
        n2516), .S2(n2610), .D3(n2512), .S3(n2613), .Z(n2960) );
  HS65_LHS_XOR2X3 U2712 ( .A(n2647), .B(n2961), .Z(n1184) );
  HS65_LH_MX41X4 U2713 ( .D0(n2934), .S0(n1014), .D1(n2520), .S1(n2610), .D2(
        n2516), .S2(n2612), .D3(n2512), .S3(n2615), .Z(n2961) );
  HS65_LHS_XOR2X3 U2714 ( .A(n2647), .B(n2962), .Z(n1183) );
  HS65_LH_MX41X4 U2715 ( .D0(n2934), .S0(n1013), .D1(n2520), .S1(n2612), .D2(
        n2517), .S2(n2614), .D3(n2512), .S3(n2617), .Z(n2962) );
  HS65_LHS_XOR2X3 U2716 ( .A(n2647), .B(n2963), .Z(n1182) );
  HS65_LH_MX41X4 U2717 ( .D0(n2934), .S0(n1012), .D1(n2521), .S1(n2614), .D2(
        n2517), .S2(n2616), .D3(n2512), .S3(n2618), .Z(n2963) );
  HS65_LHS_XOR2X3 U2718 ( .A(n2647), .B(n2964), .Z(n1181) );
  HS65_LH_MX41X4 U2719 ( .D0(n2934), .S0(n1011), .D1(n2521), .S1(n2616), .D2(
        n2517), .S2(n2618), .D3(n2512), .S3(n2620), .Z(n2964) );
  HS65_LHS_XOR2X3 U2720 ( .A(n2647), .B(n2965), .Z(n1180) );
  HS65_LH_MX41X4 U2721 ( .D0(n2934), .S0(n1010), .D1(n2521), .S1(n2618), .D2(
        n2517), .S2(n2620), .D3(n2512), .S3(n2622), .Z(n2965) );
  HS65_LHS_XOR2X3 U2722 ( .A(n2647), .B(n2966), .Z(n1179) );
  HS65_LH_MX41X4 U2723 ( .D0(n2934), .S0(n1009), .D1(n2521), .S1(n2620), .D2(
        n2517), .S2(n2622), .D3(n2512), .S3(n2624), .Z(n2966) );
  HS65_LHS_XOR2X3 U2724 ( .A(n2647), .B(n2967), .Z(n1178) );
  HS65_LH_MX41X4 U2725 ( .D0(n2934), .S0(n1008), .D1(n2521), .S1(n2622), .D2(
        n2515), .S2(n2624), .D3(n2512), .S3(n2626), .Z(n2967) );
  HS65_LH_AND2X4 U2726 ( .A(n2968), .B(n2969), .Z(n2933) );
  HS65_LHS_XOR2X3 U2727 ( .A(n2647), .B(n2970), .Z(n1177) );
  HS65_LH_OAI12X2 U2728 ( .A(n2667), .B(n2514), .C(n2971), .Z(n2970) );
  HS65_LH_OAI22X1 U2729 ( .A(n2625), .B(n2972), .C(n2519), .D(n2972), .Z(n2971) );
  HS65_LH_AND2X4 U2730 ( .A(n2515), .B(n2626), .Z(n2972) );
  HS65_LH_NOR2X2 U2731 ( .A(n2968), .B(n2973), .Z(n2936) );
  HS65_LHS_XOR2X3 U2732 ( .A(n2648), .B(n2974), .Z(n1176) );
  HS65_LH_AOI22X1 U2733 ( .A(n2934), .B(n1006), .C(n2521), .D(n2627), .Z(n2974) );
  HS65_LH_NOR3AX2 U2734 ( .A(n2973), .B(n2969), .C(n2968), .Z(n2938) );
  HS65_LHS_XNOR2X3 U2735 ( .A(a[19]), .B(a[18]), .Z(n2973) );
  HS65_LH_NOR2AX3 U2736 ( .A(n2968), .B(n2969), .Z(n2934) );
  HS65_LHS_XNOR2X3 U2737 ( .A(n2647), .B(a[19]), .Z(n2969) );
  HS65_LHS_XOR2X3 U2738 ( .A(n2643), .B(a[18]), .Z(n2968) );
  HS65_LHS_XOR2X3 U2739 ( .A(n2649), .B(n2975), .Z(n1174) );
  HS65_LH_AO22X4 U2740 ( .A(n2565), .B(n2524), .C(n2564), .D(n2977), .Z(n2975)
         );
  HS65_LHS_XOR2X3 U2741 ( .A(n2649), .B(n2978), .Z(n1173) );
  HS65_LH_AO222X4 U2742 ( .A(n2567), .B(n2524), .C(n2563), .D(n2528), .E(n1038), .F(n2526), .Z(n2978) );
  HS65_LHS_XOR2X3 U2743 ( .A(n2649), .B(n2980), .Z(n1172) );
  HS65_LH_MX41X4 U2744 ( .D0(n2526), .S0(n1037), .D1(n2524), .S1(n2568), .D2(
        n2533), .S2(n2563), .D3(n2528), .S3(n2566), .Z(n2980) );
  HS65_LHS_XOR2X3 U2745 ( .A(n2649), .B(n2982), .Z(n1171) );
  HS65_LH_MX41X4 U2746 ( .D0(n2526), .S0(n1036), .D1(n2524), .S1(n2570), .D2(
        n2532), .S2(n2566), .D3(n2528), .S3(n2568), .Z(n2982) );
  HS65_LHS_XOR2X3 U2747 ( .A(n2649), .B(n2983), .Z(n1170) );
  HS65_LH_MX41X4 U2748 ( .D0(n2526), .S0(n1035), .D1(n2524), .S1(n2572), .D2(
        n2532), .S2(n2568), .D3(n2528), .S3(n2570), .Z(n2983) );
  HS65_LHS_XOR2X3 U2749 ( .A(n2649), .B(n2984), .Z(n1169) );
  HS65_LH_MX41X4 U2750 ( .D0(n2526), .S0(n1034), .D1(n2524), .S1(n2574), .D2(
        n2532), .S2(n2570), .D3(n2528), .S3(n2572), .Z(n2984) );
  HS65_LHS_XOR2X3 U2751 ( .A(n2649), .B(n2985), .Z(n1168) );
  HS65_LH_MX41X4 U2752 ( .D0(n2526), .S0(n1033), .D1(n2524), .S1(n2576), .D2(
        n2532), .S2(n2572), .D3(n2528), .S3(n2574), .Z(n2985) );
  HS65_LHS_XOR2X3 U2753 ( .A(n2649), .B(n2986), .Z(n1167) );
  HS65_LH_MX41X4 U2754 ( .D0(n2526), .S0(n1032), .D1(n2524), .S1(n2578), .D2(
        n2532), .S2(n2574), .D3(n2528), .S3(n2576), .Z(n2986) );
  HS65_LHS_XOR2X3 U2755 ( .A(n2649), .B(n2987), .Z(n1166) );
  HS65_LH_MX41X4 U2756 ( .D0(n2526), .S0(n1031), .D1(n2524), .S1(n2580), .D2(
        n2532), .S2(n2576), .D3(n2528), .S3(n2578), .Z(n2987) );
  HS65_LHS_XOR2X3 U2757 ( .A(n2649), .B(n2988), .Z(n1165) );
  HS65_LH_MX41X4 U2758 ( .D0(n2526), .S0(n1030), .D1(n2524), .S1(n2582), .D2(
        n2532), .S2(n2578), .D3(n2529), .S3(n2580), .Z(n2988) );
  HS65_LHS_XOR2X3 U2759 ( .A(n2649), .B(n2989), .Z(n1164) );
  HS65_LH_MX41X4 U2760 ( .D0(n2526), .S0(n1029), .D1(n2524), .S1(n2584), .D2(
        n2532), .S2(n2580), .D3(n2528), .S3(n2582), .Z(n2989) );
  HS65_LHS_XOR2X3 U2761 ( .A(n2649), .B(n2990), .Z(n1163) );
  HS65_LH_MX41X4 U2762 ( .D0(n2526), .S0(n1028), .D1(n2524), .S1(n2586), .D2(
        n2532), .S2(n2582), .D3(n2528), .S3(n2584), .Z(n2990) );
  HS65_LHS_XOR2X3 U2763 ( .A(n2649), .B(n2991), .Z(n1162) );
  HS65_LH_MX41X4 U2764 ( .D0(n2526), .S0(n1027), .D1(n2524), .S1(n2588), .D2(
        n2532), .S2(n2584), .D3(n2528), .S3(n2586), .Z(n2991) );
  HS65_LHS_XOR2X3 U2765 ( .A(n2649), .B(n2992), .Z(n1161) );
  HS65_LH_MX41X4 U2766 ( .D0(n2526), .S0(n1026), .D1(n2524), .S1(n2590), .D2(
        n2532), .S2(n2586), .D3(n2529), .S3(n2588), .Z(n2992) );
  HS65_LHS_XOR2X3 U2767 ( .A(n2649), .B(n2993), .Z(n1160) );
  HS65_LH_MX41X4 U2768 ( .D0(n2526), .S0(n1025), .D1(n2524), .S1(n2592), .D2(
        n2532), .S2(n2588), .D3(n2529), .S3(n2590), .Z(n2993) );
  HS65_LHS_XOR2X3 U2769 ( .A(n2649), .B(n2994), .Z(n1159) );
  HS65_LH_MX41X4 U2770 ( .D0(n2526), .S0(n1024), .D1(n2524), .S1(n2594), .D2(
        n2533), .S2(n2590), .D3(n2529), .S3(n2592), .Z(n2994) );
  HS65_LHS_XOR2X3 U2771 ( .A(n2649), .B(n2995), .Z(n1158) );
  HS65_LH_MX41X4 U2772 ( .D0(n2526), .S0(n1023), .D1(n2525), .S1(n2596), .D2(
        n2533), .S2(n2592), .D3(n2529), .S3(n2594), .Z(n2995) );
  HS65_LHS_XOR2X3 U2773 ( .A(n2649), .B(n2996), .Z(n1157) );
  HS65_LH_MX41X4 U2774 ( .D0(n2526), .S0(n1022), .D1(n2525), .S1(n2598), .D2(
        n2533), .S2(n2594), .D3(n2529), .S3(n2596), .Z(n2996) );
  HS65_LHS_XOR2X3 U2775 ( .A(n2649), .B(n2997), .Z(n1156) );
  HS65_LH_MX41X4 U2776 ( .D0(n2526), .S0(n1021), .D1(n2525), .S1(n2600), .D2(
        n2533), .S2(n2596), .D3(n2529), .S3(n2598), .Z(n2997) );
  HS65_LHS_XOR2X3 U2777 ( .A(n91), .B(n2998), .Z(n1155) );
  HS65_LH_MX41X4 U2778 ( .D0(n2526), .S0(n1020), .D1(n2525), .S1(n2602), .D2(
        n2533), .S2(n2598), .D3(n2529), .S3(n2600), .Z(n2998) );
  HS65_LHS_XOR2X3 U2779 ( .A(n91), .B(n2999), .Z(n1154) );
  HS65_LH_MX41X4 U2780 ( .D0(n2526), .S0(n1019), .D1(n2525), .S1(n2604), .D2(
        n2533), .S2(n2600), .D3(n2529), .S3(n2602), .Z(n2999) );
  HS65_LHS_XOR2X3 U2781 ( .A(n91), .B(n3000), .Z(n1153) );
  HS65_LH_MX41X4 U2782 ( .D0(n2977), .S0(n1018), .D1(n2525), .S1(n2606), .D2(
        n2533), .S2(n2602), .D3(n2529), .S3(n2604), .Z(n3000) );
  HS65_LHS_XOR2X3 U2783 ( .A(n91), .B(n3001), .Z(n1152) );
  HS65_LH_MX41X4 U2784 ( .D0(n2977), .S0(n1017), .D1(n2525), .S1(n2608), .D2(
        n2533), .S2(n2604), .D3(n2529), .S3(n2606), .Z(n3001) );
  HS65_LHS_XOR2X3 U2785 ( .A(n2650), .B(n3002), .Z(n1151) );
  HS65_LH_MX41X4 U2786 ( .D0(n2977), .S0(n1016), .D1(n2525), .S1(n2610), .D2(
        n2533), .S2(n2606), .D3(n2529), .S3(n2608), .Z(n3002) );
  HS65_LHS_XOR2X3 U2787 ( .A(n2650), .B(n3003), .Z(n1150) );
  HS65_LH_MX41X4 U2788 ( .D0(n2977), .S0(n1015), .D1(n2525), .S1(n2612), .D2(
        n2533), .S2(n2608), .D3(n2529), .S3(n2610), .Z(n3003) );
  HS65_LHS_XOR2X3 U2789 ( .A(n2650), .B(n3004), .Z(n1149) );
  HS65_LH_MX41X4 U2790 ( .D0(n2977), .S0(n1014), .D1(n2525), .S1(n2614), .D2(
        n2533), .S2(n2610), .D3(n2529), .S3(n2612), .Z(n3004) );
  HS65_LHS_XOR2X3 U2791 ( .A(n2650), .B(n3005), .Z(n1148) );
  HS65_LH_MX41X4 U2792 ( .D0(n2977), .S0(n1013), .D1(n2525), .S1(n2616), .D2(
        n2533), .S2(n2612), .D3(n2530), .S3(n2614), .Z(n3005) );
  HS65_LHS_XOR2X3 U2793 ( .A(n2650), .B(n3006), .Z(n1147) );
  HS65_LH_MX41X4 U2794 ( .D0(n2977), .S0(n1012), .D1(n2525), .S1(n2618), .D2(
        n2533), .S2(n2614), .D3(n2530), .S3(n2616), .Z(n3006) );
  HS65_LHS_XOR2X3 U2795 ( .A(n2650), .B(n3007), .Z(n1146) );
  HS65_LH_MX41X4 U2796 ( .D0(n2977), .S0(n1011), .D1(n2525), .S1(n2620), .D2(
        n2534), .S2(n2616), .D3(n2530), .S3(n2618), .Z(n3007) );
  HS65_LHS_XOR2X3 U2797 ( .A(n2650), .B(n3008), .Z(n1145) );
  HS65_LH_MX41X4 U2798 ( .D0(n2977), .S0(n1010), .D1(n2525), .S1(n2622), .D2(
        n2534), .S2(n2618), .D3(n2530), .S3(n2620), .Z(n3008) );
  HS65_LHS_XOR2X3 U2799 ( .A(n2650), .B(n3009), .Z(n1144) );
  HS65_LH_MX41X4 U2800 ( .D0(n2977), .S0(n1009), .D1(n2525), .S1(n2624), .D2(
        n2534), .S2(n2620), .D3(n2530), .S3(n2622), .Z(n3009) );
  HS65_LHS_XOR2X3 U2801 ( .A(n2650), .B(n3010), .Z(n1143) );
  HS65_LH_MX41X4 U2802 ( .D0(n2977), .S0(n1008), .D1(n2525), .S1(n2626), .D2(
        n2534), .S2(n2622), .D3(n2528), .S3(n2624), .Z(n3010) );
  HS65_LH_AND2X4 U2803 ( .A(n3011), .B(n3012), .Z(n2976) );
  HS65_LHS_XOR2X3 U2804 ( .A(n2650), .B(n3013), .Z(n1142) );
  HS65_LH_OAI12X2 U2805 ( .A(n2667), .B(n2527), .C(n3014), .Z(n3013) );
  HS65_LH_OAI22X1 U2806 ( .A(n2625), .B(n3015), .C(n2532), .D(n3015), .Z(n3014) );
  HS65_LH_AND2X4 U2807 ( .A(n2528), .B(n2626), .Z(n3015) );
  HS65_LH_NOR2X2 U2808 ( .A(n3011), .B(n3016), .Z(n2979) );
  HS65_LHS_XOR2X3 U2809 ( .A(n2651), .B(n3017), .Z(n1141) );
  HS65_LH_AOI22X1 U2810 ( .A(n2977), .B(n1006), .C(n2534), .D(n2627), .Z(n3017) );
  HS65_LH_NOR3AX2 U2811 ( .A(n3016), .B(n3012), .C(n3011), .Z(n2981) );
  HS65_LHS_XNOR2X3 U2812 ( .A(a[22]), .B(a[21]), .Z(n3016) );
  HS65_LH_NOR2AX3 U2813 ( .A(n3011), .B(n3012), .Z(n2977) );
  HS65_LHS_XNOR2X3 U2814 ( .A(n2650), .B(a[22]), .Z(n3012) );
  HS65_LHS_XOR2X3 U2815 ( .A(n2646), .B(a[21]), .Z(n3011) );
  HS65_LHS_XOR2X3 U2816 ( .A(n2652), .B(n3018), .Z(n1139) );
  HS65_LH_AO22X4 U2817 ( .A(n2565), .B(n2537), .C(n2564), .D(n3020), .Z(n3018)
         );
  HS65_LHS_XOR2X3 U2818 ( .A(n2652), .B(n3021), .Z(n1138) );
  HS65_LH_AO222X4 U2819 ( .A(n2567), .B(n2537), .C(n2563), .D(n2541), .E(n1038), .F(n2539), .Z(n3021) );
  HS65_LHS_XOR2X3 U2820 ( .A(n2652), .B(n3023), .Z(n1137) );
  HS65_LH_MX41X4 U2821 ( .D0(n2539), .S0(n1037), .D1(n2546), .S1(n2563), .D2(
        n2541), .S2(n2566), .D3(n2537), .S3(n2568), .Z(n3023) );
  HS65_LHS_XOR2X3 U2822 ( .A(n2652), .B(n3025), .Z(n1136) );
  HS65_LH_MX41X4 U2823 ( .D0(n2539), .S0(n1036), .D1(n2545), .S1(n2567), .D2(
        n2541), .S2(n2568), .D3(n2537), .S3(n2570), .Z(n3025) );
  HS65_LHS_XOR2X3 U2824 ( .A(n2652), .B(n3026), .Z(n1135) );
  HS65_LH_MX41X4 U2825 ( .D0(n2539), .S0(n1035), .D1(n2545), .S1(n2568), .D2(
        n2541), .S2(n2570), .D3(n2537), .S3(n2572), .Z(n3026) );
  HS65_LHS_XOR2X3 U2826 ( .A(n2652), .B(n3027), .Z(n1134) );
  HS65_LH_MX41X4 U2827 ( .D0(n2539), .S0(n1034), .D1(n2545), .S1(n2570), .D2(
        n2541), .S2(n2572), .D3(n2537), .S3(n2574), .Z(n3027) );
  HS65_LHS_XOR2X3 U2828 ( .A(n2652), .B(n3028), .Z(n1133) );
  HS65_LH_MX41X4 U2829 ( .D0(n2539), .S0(n1033), .D1(n2545), .S1(n2572), .D2(
        n2541), .S2(n2574), .D3(n2537), .S3(n2576), .Z(n3028) );
  HS65_LHS_XOR2X3 U2830 ( .A(n2652), .B(n3029), .Z(n1132) );
  HS65_LH_MX41X4 U2831 ( .D0(n2539), .S0(n1032), .D1(n2545), .S1(n2574), .D2(
        n2541), .S2(n2576), .D3(n2537), .S3(n2578), .Z(n3029) );
  HS65_LHS_XOR2X3 U2832 ( .A(n2652), .B(n3030), .Z(n1131) );
  HS65_LH_MX41X4 U2833 ( .D0(n2539), .S0(n1031), .D1(n2545), .S1(n2576), .D2(
        n2541), .S2(n2578), .D3(n2537), .S3(n2580), .Z(n3030) );
  HS65_LHS_XOR2X3 U2834 ( .A(n2652), .B(n3031), .Z(n1130) );
  HS65_LH_MX41X4 U2835 ( .D0(n2539), .S0(n1030), .D1(n2545), .S1(n2578), .D2(
        n2542), .S2(n2580), .D3(n2537), .S3(n2582), .Z(n3031) );
  HS65_LHS_XOR2X3 U2836 ( .A(n2652), .B(n3032), .Z(n1129) );
  HS65_LH_MX41X4 U2837 ( .D0(n2539), .S0(n1029), .D1(n2545), .S1(n2580), .D2(
        n2541), .S2(n2582), .D3(n2537), .S3(n2584), .Z(n3032) );
  HS65_LHS_XOR2X3 U2838 ( .A(n2652), .B(n3033), .Z(n1128) );
  HS65_LH_MX41X4 U2839 ( .D0(n2539), .S0(n1028), .D1(n2545), .S1(n2582), .D2(
        n2541), .S2(n2584), .D3(n2537), .S3(n2586), .Z(n3033) );
  HS65_LHS_XOR2X3 U2840 ( .A(n2652), .B(n3034), .Z(n1127) );
  HS65_LH_MX41X4 U2841 ( .D0(n2539), .S0(n1027), .D1(n2545), .S1(n2584), .D2(
        n2541), .S2(n2586), .D3(n2537), .S3(n2588), .Z(n3034) );
  HS65_LHS_XOR2X3 U2842 ( .A(n2652), .B(n3035), .Z(n1126) );
  HS65_LH_MX41X4 U2843 ( .D0(n2539), .S0(n1026), .D1(n2545), .S1(n2586), .D2(
        n2542), .S2(n2588), .D3(n2537), .S3(n2590), .Z(n3035) );
  HS65_LHS_XOR2X3 U2844 ( .A(n2652), .B(n3036), .Z(n1125) );
  HS65_LH_MX41X4 U2845 ( .D0(n2539), .S0(n1025), .D1(n2545), .S1(n2588), .D2(
        n2542), .S2(n2590), .D3(n2537), .S3(n2592), .Z(n3036) );
  HS65_LHS_XOR2X3 U2846 ( .A(n2652), .B(n3037), .Z(n1124) );
  HS65_LH_MX41X4 U2847 ( .D0(n2539), .S0(n1024), .D1(n2546), .S1(n2590), .D2(
        n2542), .S2(n2592), .D3(n2537), .S3(n2594), .Z(n3037) );
  HS65_LHS_XOR2X3 U2848 ( .A(n2652), .B(n3038), .Z(n1123) );
  HS65_LH_MX41X4 U2849 ( .D0(n2539), .S0(n1023), .D1(n2546), .S1(n2592), .D2(
        n2542), .S2(n2594), .D3(n2537), .S3(n2596), .Z(n3038) );
  HS65_LHS_XOR2X3 U2850 ( .A(n2652), .B(n3039), .Z(n1122) );
  HS65_LH_MX41X4 U2851 ( .D0(n2539), .S0(n1022), .D1(n2546), .S1(n2594), .D2(
        n2542), .S2(n2596), .D3(n2538), .S3(n2598), .Z(n3039) );
  HS65_LHS_XOR2X3 U2852 ( .A(n2652), .B(n3040), .Z(n1121) );
  HS65_LH_MX41X4 U2853 ( .D0(n2539), .S0(n1021), .D1(n2546), .S1(n2596), .D2(
        n2542), .S2(n2598), .D3(n2538), .S3(n2600), .Z(n3040) );
  HS65_LHS_XOR2X3 U2854 ( .A(n103), .B(n3041), .Z(n1120) );
  HS65_LH_MX41X4 U2855 ( .D0(n2539), .S0(n1020), .D1(n2546), .S1(n2598), .D2(
        n2542), .S2(n2600), .D3(n2538), .S3(n2602), .Z(n3041) );
  HS65_LHS_XOR2X3 U2856 ( .A(n103), .B(n3042), .Z(n1119) );
  HS65_LH_MX41X4 U2857 ( .D0(n2539), .S0(n1019), .D1(n2546), .S1(n2600), .D2(
        n2542), .S2(n2602), .D3(n2538), .S3(n2604), .Z(n3042) );
  HS65_LHS_XOR2X3 U2858 ( .A(n103), .B(n3043), .Z(n1118) );
  HS65_LH_MX41X4 U2859 ( .D0(n3020), .S0(n1018), .D1(n2546), .S1(n2602), .D2(
        n2542), .S2(n2604), .D3(n2538), .S3(n2606), .Z(n3043) );
  HS65_LHS_XOR2X3 U2860 ( .A(n103), .B(n3044), .Z(n1117) );
  HS65_LH_MX41X4 U2861 ( .D0(n3020), .S0(n1017), .D1(n2546), .S1(n2604), .D2(
        n2542), .S2(n2606), .D3(n2538), .S3(n2608), .Z(n3044) );
  HS65_LHS_XOR2X3 U2862 ( .A(n2653), .B(n3045), .Z(n1116) );
  HS65_LH_MX41X4 U2863 ( .D0(n3020), .S0(n1016), .D1(n2546), .S1(n2606), .D2(
        n2542), .S2(n2608), .D3(n2538), .S3(n2610), .Z(n3045) );
  HS65_LHS_XOR2X3 U2864 ( .A(n2653), .B(n3046), .Z(n1115) );
  HS65_LH_MX41X4 U2865 ( .D0(n3020), .S0(n1015), .D1(n2546), .S1(n2608), .D2(
        n2542), .S2(n2610), .D3(n2538), .S3(n2612), .Z(n3046) );
  HS65_LHS_XOR2X3 U2866 ( .A(n2653), .B(n3047), .Z(n1114) );
  HS65_LH_MX41X4 U2867 ( .D0(n3020), .S0(n1014), .D1(n2546), .S1(n2610), .D2(
        n2542), .S2(n2612), .D3(n2538), .S3(n2614), .Z(n3047) );
  HS65_LHS_XOR2X3 U2868 ( .A(n2653), .B(n3048), .Z(n1113) );
  HS65_LH_MX41X4 U2869 ( .D0(n3020), .S0(n1013), .D1(n2546), .S1(n2612), .D2(
        n2543), .S2(n2614), .D3(n2538), .S3(n2616), .Z(n3048) );
  HS65_LHS_XOR2X3 U2870 ( .A(n2653), .B(n3049), .Z(n1112) );
  HS65_LH_MX41X4 U2871 ( .D0(n3020), .S0(n1012), .D1(n2547), .S1(n2614), .D2(
        n2543), .S2(n2616), .D3(n2538), .S3(n2618), .Z(n3049) );
  HS65_LHS_XOR2X3 U2872 ( .A(n2653), .B(n3050), .Z(n1111) );
  HS65_LH_MX41X4 U2873 ( .D0(n3020), .S0(n1011), .D1(n2547), .S1(n2616), .D2(
        n2543), .S2(n2618), .D3(n2538), .S3(n2620), .Z(n3050) );
  HS65_LHS_XOR2X3 U2874 ( .A(n2653), .B(n3051), .Z(n1110) );
  HS65_LH_MX41X4 U2875 ( .D0(n3020), .S0(n1010), .D1(n2547), .S1(n2618), .D2(
        n2543), .S2(n2620), .D3(n2538), .S3(n2622), .Z(n3051) );
  HS65_LHS_XOR2X3 U2876 ( .A(n2653), .B(n3052), .Z(n1109) );
  HS65_LH_MX41X4 U2877 ( .D0(n3020), .S0(n1009), .D1(n2547), .S1(n2620), .D2(
        n2543), .S2(n2622), .D3(n2538), .S3(n2624), .Z(n3052) );
  HS65_LHS_XOR2X3 U2878 ( .A(n2653), .B(n3053), .Z(n1108) );
  HS65_LH_MX41X4 U2879 ( .D0(n3020), .S0(n1008), .D1(n2547), .S1(n2622), .D2(
        n2541), .S2(n2624), .D3(n2538), .S3(n2626), .Z(n3053) );
  HS65_LH_AND2X4 U2880 ( .A(n3054), .B(n3055), .Z(n3019) );
  HS65_LHS_XOR2X3 U2881 ( .A(n2653), .B(n3056), .Z(n1107) );
  HS65_LH_OAI12X2 U2882 ( .A(n2667), .B(n2540), .C(n3057), .Z(n3056) );
  HS65_LH_OAI22X1 U2883 ( .A(n2625), .B(n3058), .C(n2545), .D(n3058), .Z(n3057) );
  HS65_LH_AND2X4 U2884 ( .A(n2541), .B(n2626), .Z(n3058) );
  HS65_LH_NOR2X2 U2885 ( .A(n3054), .B(n3059), .Z(n3022) );
  HS65_LHS_XOR2X3 U2886 ( .A(n2654), .B(n3060), .Z(n1106) );
  HS65_LH_AOI22X1 U2887 ( .A(n3020), .B(n1006), .C(n2547), .D(n2627), .Z(n3060) );
  HS65_LH_NOR3AX2 U2888 ( .A(n3059), .B(n3055), .C(n3054), .Z(n3024) );
  HS65_LHS_XNOR2X3 U2889 ( .A(a[25]), .B(a[24]), .Z(n3059) );
  HS65_LH_NOR2AX3 U2890 ( .A(n3054), .B(n3055), .Z(n3020) );
  HS65_LHS_XNOR2X3 U2891 ( .A(n2653), .B(a[25]), .Z(n3055) );
  HS65_LHS_XOR2X3 U2892 ( .A(n2649), .B(a[24]), .Z(n3054) );
  HS65_LHS_XOR2X3 U2893 ( .A(n2655), .B(n3061), .Z(n1104) );
  HS65_LH_AO22X4 U2894 ( .A(n2565), .B(n2550), .C(n2564), .D(n3063), .Z(n3061)
         );
  HS65_LHS_XOR2X3 U2895 ( .A(n2655), .B(n3064), .Z(n1103) );
  HS65_LH_AO222X4 U2896 ( .A(n2567), .B(n2550), .C(n2563), .D(n2554), .E(n1038), .F(n2552), .Z(n3064) );
  HS65_LHS_XOR2X3 U2897 ( .A(n2655), .B(n3066), .Z(n1102) );
  HS65_LH_MX41X4 U2898 ( .D0(n2552), .S0(n1037), .D1(n2559), .S1(n2563), .D2(
        n2554), .S2(n2566), .D3(n2550), .S3(n2568), .Z(n3066) );
  HS65_LHS_XOR2X3 U2899 ( .A(n2655), .B(n3068), .Z(n1101) );
  HS65_LH_MX41X4 U2900 ( .D0(n2552), .S0(n1036), .D1(n2558), .S1(n2567), .D2(
        n2554), .S2(n2568), .D3(n2550), .S3(n2570), .Z(n3068) );
  HS65_LHS_XOR2X3 U2901 ( .A(n2655), .B(n3069), .Z(n1100) );
  HS65_LH_MX41X4 U2902 ( .D0(n2552), .S0(n1035), .D1(n2558), .S1(n2568), .D2(
        n2554), .S2(n2570), .D3(n2550), .S3(n2572), .Z(n3069) );
  HS65_LHS_XOR2X3 U2903 ( .A(n2655), .B(n3070), .Z(n1099) );
  HS65_LH_MX41X4 U2904 ( .D0(n2552), .S0(n1034), .D1(n2558), .S1(n2570), .D2(
        n2554), .S2(n2572), .D3(n2550), .S3(n2574), .Z(n3070) );
  HS65_LHS_XOR2X3 U2905 ( .A(n2655), .B(n3071), .Z(n1098) );
  HS65_LH_MX41X4 U2906 ( .D0(n2552), .S0(n1033), .D1(n2558), .S1(n2572), .D2(
        n2554), .S2(n2574), .D3(n2550), .S3(n2576), .Z(n3071) );
  HS65_LHS_XOR2X3 U2907 ( .A(n2655), .B(n3072), .Z(n1097) );
  HS65_LH_MX41X4 U2908 ( .D0(n2552), .S0(n1032), .D1(n2558), .S1(n2574), .D2(
        n2554), .S2(n2576), .D3(n2550), .S3(n2578), .Z(n3072) );
  HS65_LHS_XOR2X3 U2909 ( .A(n2655), .B(n3073), .Z(n1096) );
  HS65_LH_MX41X4 U2910 ( .D0(n2552), .S0(n1031), .D1(n2558), .S1(n2576), .D2(
        n2554), .S2(n2578), .D3(n2550), .S3(n2580), .Z(n3073) );
  HS65_LHS_XOR2X3 U2911 ( .A(n2655), .B(n3074), .Z(n1095) );
  HS65_LH_MX41X4 U2912 ( .D0(n2552), .S0(n1030), .D1(n2558), .S1(n2578), .D2(
        n2555), .S2(n2580), .D3(n2550), .S3(n2582), .Z(n3074) );
  HS65_LHS_XOR2X3 U2913 ( .A(n2655), .B(n3075), .Z(n1094) );
  HS65_LH_MX41X4 U2914 ( .D0(n2552), .S0(n1029), .D1(n2558), .S1(n2580), .D2(
        n2554), .S2(n2582), .D3(n2550), .S3(n2584), .Z(n3075) );
  HS65_LHS_XOR2X3 U2915 ( .A(n2655), .B(n3076), .Z(n1093) );
  HS65_LH_MX41X4 U2916 ( .D0(n2552), .S0(n1028), .D1(n2558), .S1(n2582), .D2(
        n2554), .S2(n2584), .D3(n2550), .S3(n2586), .Z(n3076) );
  HS65_LHS_XOR2X3 U2917 ( .A(n2655), .B(n3077), .Z(n1092) );
  HS65_LH_MX41X4 U2918 ( .D0(n2552), .S0(n1027), .D1(n2558), .S1(n2584), .D2(
        n2554), .S2(n2586), .D3(n2550), .S3(n2588), .Z(n3077) );
  HS65_LHS_XOR2X3 U2919 ( .A(n2655), .B(n3078), .Z(n1091) );
  HS65_LH_MX41X4 U2920 ( .D0(n2552), .S0(n1026), .D1(n2558), .S1(n2586), .D2(
        n2555), .S2(n2588), .D3(n2550), .S3(n2590), .Z(n3078) );
  HS65_LHS_XOR2X3 U2921 ( .A(n2655), .B(n3079), .Z(n1090) );
  HS65_LH_MX41X4 U2922 ( .D0(n2552), .S0(n1025), .D1(n2558), .S1(n2588), .D2(
        n2555), .S2(n2590), .D3(n2550), .S3(n2592), .Z(n3079) );
  HS65_LHS_XOR2X3 U2923 ( .A(n2655), .B(n3080), .Z(n1089) );
  HS65_LH_MX41X4 U2924 ( .D0(n2552), .S0(n1024), .D1(n2559), .S1(n2590), .D2(
        n2555), .S2(n2592), .D3(n2550), .S3(n2594), .Z(n3080) );
  HS65_LHS_XOR2X3 U2925 ( .A(n2655), .B(n3081), .Z(n1088) );
  HS65_LH_MX41X4 U2926 ( .D0(n2552), .S0(n1023), .D1(n2559), .S1(n2592), .D2(
        n2555), .S2(n2594), .D3(n2550), .S3(n2596), .Z(n3081) );
  HS65_LHS_XOR2X3 U2927 ( .A(n2655), .B(n3082), .Z(n1087) );
  HS65_LH_MX41X4 U2928 ( .D0(n2552), .S0(n1022), .D1(n2559), .S1(n2594), .D2(
        n2555), .S2(n2596), .D3(n2551), .S3(n2598), .Z(n3082) );
  HS65_LHS_XOR2X3 U2929 ( .A(n2655), .B(n3083), .Z(n1086) );
  HS65_LH_MX41X4 U2930 ( .D0(n2552), .S0(n1021), .D1(n2559), .S1(n2596), .D2(
        n2555), .S2(n2598), .D3(n2551), .S3(n2600), .Z(n3083) );
  HS65_LHS_XOR2X3 U2931 ( .A(n115), .B(n3084), .Z(n1085) );
  HS65_LH_MX41X4 U2932 ( .D0(n2552), .S0(n1020), .D1(n2559), .S1(n2598), .D2(
        n2555), .S2(n2600), .D3(n2551), .S3(n2602), .Z(n3084) );
  HS65_LHS_XOR2X3 U2933 ( .A(n115), .B(n3085), .Z(n1084) );
  HS65_LH_MX41X4 U2934 ( .D0(n2552), .S0(n1019), .D1(n2559), .S1(n2600), .D2(
        n2555), .S2(n2602), .D3(n2551), .S3(n2604), .Z(n3085) );
  HS65_LHS_XOR2X3 U2935 ( .A(n115), .B(n3086), .Z(n1083) );
  HS65_LH_MX41X4 U2936 ( .D0(n3063), .S0(n1018), .D1(n2559), .S1(n2602), .D2(
        n2555), .S2(n2604), .D3(n2551), .S3(n2606), .Z(n3086) );
  HS65_LHS_XOR2X3 U2937 ( .A(n115), .B(n3087), .Z(n1082) );
  HS65_LH_MX41X4 U2938 ( .D0(n3063), .S0(n1017), .D1(n2559), .S1(n2604), .D2(
        n2555), .S2(n2606), .D3(n2551), .S3(n2608), .Z(n3087) );
  HS65_LHS_XOR2X3 U2939 ( .A(n2656), .B(n3088), .Z(n1081) );
  HS65_LH_MX41X4 U2940 ( .D0(n3063), .S0(n1016), .D1(n2559), .S1(n2606), .D2(
        n2555), .S2(n2608), .D3(n2551), .S3(n2610), .Z(n3088) );
  HS65_LHS_XOR2X3 U2941 ( .A(n2656), .B(n3089), .Z(n1080) );
  HS65_LH_MX41X4 U2942 ( .D0(n3063), .S0(n1015), .D1(n2559), .S1(n2608), .D2(
        n2555), .S2(n2610), .D3(n2551), .S3(n2612), .Z(n3089) );
  HS65_LHS_XOR2X3 U2943 ( .A(n2656), .B(n3090), .Z(n1079) );
  HS65_LH_MX41X4 U2944 ( .D0(n3063), .S0(n1014), .D1(n2559), .S1(n2610), .D2(
        n2555), .S2(n2612), .D3(n2551), .S3(n2614), .Z(n3090) );
  HS65_LHS_XOR2X3 U2945 ( .A(n2656), .B(n3091), .Z(n1078) );
  HS65_LH_MX41X4 U2946 ( .D0(n3063), .S0(n1013), .D1(n2559), .S1(n2612), .D2(
        n2556), .S2(n2614), .D3(n2551), .S3(n2616), .Z(n3091) );
  HS65_LHS_XOR2X3 U2947 ( .A(n2656), .B(n3092), .Z(n1077) );
  HS65_LH_MX41X4 U2948 ( .D0(n3063), .S0(n1012), .D1(n2560), .S1(n2614), .D2(
        n2556), .S2(n2616), .D3(n2551), .S3(n2618), .Z(n3092) );
  HS65_LHS_XOR2X3 U2949 ( .A(n2656), .B(n3093), .Z(n1076) );
  HS65_LH_MX41X4 U2950 ( .D0(n3063), .S0(n1011), .D1(n2560), .S1(n2616), .D2(
        n2556), .S2(n2618), .D3(n2551), .S3(n2620), .Z(n3093) );
  HS65_LHS_XOR2X3 U2951 ( .A(n2656), .B(n3094), .Z(n1075) );
  HS65_LH_MX41X4 U2952 ( .D0(n3063), .S0(n1010), .D1(n2560), .S1(n2618), .D2(
        n2556), .S2(n2620), .D3(n2551), .S3(n2622), .Z(n3094) );
  HS65_LHS_XOR2X3 U2953 ( .A(n2656), .B(n3095), .Z(n1074) );
  HS65_LH_MX41X4 U2954 ( .D0(n3063), .S0(n1009), .D1(n2560), .S1(n2620), .D2(
        n2556), .S2(n2622), .D3(n2551), .S3(n2624), .Z(n3095) );
  HS65_LHS_XOR2X3 U2955 ( .A(n2656), .B(n3096), .Z(n1073) );
  HS65_LH_MX41X4 U2956 ( .D0(n3063), .S0(n1008), .D1(n2560), .S1(n2622), .D2(
        n2554), .S2(n2624), .D3(n2551), .S3(n2626), .Z(n3096) );
  HS65_LH_AND2X4 U2957 ( .A(n3097), .B(n3098), .Z(n3062) );
  HS65_LHS_XOR2X3 U2958 ( .A(n2656), .B(n3099), .Z(n1072) );
  HS65_LH_OAI12X2 U2959 ( .A(n2667), .B(n2553), .C(n3100), .Z(n3099) );
  HS65_LH_OAI22X1 U2960 ( .A(n2625), .B(n3101), .C(n2558), .D(n3101), .Z(n3100) );
  HS65_LH_AND2X4 U2961 ( .A(n2554), .B(n2626), .Z(n3101) );
  HS65_LH_NOR2X2 U2962 ( .A(n3097), .B(n3102), .Z(n3065) );
  HS65_LHS_XOR2X3 U2963 ( .A(n2657), .B(n3103), .Z(n1071) );
  HS65_LH_AOI22X1 U2964 ( .A(n3063), .B(n1006), .C(n2560), .D(n2627), .Z(n3103) );
  HS65_LH_NOR3AX2 U2965 ( .A(n3102), .B(n3098), .C(n3097), .Z(n3067) );
  HS65_LHS_XNOR2X3 U2966 ( .A(a[28]), .B(a[27]), .Z(n3102) );
  HS65_LH_NOR2AX3 U2967 ( .A(n3097), .B(n3098), .Z(n3063) );
  HS65_LHS_XNOR2X3 U2968 ( .A(n2656), .B(a[28]), .Z(n3098) );
  HS65_LHS_XOR2X3 U2969 ( .A(n2652), .B(a[27]), .Z(n3097) );
  HS65_LH_AO22X4 U2970 ( .A(n2428), .B(n2563), .C(n2419), .D(n2564), .Z(n1069)
         );
  HS65_LH_AO222X4 U2971 ( .A(n2428), .B(n2566), .C(n2432), .D(n2563), .E(n2419), .F(n1038), .Z(n1068) );
  HS65_LH_MX41X4 U2972 ( .D0(n1037), .S0(n2419), .D1(n2569), .S1(n2426), .D2(
        n2567), .S2(n2430), .D3(n2564), .S3(n2423), .Z(n1067) );
  HS65_LH_MX41X4 U2973 ( .D0(n1036), .S0(n2419), .D1(n2571), .S1(n2426), .D2(
        n2569), .S2(n2430), .D3(n2567), .S3(n2423), .Z(n1066) );
  HS65_LH_MX41X4 U2974 ( .D0(n1035), .S0(n2419), .D1(n2573), .S1(n2426), .D2(
        n2571), .S2(n2430), .D3(n2569), .S3(n2423), .Z(n1065) );
  HS65_LH_MX41X4 U2975 ( .D0(n1034), .S0(n2418), .D1(n2575), .S1(n2426), .D2(
        n2573), .S2(n2430), .D3(n2571), .S3(n2423), .Z(n1064) );
  HS65_LH_MX41X4 U2976 ( .D0(n1033), .S0(n2418), .D1(n2577), .S1(n2426), .D2(
        n2575), .S2(n2430), .D3(n2573), .S3(n2423), .Z(n1063) );
  HS65_LH_MX41X4 U2977 ( .D0(n1032), .S0(n2418), .D1(n2579), .S1(n2426), .D2(
        n2577), .S2(n2430), .D3(n2575), .S3(n2423), .Z(n1062) );
  HS65_LH_MX41X4 U2978 ( .D0(n1031), .S0(n2418), .D1(n2581), .S1(n2426), .D2(
        n2579), .S2(n2430), .D3(n2577), .S3(n2423), .Z(n1061) );
  HS65_LH_MX41X4 U2979 ( .D0(n1030), .S0(n2418), .D1(n2583), .S1(n2426), .D2(
        n2581), .S2(n2430), .D3(n2579), .S3(n2423), .Z(n1060) );
  HS65_LH_MX41X4 U2980 ( .D0(n1029), .S0(n2418), .D1(n2585), .S1(n2426), .D2(
        n2583), .S2(n2430), .D3(n2581), .S3(n2423), .Z(n1059) );
  HS65_LH_MX41X4 U2981 ( .D0(n1028), .S0(n2418), .D1(n2587), .S1(n2426), .D2(
        n2585), .S2(n2431), .D3(n2583), .S3(n2424), .Z(n1058) );
  HS65_LH_MX41X4 U2982 ( .D0(n1027), .S0(n2418), .D1(n2428), .S1(n2588), .D2(
        n2587), .S2(n2431), .D3(n2585), .S3(n2424), .Z(n1057) );
  HS65_LH_MX41X4 U2983 ( .D0(n1026), .S0(n2418), .D1(n2428), .S1(n2590), .D2(
        n2589), .S2(n2431), .D3(n2587), .S3(n2424), .Z(n1056) );
  HS65_LH_MX41X4 U2984 ( .D0(n1024), .S0(n2418), .D1(n2593), .S1(n2432), .D2(
        n2591), .S2(n2423), .D3(n2595), .S3(n2426), .Z(n1055) );
  HS65_LH_MX41X4 U2985 ( .D0(n1023), .S0(n2418), .D1(n2593), .S1(n2424), .D2(
        n2595), .S2(n2431), .D3(n2597), .S3(n2427), .Z(n1054) );
  HS65_LH_MX41X4 U2986 ( .D0(n1022), .S0(n2417), .D1(n2595), .S1(n2424), .D2(
        n2597), .S2(n2431), .D3(n2599), .S3(n2427), .Z(n1053) );
  HS65_LH_MX41X4 U2987 ( .D0(n1021), .S0(n2417), .D1(n2597), .S1(n2424), .D2(
        n2599), .S2(n2431), .D3(n2601), .S3(n2427), .Z(n1052) );
  HS65_LH_MX41X4 U2988 ( .D0(n1020), .S0(n2417), .D1(n2599), .S1(n2424), .D2(
        n2601), .S2(n2431), .D3(n2603), .S3(n2427), .Z(n1051) );
  HS65_LH_MX41X4 U2989 ( .D0(n1018), .S0(n2417), .D1(n2603), .S1(n2424), .D2(
        n2605), .S2(n2431), .D3(n2607), .S3(n2427), .Z(n1050) );
  HS65_LH_MX41X4 U2990 ( .D0(n1017), .S0(n2417), .D1(n2605), .S1(n2424), .D2(
        n2607), .S2(n2431), .D3(n2609), .S3(n2427), .Z(n1049) );
  HS65_LH_MX41X4 U2991 ( .D0(n1016), .S0(n2417), .D1(n2607), .S1(n2424), .D2(
        n2609), .S2(n2431), .D3(n2611), .S3(n2427), .Z(n1048) );
  HS65_LH_MX41X4 U2992 ( .D0(n1015), .S0(n2417), .D1(n2609), .S1(n2424), .D2(
        n2611), .S2(n2431), .D3(n2613), .S3(n2427), .Z(n1047) );
  HS65_LH_MX41X4 U2993 ( .D0(n1014), .S0(n2417), .D1(n2611), .S1(n2424), .D2(
        n2613), .S2(n2432), .D3(n2615), .S3(n2427), .Z(n1046) );
  HS65_LH_MX41X4 U2994 ( .D0(n1012), .S0(n2417), .D1(n2615), .S1(n2424), .D2(
        n2617), .S2(n2432), .D3(n2619), .S3(n2427), .Z(n1045) );
  HS65_LH_MX41X4 U2995 ( .D0(n1011), .S0(n2417), .D1(n2617), .S1(n2424), .D2(
        n2619), .S2(n2432), .D3(n2621), .S3(n2427), .Z(n1044) );
  HS65_LH_MX41X4 U2996 ( .D0(n1010), .S0(n2417), .D1(n2619), .S1(n2424), .D2(
        n2621), .S2(n2432), .D3(n2623), .S3(n2427), .Z(n1043) );
  HS65_LH_MX41X4 U2997 ( .D0(n1009), .S0(n2417), .D1(n2621), .S1(n2423), .D2(
        n2623), .S2(n2431), .D3(n2625), .S3(n2428), .Z(n1042) );
  HS65_LH_MX41X4 U2998 ( .D0(n1008), .S0(n2418), .D1(n2623), .S1(n2424), .D2(
        n2625), .S2(n2430), .D3(n2428), .S3(n2626), .Z(n1041) );
  HS65_LH_NOR2AX3 U2999 ( .A(n3104), .B(a[31]), .Z(n2671) );
  HS65_LH_NOR2AX3 U3000 ( .A(n3105), .B(n3104), .Z(n2672) );
  HS65_LH_NOR3AX2 U3001 ( .A(a[31]), .B(n3105), .C(n3104), .Z(n2670) );
  HS65_LHS_XOR2X3 U3002 ( .A(a[31]), .B(a[30]), .Z(n3105) );
  HS65_LH_NAND2X2 U3003 ( .A(a[31]), .B(n3104), .Z(n2673) );
  HS65_LHS_XOR2X3 U3004 ( .A(n2655), .B(a[30]), .Z(n3104) );
endmodule


module alu ( clk, rst_n, .alu_i({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , 
        \alu_i[SRC_B][31] , \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , 
        \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , 
        \alu_i[SRC_B][25] , \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , 
        \alu_i[SRC_B][22] , \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , 
        \alu_i[SRC_B][19] , \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , 
        \alu_i[SRC_B][16] , \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , 
        \alu_i[SRC_B][13] , \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , 
        \alu_i[SRC_B][10] , \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , 
        \alu_i[SRC_B][7] , \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , 
        \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , 
        \alu_i[SRC_B][1] , \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , 
        \alu_i[OP][2] , \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , 
        \alu_i[SHAMT][3] , \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , 
        \alu_i[SHAMT][0] }), .alu_o({\alu_o[BRANCH] , \alu_o[RESULT][31] , 
        \alu_o[RESULT][30] , \alu_o[RESULT][29] , \alu_o[RESULT][28] , 
        \alu_o[RESULT][27] , \alu_o[RESULT][26] , \alu_o[RESULT][25] , 
        \alu_o[RESULT][24] , \alu_o[RESULT][23] , \alu_o[RESULT][22] , 
        \alu_o[RESULT][21] , \alu_o[RESULT][20] , \alu_o[RESULT][19] , 
        \alu_o[RESULT][18] , \alu_o[RESULT][17] , \alu_o[RESULT][16] , 
        \alu_o[RESULT][15] , \alu_o[RESULT][14] , \alu_o[RESULT][13] , 
        \alu_o[RESULT][12] , \alu_o[RESULT][11] , \alu_o[RESULT][10] , 
        \alu_o[RESULT][9] , \alu_o[RESULT][8] , \alu_o[RESULT][7] , 
        \alu_o[RESULT][6] , \alu_o[RESULT][5] , \alu_o[RESULT][4] , 
        \alu_o[RESULT][3] , \alu_o[RESULT][2] , \alu_o[RESULT][1] , 
        \alu_o[RESULT][0] }) );
  input clk, rst_n, \alu_i[SRC_A][31] , \alu_i[SRC_A][30] , \alu_i[SRC_A][29] ,
         \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , \alu_i[SRC_A][26] ,
         \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , \alu_i[SRC_A][23] ,
         \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , \alu_i[SRC_A][20] ,
         \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , \alu_i[SRC_A][17] ,
         \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , \alu_i[SRC_A][14] ,
         \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , \alu_i[SRC_A][11] ,
         \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , \alu_i[SRC_A][8] ,
         \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , \alu_i[SRC_A][5] ,
         \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , \alu_i[SRC_A][2] ,
         \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , \alu_i[SRC_B][31] ,
         \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , \alu_i[SRC_B][28] ,
         \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , \alu_i[SRC_B][25] ,
         \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , \alu_i[SRC_B][22] ,
         \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , \alu_i[SRC_B][19] ,
         \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , \alu_i[SRC_B][16] ,
         \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , \alu_i[SRC_B][13] ,
         \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , \alu_i[SRC_B][10] ,
         \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , \alu_i[SRC_B][7] ,
         \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , \alu_i[SRC_B][4] ,
         \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , \alu_i[SRC_B][1] ,
         \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , \alu_i[OP][2] ,
         \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , \alu_i[SHAMT][3] ,
         \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , \alu_i[SHAMT][0] ;
  output \alu_o[BRANCH] , \alu_o[RESULT][31] , \alu_o[RESULT][30] ,
         \alu_o[RESULT][29] , \alu_o[RESULT][28] , \alu_o[RESULT][27] ,
         \alu_o[RESULT][26] , \alu_o[RESULT][25] , \alu_o[RESULT][24] ,
         \alu_o[RESULT][23] , \alu_o[RESULT][22] , \alu_o[RESULT][21] ,
         \alu_o[RESULT][20] , \alu_o[RESULT][19] , \alu_o[RESULT][18] ,
         \alu_o[RESULT][17] , \alu_o[RESULT][16] , \alu_o[RESULT][15] ,
         \alu_o[RESULT][14] , \alu_o[RESULT][13] , \alu_o[RESULT][12] ,
         \alu_o[RESULT][11] , \alu_o[RESULT][10] , \alu_o[RESULT][9] ,
         \alu_o[RESULT][8] , \alu_o[RESULT][7] , \alu_o[RESULT][6] ,
         \alu_o[RESULT][5] , \alu_o[RESULT][4] , \alu_o[RESULT][3] ,
         \alu_o[RESULT][2] , \alu_o[RESULT][1] , \alu_o[RESULT][0] ;
  wire   \HI_LO_c[HI][31] , \HI_LO_c[HI][30] , \HI_LO_c[HI][29] ,
         \HI_LO_c[HI][28] , \HI_LO_c[HI][27] , \HI_LO_c[HI][26] ,
         \HI_LO_c[HI][25] , \HI_LO_c[HI][24] , \HI_LO_c[HI][23] ,
         \HI_LO_c[HI][22] , \HI_LO_c[HI][21] , \HI_LO_c[HI][20] ,
         \HI_LO_c[HI][19] , \HI_LO_c[HI][18] , \HI_LO_c[HI][17] ,
         \HI_LO_c[HI][16] , \HI_LO_c[HI][15] , \HI_LO_c[HI][14] ,
         \HI_LO_c[HI][13] , \HI_LO_c[HI][12] , \HI_LO_c[HI][11] ,
         \HI_LO_c[HI][10] , \HI_LO_c[HI][9] , \HI_LO_c[HI][8] ,
         \HI_LO_c[HI][7] , \HI_LO_c[HI][6] , \HI_LO_c[HI][5] ,
         \HI_LO_c[HI][4] , \HI_LO_c[HI][3] , \HI_LO_c[HI][2] ,
         \HI_LO_c[HI][1] , \HI_LO_c[HI][0] , \HI_LO_c[LO][31] ,
         \HI_LO_c[LO][30] , \HI_LO_c[LO][29] , \HI_LO_c[LO][28] ,
         \HI_LO_c[LO][27] , \HI_LO_c[LO][26] , \HI_LO_c[LO][25] ,
         \HI_LO_c[LO][24] , \HI_LO_c[LO][23] , \HI_LO_c[LO][22] ,
         \HI_LO_c[LO][21] , \HI_LO_c[LO][20] , \HI_LO_c[LO][19] ,
         \HI_LO_c[LO][18] , \HI_LO_c[LO][17] , \HI_LO_c[LO][16] ,
         \HI_LO_c[LO][15] , \HI_LO_c[LO][14] , \HI_LO_c[LO][13] ,
         \HI_LO_c[LO][12] , \HI_LO_c[LO][11] , \HI_LO_c[LO][10] ,
         \HI_LO_c[LO][9] , \HI_LO_c[LO][8] , \HI_LO_c[LO][7] ,
         \HI_LO_c[LO][6] , \HI_LO_c[LO][5] , \HI_LO_c[LO][4] ,
         \HI_LO_c[LO][3] , \HI_LO_c[LO][2] , \HI_LO_c[LO][1] ,
         \HI_LO_c[LO][0] , N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N648, N649,
         N714, N715, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n300, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612;

  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][31]  ( .D(n516), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][30]  ( .D(n515), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][29]  ( .D(n514), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][28]  ( .D(n513), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][27]  ( .D(n512), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][26]  ( .D(n511), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][25]  ( .D(n510), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][24]  ( .D(n509), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][23]  ( .D(n508), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][22]  ( .D(n507), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][21]  ( .D(n506), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][20]  ( .D(n505), .CP(clk), .RN(n556), .Q(
        \HI_LO_c[HI][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][19]  ( .D(n504), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][18]  ( .D(n503), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][17]  ( .D(n502), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][16]  ( .D(n501), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][15]  ( .D(n500), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][14]  ( .D(n499), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][13]  ( .D(n498), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][12]  ( .D(n497), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][11]  ( .D(n496), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][10]  ( .D(n495), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][9]  ( .D(n494), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][8]  ( .D(n493), .CP(clk), .RN(n557), .Q(
        \HI_LO_c[HI][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][7]  ( .D(n492), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][6]  ( .D(n491), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][5]  ( .D(n490), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][4]  ( .D(n489), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][3]  ( .D(n488), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][2]  ( .D(n487), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][1]  ( .D(n486), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][0]  ( .D(n485), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[HI][0] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][31]  ( .D(n484), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[LO][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][30]  ( .D(n483), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[LO][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][29]  ( .D(n482), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[LO][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][28]  ( .D(n481), .CP(clk), .RN(n558), .Q(
        \HI_LO_c[LO][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][27]  ( .D(n480), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][26]  ( .D(n479), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][25]  ( .D(n478), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][24]  ( .D(n477), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][23]  ( .D(n476), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][22]  ( .D(n475), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][21]  ( .D(n474), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][20]  ( .D(n473), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][19]  ( .D(n472), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][18]  ( .D(n471), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][17]  ( .D(n470), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][16]  ( .D(n469), .CP(clk), .RN(n559), .Q(
        \HI_LO_c[LO][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][15]  ( .D(n468), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][14]  ( .D(n467), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][13]  ( .D(n466), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][12]  ( .D(n465), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][11]  ( .D(n464), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][10]  ( .D(n463), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][9]  ( .D(n462), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][8]  ( .D(n461), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][7]  ( .D(n460), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][6]  ( .D(n459), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][5]  ( .D(n458), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][4]  ( .D(n457), .CP(clk), .RN(n560), .Q(
        \HI_LO_c[LO][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][3]  ( .D(n456), .CP(clk), .RN(n561), .Q(
        \HI_LO_c[LO][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][2]  ( .D(n455), .CP(clk), .RN(n561), .Q(
        \HI_LO_c[LO][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][1]  ( .D(n454), .CP(clk), .RN(n561), .Q(
        \HI_LO_c[LO][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][0]  ( .D(n453), .CP(clk), .RN(n561), .Q(
        \HI_LO_c[LO][0] ) );
  alu_DW_cmp_0 lt_136 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , n552, 
        \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , n550, \alu_i[SRC_A][25] , 
        \alu_i[SRC_A][24] , n548, \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , n546, 
        \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , n544, \alu_i[SRC_A][16] , 
        \alu_i[SRC_A][15] , n542, \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , n540, 
        \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , n538, \alu_i[SRC_A][7] , 
        \alu_i[SRC_A][6] , n536, \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n534, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({n532, n531, n530, n528, 
        n526, n525, n524, n523, n522, n521, n520, n518, n517, n300, n90, n89, 
        n88, n87, n86, n85, n83, n82, n81, n80, n79, n78, n77, n75, n73, n71, 
        n70, n69}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(
        N648) );
  alu_DW01_sub_0 sub_68 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , n552, 
        \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , n550, \alu_i[SRC_A][25] , 
        \alu_i[SRC_A][24] , n548, \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , n546, 
        \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , n544, \alu_i[SRC_A][16] , 
        \alu_i[SRC_A][15] , n542, \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , n540, 
        \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , n538, \alu_i[SRC_A][7] , 
        \alu_i[SRC_A][6] , n536, \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n534, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({n532, n531, n530, n528, 
        n526, n525, n524, n523, n522, n521, n520, n518, n517, n300, n90, n89, 
        n88, n87, n86, n85, n83, n82, n81, n80, n79, n78, n77, n75, n73, n71, 
        n70, n69}), .CI(1'b0), .DIFF({N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131}) );
  alu_DW01_cmp6_0 r325 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , n552, 
        \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , n550, \alu_i[SRC_A][25] , 
        \alu_i[SRC_A][24] , n548, \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , n546, 
        \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , n544, \alu_i[SRC_A][16] , 
        \alu_i[SRC_A][15] , n542, \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , n540, 
        \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , n538, \alu_i[SRC_A][7] , 
        \alu_i[SRC_A][6] , n536, \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n534, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({n532, n531, n530, n528, 
        n526, n525, n524, n523, n522, n521, n520, n518, n517, n300, n90, n89, 
        n88, n87, n86, n85, n83, n82, n81, n80, n79, n78, n77, n75, n73, n71, 
        n70, n69}), .TC(1'b0), .LT(N649), .EQ(N714), .NE(N715) );
  alu_DW01_add_0 r321 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , n552, 
        \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , n550, \alu_i[SRC_A][25] , 
        \alu_i[SRC_A][24] , n548, \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , n546, 
        \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , n544, \alu_i[SRC_A][16] , 
        \alu_i[SRC_A][15] , n542, \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , n540, 
        \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , n538, \alu_i[SRC_A][7] , 
        \alu_i[SRC_A][6] , n536, \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n534, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({n532, n531, n530, n528, 
        n526, n525, n524, n523, n522, n521, n520, n518, n517, n300, n90, n89, 
        n88, n87, n86, n85, n83, n82, n81, n80, n79, n78, n77, n75, n73, n71, 
        n70, n69}), .CI(1'b0), .SUM({N130, N129, N128, N127, N126, N125, N124, 
        N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, 
        N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, 
        N99}) );
  alu_DW_mult_uns_0 mult_71 ( .a({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , n552, 
        \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , n550, \alu_i[SRC_A][25] , 
        \alu_i[SRC_A][24] , n548, \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , n546, 
        \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , n544, \alu_i[SRC_A][16] , 
        \alu_i[SRC_A][15] , n542, \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , n540, 
        \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , n538, \alu_i[SRC_A][7] , 
        \alu_i[SRC_A][6] , n536, \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , n534, 
        \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .b({n532, n531, n530, n528, 
        n526, n525, n524, n523, n522, n521, n520, n518, n517, n300, n90, n89, 
        n88, n87, n86, n85, n83, n82, n81, n80, n79, n78, n77, n75, n73, n71, 
        n70, n69}), .product({N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163}) );
  HS65_LH_NOR4ABX2 U3 ( .A(n92), .B(n93), .C(n94), .D(n95), .Z(n91) );
  HS65_LH_IVX9 U4 ( .A(n537), .Z(n536) );
  HS65_LH_IVX9 U5 ( .A(n76), .Z(n75) );
  HS65_LH_IVX9 U6 ( .A(n74), .Z(n73) );
  HS65_LH_IVX9 U7 ( .A(n541), .Z(n540) );
  HS65_LH_IVX9 U13 ( .A(n545), .Z(n544) );
  HS65_LH_IVX9 U14 ( .A(n539), .Z(n538) );
  HS65_LH_IVX9 U15 ( .A(n543), .Z(n542) );
  HS65_LH_IVX9 U16 ( .A(n72), .Z(n71) );
  HS65_LH_IVX9 U17 ( .A(n84), .Z(n83) );
  HS65_LH_IVX9 U18 ( .A(n547), .Z(n546) );
  HS65_LH_IVX9 U19 ( .A(n551), .Z(n550) );
  HS65_LH_IVX9 U20 ( .A(n553), .Z(n552) );
  HS65_LH_IVX9 U21 ( .A(n519), .Z(n518) );
  HS65_LH_IVX9 U22 ( .A(n527), .Z(n526) );
  HS65_LH_IVX9 U23 ( .A(n529), .Z(n528) );
  HS65_LH_IVX9 U24 ( .A(n533), .Z(n532) );
  HS65_LH_NOR4ABX4 U25 ( .A(n612), .B(n435), .C(\alu_i[OP][3] ), .D(
        \alu_i[OP][2] ), .Z(n180) );
  HS65_LH_BFX9 U26 ( .A(\alu_i[SRC_B][1] ), .Z(n70) );
  HS65_LH_BFX9 U27 ( .A(\alu_i[SRC_B][8] ), .Z(n80) );
  HS65_LH_BFX9 U28 ( .A(\alu_i[SRC_B][5] ), .Z(n77) );
  HS65_LH_BFX9 U29 ( .A(\alu_i[SRC_B][6] ), .Z(n78) );
  HS65_LH_BFX9 U30 ( .A(\alu_i[SRC_B][7] ), .Z(n79) );
  HS65_LH_BFX9 U31 ( .A(\alu_i[SRC_B][10] ), .Z(n82) );
  HS65_LH_BFX9 U32 ( .A(\alu_i[SRC_B][12] ), .Z(n85) );
  HS65_LH_BFX9 U33 ( .A(\alu_i[SRC_B][13] ), .Z(n86) );
  HS65_LH_BFX9 U34 ( .A(\alu_i[SRC_B][14] ), .Z(n87) );
  HS65_LH_BFX9 U35 ( .A(\alu_i[SRC_B][15] ), .Z(n88) );
  HS65_LH_BFX9 U36 ( .A(\alu_i[SRC_B][9] ), .Z(n81) );
  HS65_LH_BFX9 U37 ( .A(\alu_i[SRC_B][19] ), .Z(n517) );
  HS65_LH_BFX9 U38 ( .A(\alu_i[SRC_B][16] ), .Z(n89) );
  HS65_LH_BFX9 U39 ( .A(\alu_i[SRC_B][17] ), .Z(n90) );
  HS65_LH_BFX9 U40 ( .A(\alu_i[SRC_B][18] ), .Z(n300) );
  HS65_LH_BFX9 U41 ( .A(\alu_i[SRC_B][21] ), .Z(n520) );
  HS65_LH_BFX9 U42 ( .A(\alu_i[SRC_B][23] ), .Z(n522) );
  HS65_LH_BFX9 U43 ( .A(\alu_i[SRC_B][25] ), .Z(n524) );
  HS65_LH_BFX9 U44 ( .A(\alu_i[SRC_B][22] ), .Z(n521) );
  HS65_LH_BFX9 U45 ( .A(\alu_i[SRC_B][24] ), .Z(n523) );
  HS65_LH_BFX9 U46 ( .A(\alu_i[SRC_B][26] ), .Z(n525) );
  HS65_LH_BFX9 U47 ( .A(\alu_i[SRC_B][29] ), .Z(n530) );
  HS65_LH_BFX9 U48 ( .A(\alu_i[SRC_B][30] ), .Z(n531) );
  HS65_LH_NOR2X6 U49 ( .A(n98), .B(\alu_i[SHAMT][4] ), .Z(n284) );
  HS65_LH_IVX9 U50 ( .A(n61), .Z(n60) );
  HS65_LH_IVX9 U51 ( .A(n61), .Z(n59) );
  HS65_LH_IVX9 U52 ( .A(n62), .Z(n58) );
  HS65_LH_IVX9 U53 ( .A(n62), .Z(n57) );
  HS65_LH_IVX9 U54 ( .A(n98), .Z(n605) );
  HS65_LH_IVX9 U55 ( .A(n56), .Z(n55) );
  HS65_LH_IVX9 U56 ( .A(n42), .Z(n41) );
  HS65_LH_IVX9 U57 ( .A(n42), .Z(n40) );
  HS65_LH_BFX9 U58 ( .A(n68), .Z(n61) );
  HS65_LH_BFX9 U59 ( .A(n68), .Z(n62) );
  HS65_LH_BFX9 U60 ( .A(n604), .Z(n12) );
  HS65_LH_BFX9 U61 ( .A(n604), .Z(n11) );
  HS65_LH_BFX9 U62 ( .A(n603), .Z(n8) );
  HS65_LH_BFX9 U63 ( .A(n603), .Z(n9) );
  HS65_LH_BFX9 U64 ( .A(n67), .Z(n65) );
  HS65_LH_BFX9 U65 ( .A(n67), .Z(n64) );
  HS65_LH_BFX9 U66 ( .A(n68), .Z(n63) );
  HS65_LH_BFX9 U67 ( .A(n604), .Z(n13) );
  HS65_LH_BFX9 U68 ( .A(n603), .Z(n10) );
  HS65_LH_BFX9 U69 ( .A(n67), .Z(n66) );
  HS65_LH_BFX9 U70 ( .A(n555), .Z(n560) );
  HS65_LH_BFX9 U71 ( .A(n555), .Z(n559) );
  HS65_LH_BFX9 U72 ( .A(n554), .Z(n558) );
  HS65_LH_BFX9 U73 ( .A(n554), .Z(n557) );
  HS65_LH_BFX9 U74 ( .A(n554), .Z(n556) );
  HS65_LH_BFX9 U75 ( .A(n555), .Z(n561) );
  HS65_LH_IVX9 U76 ( .A(n101), .Z(n603) );
  HS65_LH_IVX9 U77 ( .A(n100), .Z(n604) );
  HS65_LH_NAND2X7 U78 ( .A(n442), .B(n435), .Z(n98) );
  HS65_LH_IVX9 U79 ( .A(n96), .Z(n606) );
  HS65_LH_NOR3X4 U80 ( .A(n48), .B(n45), .C(n106), .Z(n92) );
  HS65_LH_IVX9 U81 ( .A(n176), .Z(n597) );
  HS65_LH_IVX9 U82 ( .A(n281), .Z(n598) );
  HS65_LH_IVX9 U83 ( .A(n54), .Z(n56) );
  HS65_LH_IVX9 U84 ( .A(n39), .Z(n42) );
  HS65_LH_BFX9 U85 ( .A(n43), .Z(n44) );
  HS65_LH_BFX9 U86 ( .A(n91), .Z(n68) );
  HS65_LH_BFX9 U87 ( .A(n91), .Z(n67) );
  HS65_LH_BFX9 U88 ( .A(n50), .Z(n52) );
  HS65_LH_BFX9 U89 ( .A(n50), .Z(n51) );
  HS65_LH_BFX9 U90 ( .A(n608), .Z(n15) );
  HS65_LH_BFX9 U91 ( .A(n608), .Z(n14) );
  HS65_LH_BFX9 U92 ( .A(n43), .Z(n45) );
  HS65_LH_BFX9 U93 ( .A(n50), .Z(n53) );
  HS65_LH_BFX9 U94 ( .A(rst_n), .Z(n555) );
  HS65_LH_BFX9 U95 ( .A(rst_n), .Z(n554) );
  HS65_LH_IVX9 U96 ( .A(n237), .Z(n592) );
  HS65_LH_AO222X4 U97 ( .A(n128), .B(n115), .C(n133), .D(n118), .E(n174), .F(
        n117), .Z(n170) );
  HS65_LH_IVX9 U98 ( .A(n317), .Z(n582) );
  HS65_LH_IVX9 U99 ( .A(n144), .Z(n572) );
  HS65_LH_IVX9 U100 ( .A(n130), .Z(n579) );
  HS65_LH_IVX9 U101 ( .A(n212), .Z(n575) );
  HS65_LH_NOR4ABX2 U102 ( .A(n100), .B(n101), .C(n102), .D(n103), .Z(n93) );
  HS65_LH_NAND3X5 U103 ( .A(n96), .B(n54), .C(n98), .Z(n95) );
  HS65_LH_NAND4ABX3 U104 ( .A(n42), .B(n53), .C(n612), .D(n15), .Z(n94) );
  HS65_LH_NOR2X6 U105 ( .A(n96), .B(n189), .Z(n279) );
  HS65_LH_IVX9 U106 ( .A(n180), .Z(n608) );
  HS65_LH_NAND2X7 U107 ( .A(n436), .B(n442), .Z(n96) );
  HS65_LH_NOR2X6 U108 ( .A(n189), .B(n98), .Z(n115) );
  HS65_LH_NOR2X6 U109 ( .A(n611), .B(n609), .Z(n435) );
  HS65_LH_IVX9 U110 ( .A(n208), .Z(n600) );
  HS65_LH_AND2X4 U111 ( .A(n390), .B(n391), .Z(n106) );
  HS65_LH_IVX9 U112 ( .A(n186), .Z(n599) );
  HS65_LH_NAND2X7 U113 ( .A(n195), .B(n605), .Z(n176) );
  HS65_LH_AND2X4 U114 ( .A(n445), .B(n607), .Z(n442) );
  HS65_LH_NAND2X7 U115 ( .A(n606), .B(n195), .Z(n281) );
  HS65_LH_IVX9 U116 ( .A(n189), .Z(n595) );
  HS65_LH_NAND2X7 U117 ( .A(n434), .B(n438), .Z(n101) );
  HS65_LH_AND2X4 U118 ( .A(n275), .B(n16), .Z(n368) );
  HS65_LH_AND2X4 U119 ( .A(n117), .B(n16), .Z(n397) );
  HS65_LH_NAND2X7 U120 ( .A(n434), .B(n435), .Z(n100) );
  HS65_LH_BFX9 U121 ( .A(n123), .Z(n39) );
  HS65_LH_NAND2X7 U122 ( .A(n438), .B(n442), .Z(n123) );
  HS65_LH_BFX9 U123 ( .A(n97), .Z(n54) );
  HS65_LH_NAND2X7 U124 ( .A(n391), .B(n442), .Z(n97) );
  HS65_LH_IVX9 U125 ( .A(n438), .Z(n610) );
  HS65_LH_BFX9 U126 ( .A(n105), .Z(n43) );
  HS65_LH_NOR2AX3 U127 ( .A(n390), .B(n610), .Z(n105) );
  HS65_LH_BFX9 U128 ( .A(n99), .Z(n50) );
  HS65_LH_NOR2X6 U129 ( .A(n609), .B(n437), .Z(n99) );
  HS65_LH_IVX9 U130 ( .A(n38), .Z(n36) );
  HS65_LH_BFX9 U131 ( .A(n46), .Z(n48) );
  HS65_LH_BFX9 U132 ( .A(n46), .Z(n47) );
  HS65_LH_AND2X4 U133 ( .A(n434), .B(n391), .Z(n102) );
  HS65_LH_BFX9 U134 ( .A(n29), .Z(n31) );
  HS65_LH_BFX9 U135 ( .A(n29), .Z(n32) );
  HS65_LH_BFX9 U136 ( .A(n30), .Z(n33) );
  HS65_LH_IVX9 U137 ( .A(n38), .Z(n37) );
  HS65_LH_AND2X4 U138 ( .A(n434), .B(n436), .Z(n103) );
  HS65_LH_BFX9 U139 ( .A(n18), .Z(n20) );
  HS65_LH_BFX9 U140 ( .A(n18), .Z(n22) );
  HS65_LH_BFX9 U141 ( .A(n18), .Z(n21) );
  HS65_LH_BFX9 U142 ( .A(n19), .Z(n23) );
  HS65_LH_BFX9 U143 ( .A(n19), .Z(n24) );
  HS65_LH_BFX9 U144 ( .A(n46), .Z(n49) );
  HS65_LH_BFX9 U145 ( .A(n30), .Z(n34) );
  HS65_LH_IVX9 U146 ( .A(n535), .Z(n534) );
  HS65_LH_IVX9 U147 ( .A(n549), .Z(n548) );
  HS65_LH_AO112X9 U148 ( .A(N714), .B(n450), .C(n451), .D(n452), .Z(
        \alu_o[BRANCH] ) );
  HS65_LH_AO222X4 U149 ( .A(n391), .B(n450), .C(n438), .D(n450), .E(n436), .F(
        n450), .Z(n452) );
  HS65_LH_NOR3X4 U150 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][3] ), .C(n612), .Z(
        n450) );
  HS65_LH_NOR4ABX2 U151 ( .A(N715), .B(n607), .C(n612), .D(n610), .Z(n451) );
  HS65_LH_AOI222X2 U152 ( .A(n31), .B(n70), .C(n26), .D(n69), .E(n35), .F(n71), 
        .Z(n237) );
  HS65_LH_AOI212X4 U153 ( .A(\alu_i[SRC_A][4] ), .B(n180), .C(n56), .D(n589), 
        .E(n42), .Z(n175) );
  HS65_LH_IVX9 U154 ( .A(\alu_i[SRC_A][4] ), .Z(n589) );
  HS65_LH_AOI212X4 U155 ( .A(n540), .B(n180), .C(n56), .D(n541), .E(n42), .Z(
        n421) );
  HS65_LH_AOI212X4 U156 ( .A(n546), .B(n180), .C(n56), .D(n547), .E(n42), .Z(
        n350) );
  HS65_LH_AOI212X4 U157 ( .A(\alu_i[SRC_A][27] ), .B(n180), .C(n56), .D(n567), 
        .E(n42), .Z(n280) );
  HS65_LH_IVX9 U158 ( .A(\alu_i[SRC_A][27] ), .Z(n567) );
  HS65_LH_OAI212X5 U159 ( .A(n585), .B(n189), .C(n190), .D(n596), .E(n191), 
        .Z(n183) );
  HS65_LH_IVX9 U160 ( .A(n140), .Z(n585) );
  HS65_LH_AOI222X2 U161 ( .A(n192), .B(n145), .C(n193), .D(n194), .E(n195), 
        .F(n142), .Z(n191) );
  HS65_LH_MX41X7 U162 ( .D0(n73), .S0(n36), .D1(n75), .S1(n32), .D2(n77), .S2(
        n27), .D3(n78), .S3(n22), .Z(n194) );
  HS65_LH_OAI212X5 U163 ( .A(n570), .B(n189), .C(n264), .D(n596), .E(n265), 
        .Z(n259) );
  HS65_LH_IVX9 U164 ( .A(n269), .Z(n570) );
  HS65_LH_AOI222X2 U165 ( .A(n192), .B(n266), .C(n193), .D(n267), .E(n195), 
        .F(n268), .Z(n265) );
  HS65_LH_MX41X7 U166 ( .D0(n528), .S0(n196), .D1(n526), .S1(n31), .D2(n525), 
        .S2(n26), .D3(n524), .S3(n20), .Z(n267) );
  HS65_LH_OAI212X5 U167 ( .A(n236), .B(n72), .C(n237), .D(n186), .E(n238), .Z(
        n235) );
  HS65_LH_CBI4I1X5 U168 ( .A(n56), .B(n72), .C(n42), .D(n534), .Z(n238) );
  HS65_LH_AOI212X4 U169 ( .A(n534), .B(n180), .C(n56), .D(n535), .E(n42), .Z(
        n236) );
  HS65_LH_OAI212X5 U170 ( .A(n185), .B(n74), .C(n591), .D(n186), .E(n187), .Z(
        n184) );
  HS65_LH_CBI4I1X5 U171 ( .A(n56), .B(n74), .C(n42), .D(\alu_i[SRC_A][3] ), 
        .Z(n187) );
  HS65_LH_AOI212X4 U172 ( .A(\alu_i[SRC_A][3] ), .B(n180), .C(n56), .D(n590), 
        .E(n42), .Z(n185) );
  HS65_LH_IVX9 U173 ( .A(n188), .Z(n591) );
  HS65_LH_OAI212X5 U174 ( .A(n261), .B(n529), .C(n564), .D(n208), .E(n262), 
        .Z(n260) );
  HS65_LH_CBI4I1X5 U175 ( .A(n56), .B(n529), .C(n42), .D(\alu_i[SRC_A][28] ), 
        .Z(n262) );
  HS65_LH_AOI212X4 U176 ( .A(\alu_i[SRC_A][28] ), .B(n180), .C(n56), .D(n566), 
        .E(n42), .Z(n261) );
  HS65_LH_IVX9 U177 ( .A(n263), .Z(n564) );
  HS65_LH_OAI212X5 U178 ( .A(n552), .B(n97), .C(n14), .D(n553), .E(n41), .Z(
        n248) );
  HS65_LH_AOI32X5 U179 ( .A(n283), .B(n601), .C(n284), .D(\alu_i[SRC_A][27] ), 
        .E(n285), .Z(n282) );
  HS65_LH_OAI21X3 U180 ( .A(n526), .B(n55), .C(n41), .Z(n285) );
  HS65_LH_OAI212X5 U181 ( .A(\alu_i[SRC_A][16] ), .B(n55), .C(n15), .D(n577), 
        .E(n41), .Z(n388) );
  HS65_LH_IVX9 U182 ( .A(\alu_i[SRC_A][16] ), .Z(n577) );
  HS65_LH_OAI212X5 U183 ( .A(\alu_i[SRC_A][15] ), .B(n55), .C(n15), .D(n578), 
        .E(n40), .Z(n396) );
  HS65_LH_IVX9 U184 ( .A(\alu_i[SRC_A][15] ), .Z(n578) );
  HS65_LH_OAI212X5 U185 ( .A(\alu_i[SRC_A][12] ), .B(n55), .C(n15), .D(n581), 
        .E(n40), .Z(n415) );
  HS65_LH_IVX9 U186 ( .A(\alu_i[SRC_A][12] ), .Z(n581) );
  HS65_LH_OAI212X5 U187 ( .A(\alu_i[SRC_A][13] ), .B(n55), .C(n15), .D(n580), 
        .E(n40), .Z(n409) );
  HS65_LH_IVX9 U188 ( .A(\alu_i[SRC_A][13] ), .Z(n580) );
  HS65_LH_OAI212X5 U189 ( .A(n542), .B(n55), .C(n15), .D(n543), .E(n40), .Z(
        n403) );
  HS65_LH_OAI212X5 U190 ( .A(n544), .B(n55), .C(n15), .D(n545), .E(n123), .Z(
        n381) );
  HS65_LH_OAI212X5 U191 ( .A(\alu_i[SRC_A][19] ), .B(n55), .C(n15), .D(n574), 
        .E(n40), .Z(n367) );
  HS65_LH_IVX9 U192 ( .A(\alu_i[SRC_A][19] ), .Z(n574) );
  HS65_LH_OAI212X5 U193 ( .A(\alu_i[SRC_A][22] ), .B(n55), .C(n14), .D(n571), 
        .E(n41), .Z(n338) );
  HS65_LH_IVX9 U194 ( .A(\alu_i[SRC_A][22] ), .Z(n571) );
  HS65_LH_OAI212X5 U195 ( .A(n536), .B(n54), .C(n14), .D(n537), .E(n41), .Z(
        n167) );
  HS65_LH_OAI212X5 U196 ( .A(\alu_i[SRC_A][7] ), .B(n54), .C(n14), .D(n587), 
        .E(n41), .Z(n146) );
  HS65_LH_IVX9 U197 ( .A(\alu_i[SRC_A][7] ), .Z(n587) );
  HS65_LH_OAI212X5 U198 ( .A(n538), .B(n54), .C(n14), .D(n539), .E(n41), .Z(
        n134) );
  HS65_LH_OAI212X5 U199 ( .A(\alu_i[SRC_A][9] ), .B(n54), .C(n586), .D(n15), 
        .E(n41), .Z(n121) );
  HS65_LH_IVX9 U200 ( .A(\alu_i[SRC_A][9] ), .Z(n586) );
  HS65_LH_OAI212X5 U201 ( .A(n548), .B(n54), .C(n14), .D(n549), .E(n41), .Z(
        n328) );
  HS65_LH_OAI212X5 U202 ( .A(n550), .B(n54), .C(n14), .D(n551), .E(n41), .Z(
        n293) );
  HS65_LH_OAI212X5 U203 ( .A(\alu_i[SRC_A][10] ), .B(n55), .C(n15), .D(n584), 
        .E(n41), .Z(n428) );
  HS65_LH_IVX9 U204 ( .A(\alu_i[SRC_A][10] ), .Z(n584) );
  HS65_LH_OAI212X5 U205 ( .A(\alu_i[SRC_A][25] ), .B(n55), .C(n14), .D(n568), 
        .E(n41), .Z(n307) );
  HS65_LH_IVX9 U206 ( .A(\alu_i[SRC_A][25] ), .Z(n568) );
  HS65_LH_AOI32X5 U207 ( .A(n178), .B(n601), .C(n275), .D(n546), .E(n352), .Z(
        n351) );
  HS65_LH_OAI21X3 U208 ( .A(n518), .B(n55), .C(n123), .Z(n352) );
  HS65_LH_AOI32X5 U209 ( .A(n178), .B(n601), .C(n113), .D(\alu_i[SRC_A][4] ), 
        .E(n179), .Z(n177) );
  HS65_LH_OAI21X3 U210 ( .A(n75), .B(n55), .C(n39), .Z(n179) );
  HS65_LH_AOI32X5 U211 ( .A(n283), .B(n601), .C(n117), .D(n540), .E(n423), .Z(
        n422) );
  HS65_LH_OAI21X3 U212 ( .A(n83), .B(n55), .C(n40), .Z(n423) );
  HS65_LH_MX41X7 U213 ( .D0(n85), .S0(n37), .D1(n83), .S1(n33), .D2(n82), .S2(
        n28), .D3(n20), .S3(n81), .Z(n317) );
  HS65_LH_MX41X7 U214 ( .D0(n80), .S0(n37), .D1(n79), .S1(n33), .D2(n78), .S2(
        n27), .D3(n77), .S3(n22), .Z(n316) );
  HS65_LH_MX41X7 U215 ( .D0(n88), .S0(n37), .D1(n89), .S1(n33), .D2(n90), .S2(
        n28), .D3(n300), .S3(n23), .Z(n145) );
  HS65_LH_MX41X7 U216 ( .D0(n89), .S0(n36), .D1(n88), .S1(n32), .D2(n87), .S2(
        n27), .D3(n86), .S3(n21), .Z(n266) );
  HS65_LH_MX41X7 U217 ( .D0(n88), .S0(n36), .D1(n87), .S1(n32), .D2(n86), .S2(
        n27), .D3(n85), .S3(n21), .Z(n278) );
  HS65_LH_NOR2AX3 U218 ( .A(n69), .B(n38), .Z(n315) );
  HS65_LH_MX41X7 U219 ( .D0(n196), .S0(n517), .D1(n31), .S1(n518), .D2(n520), 
        .S2(n28), .D3(n521), .S3(n23), .Z(n144) );
  HS65_LH_MX41X7 U220 ( .D0(n528), .S0(n37), .D1(n530), .S1(n33), .D2(n531), 
        .S2(n28), .D3(n532), .S3(n24), .Z(n263) );
  HS65_LH_MX41X7 U221 ( .D0(n73), .S0(n37), .D1(n71), .S1(n33), .D2(n70), .S2(
        n28), .D3(n69), .S3(n23), .Z(n188) );
  HS65_LH_MX41X7 U222 ( .D0(n85), .S0(n37), .D1(n86), .S1(n33), .D2(n87), .S2(
        n28), .D3(n88), .S3(n24), .Z(n130) );
  HS65_LH_MX41X7 U223 ( .D0(n35), .S0(n517), .D1(n300), .S1(n32), .D2(n90), 
        .S2(n27), .D3(n89), .S3(n21), .Z(n212) );
  HS65_LH_MX41X7 U224 ( .D0(n522), .S0(n37), .D1(n523), .S1(n33), .D2(n524), 
        .S2(n28), .D3(n525), .S3(n23), .Z(n325) );
  HS65_LH_MX41X7 U225 ( .D0(n87), .S0(n37), .D1(n88), .S1(n33), .D2(n89), .S2(
        n28), .D3(n90), .S3(n23), .Z(n157) );
  HS65_LH_MX41X7 U226 ( .D0(n86), .S0(n36), .D1(n87), .S1(n32), .D2(n88), .S2(
        n27), .D3(n89), .S3(n22), .Z(n114) );
  HS65_LH_MX41X7 U227 ( .D0(n83), .S0(n37), .D1(n85), .S1(n33), .D2(n86), .S2(
        n28), .D3(n87), .S3(n22), .Z(n142) );
  HS65_LH_MX41X7 U228 ( .D0(n77), .S0(n36), .D1(n75), .S1(n32), .D2(n73), .S2(
        n27), .D3(n71), .S3(n22), .Z(n302) );
  HS65_LH_MX41X7 U229 ( .D0(n78), .S0(n37), .D1(n77), .S1(n33), .D2(n75), .S2(
        n28), .D3(n73), .S3(n23), .Z(n336) );
  HS65_LH_MX41X7 U230 ( .D0(n79), .S0(n37), .D1(n78), .S1(n33), .D2(n77), .S2(
        n28), .D3(n75), .S3(n23), .Z(n326) );
  HS65_LH_MX41X7 U231 ( .D0(n35), .S0(n300), .D1(n90), .S1(n32), .D2(n89), 
        .S2(n27), .D3(n88), .S3(n21), .Z(n229) );
  HS65_LH_MX41X7 U232 ( .D0(n196), .S0(n518), .D1(n31), .S1(n517), .D2(n300), 
        .S2(n27), .D3(n90), .S3(n21), .Z(n268) );
  HS65_LH_MX41X7 U233 ( .D0(n90), .S0(n36), .D1(n89), .S1(n32), .D2(n88), .S2(
        n27), .D3(n87), .S3(n21), .Z(n254) );
  HS65_LH_MX41X7 U234 ( .D0(n87), .S0(n36), .D1(n86), .S1(n32), .D2(n85), .S2(
        n27), .D3(n83), .S3(n22), .Z(n292) );
  HS65_LH_MX41X7 U235 ( .D0(n86), .S0(n36), .D1(n85), .S1(n32), .D2(n83), .S2(
        n27), .D3(n82), .S3(n22), .Z(n306) );
  HS65_LH_CBI4I6X5 U236 ( .A(n530), .B(n54), .C(n40), .D(n553), .Z(n249) );
  HS65_LH_AO222X4 U237 ( .A(n33), .B(n531), .C(n26), .D(n532), .E(n35), .F(
        n530), .Z(n247) );
  HS65_LH_NOR2X6 U238 ( .A(n533), .B(n38), .Z(n216) );
  HS65_LH_MX41X7 U239 ( .D0(n523), .S0(n37), .D1(n524), .S1(n33), .D2(n525), 
        .S2(n28), .D3(n526), .S3(n24), .Z(n313) );
  HS65_LH_MX41X7 U240 ( .D0(n196), .S0(n81), .D1(n82), .S1(n32), .D2(n83), 
        .S2(n27), .D3(n85), .S3(n21), .Z(n111) );
  HS65_LH_MX41X7 U241 ( .D0(n82), .S0(n37), .D1(n83), .S1(n33), .D2(n85), .S2(
        n28), .D3(n86), .S3(n23), .Z(n154) );
  HS65_LH_MX41X7 U242 ( .D0(n524), .S0(n36), .D1(n525), .S1(n32), .D2(n526), 
        .S2(n27), .D3(n528), .S3(n22), .Z(n299) );
  HS65_LH_MX41X7 U243 ( .D0(n525), .S0(n37), .D1(n526), .S1(n33), .D2(n528), 
        .S2(n28), .D3(n530), .S3(n23), .Z(n334) );
  HS65_LH_MX41X7 U244 ( .D0(n89), .S0(n35), .D1(n90), .S1(n33), .D2(n300), 
        .S2(n28), .D3(n517), .S3(n24), .Z(n133) );
  HS65_LH_MX41X7 U245 ( .D0(n35), .S0(n518), .D1(n520), .S1(n33), .D2(n521), 
        .S2(n28), .D3(n522), .S3(n24), .Z(n132) );
  HS65_LH_MX41X7 U246 ( .D0(n521), .S0(n36), .D1(n520), .S1(n32), .D2(n26), 
        .S2(n518), .D3(n517), .S3(n21), .Z(n231) );
  HS65_LH_MX41X7 U247 ( .D0(n521), .S0(n37), .D1(n522), .S1(n33), .D2(n523), 
        .S2(n28), .D3(n524), .S3(n23), .Z(n335) );
  HS65_LH_MX41X7 U248 ( .D0(n82), .S0(n37), .D1(n31), .S1(n81), .D2(n80), .S2(
        n28), .D3(n79), .S3(n23), .Z(n337) );
  HS65_LH_MX41X7 U249 ( .D0(n520), .S0(n36), .D1(n521), .S1(n32), .D2(n522), 
        .S2(n27), .D3(n523), .S3(n22), .Z(n119) );
  HS65_LH_MX41X7 U250 ( .D0(n520), .S0(n36), .D1(n31), .S1(n518), .D2(n517), 
        .S2(n26), .D3(n300), .S3(n21), .Z(n256) );
  HS65_LH_MX41X7 U251 ( .D0(n35), .S0(n81), .D1(n80), .S1(n32), .D2(n79), .S2(
        n27), .D3(n78), .S3(n22), .Z(n305) );
  HS65_LH_MX41X7 U252 ( .D0(n83), .S0(n37), .D1(n82), .S1(n33), .D2(n26), .S2(
        n81), .D3(n80), .S3(n22), .Z(n327) );
  HS65_LH_MX41X7 U253 ( .D0(n75), .S0(n37), .D1(n73), .S1(n32), .D2(n71), .S2(
        n27), .D3(n70), .S3(n22), .Z(n314) );
  HS65_LH_MX41X7 U254 ( .D0(n90), .S0(n36), .D1(n300), .S1(n32), .D2(n517), 
        .S2(n27), .D3(n518), .S3(n22), .Z(n120) );
  HS65_LH_MX41X7 U255 ( .D0(n196), .S0(n300), .D1(n31), .S1(n517), .D2(n26), 
        .S2(n518), .D3(n520), .S3(n23), .Z(n156) );
  HS65_LH_MX41X7 U256 ( .D0(n80), .S0(n37), .D1(n31), .S1(n81), .D2(n82), .S2(
        n28), .D3(n83), .S3(n24), .Z(n128) );
  HS65_LH_MX41X7 U257 ( .D0(n522), .S0(n36), .D1(n521), .S1(n31), .D2(n520), 
        .S2(n26), .D3(n518), .S3(n21), .Z(n214) );
  HS65_LH_MX41X7 U258 ( .D0(n79), .S0(n36), .D1(n80), .S1(n31), .D2(n26), .S2(
        n81), .D3(n82), .S3(n20), .Z(n140) );
  HS65_LH_AO22X9 U259 ( .A(n35), .B(n70), .C(n31), .D(n69), .Z(n303) );
  HS65_LH_AO22X9 U260 ( .A(n35), .B(n531), .C(n31), .D(n532), .Z(n222) );
  HS65_LH_MX41X7 U261 ( .D0(n526), .S0(n37), .D1(n528), .S1(n33), .D2(n530), 
        .S2(n28), .D3(n531), .S3(n23), .Z(n324) );
  HS65_LH_MX41X7 U262 ( .D0(n16), .S0(n133), .D1(n7), .S1(n132), .D2(n304), 
        .S2(n313), .D3(n374), .S3(n263), .Z(n387) );
  HS65_LH_MX41X7 U263 ( .D0(n16), .S0(n120), .D1(n7), .S1(n119), .D2(n304), 
        .S2(n299), .D3(n374), .S3(n247), .Z(n360) );
  HS65_LH_MX41X7 U264 ( .D0(n16), .S0(n156), .D1(n301), .S1(n335), .D2(n304), 
        .S2(n334), .D3(n374), .S3(n222), .Z(n239) );
  HS65_LH_MX41X7 U265 ( .D0(n75), .S0(n196), .D1(n77), .S1(n31), .D2(n78), 
        .S2(n26), .D3(n79), .S3(n20), .Z(n173) );
  HS65_LH_MX41X7 U266 ( .D0(n77), .S0(n36), .D1(n78), .S1(n32), .D2(n79), .S2(
        n27), .D3(n80), .S3(n21), .Z(n164) );
  HS65_LH_MX41X7 U267 ( .D0(n78), .S0(n36), .D1(n79), .S1(n31), .D2(n80), .S2(
        n26), .D3(n20), .S3(n81), .Z(n152) );
  HS65_LH_OAI21X3 U268 ( .A(n205), .B(n533), .C(n206), .Z(n204) );
  HS65_LH_AOI212X4 U269 ( .A(n56), .B(n562), .C(\alu_i[SRC_A][31] ), .D(n180), 
        .E(n207), .Z(n205) );
  HS65_LH_CBI4I1X5 U270 ( .A(n56), .B(n533), .C(n42), .D(\alu_i[SRC_A][31] ), 
        .Z(n206) );
  HS65_LH_OAI211X5 U271 ( .A(n38), .B(n208), .C(n101), .D(n39), .Z(n207) );
  HS65_LH_AO222X4 U272 ( .A(n313), .B(n7), .C(n263), .D(n304), .E(n132), .F(
        n16), .Z(n174) );
  HS65_LH_AO222X4 U273 ( .A(n326), .B(n301), .C(n188), .D(n304), .E(n327), .F(
        n16), .Z(n276) );
  HS65_LH_AO222X4 U274 ( .A(n314), .B(n7), .C(n304), .D(n315), .E(n316), .F(
        n17), .Z(n129) );
  HS65_LH_AO222X4 U275 ( .A(n302), .B(n301), .C(n303), .D(n304), .E(n305), .F(
        n17), .Z(n112) );
  HS65_LH_AO222X4 U276 ( .A(n336), .B(n301), .C(n592), .D(n304), .E(n337), .F(
        n16), .Z(n290) );
  HS65_LH_MX41X7 U277 ( .D0(n523), .S0(n196), .D1(n522), .S1(n32), .D2(n521), 
        .S2(n26), .D3(n520), .S3(n20), .Z(n269) );
  HS65_LH_AO222X4 U278 ( .A(n324), .B(n301), .C(n304), .D(n216), .E(n325), .F(
        n17), .Z(n143) );
  HS65_LH_AO222X4 U279 ( .A(n299), .B(n301), .C(n247), .D(n304), .E(n119), .F(
        n16), .Z(n166) );
  HS65_LH_AO222X4 U280 ( .A(n334), .B(n7), .C(n222), .D(n304), .E(n335), .F(
        n17), .Z(n155) );
  HS65_LH_MX41X7 U281 ( .D0(n525), .S0(n196), .D1(n524), .S1(n31), .D2(n523), 
        .S2(n26), .D3(n522), .S3(n20), .Z(n226) );
  HS65_LH_MX41X7 U282 ( .D0(n526), .S0(n196), .D1(n525), .S1(n31), .D2(n524), 
        .S2(n26), .D3(n523), .S3(n20), .Z(n209) );
  HS65_LH_MX41X7 U283 ( .D0(n524), .S0(n36), .D1(n523), .S1(n31), .D2(n522), 
        .S2(n26), .D3(n521), .S3(n21), .Z(n251) );
  HS65_LH_OAI21X3 U284 ( .A(n77), .B(n97), .C(n123), .Z(n168) );
  HS65_LH_OAI21X3 U285 ( .A(n79), .B(n97), .C(n40), .Z(n147) );
  HS65_LH_OAI21X3 U286 ( .A(n85), .B(n54), .C(n40), .Z(n416) );
  HS65_LH_OAI21X3 U287 ( .A(n86), .B(n54), .C(n40), .Z(n410) );
  HS65_LH_OAI21X3 U288 ( .A(n88), .B(n54), .C(n40), .Z(n398) );
  HS65_LH_OAI21X3 U289 ( .A(n90), .B(n97), .C(n123), .Z(n382) );
  HS65_LH_OAI21X3 U290 ( .A(n517), .B(n97), .C(n123), .Z(n369) );
  HS65_LH_OAI21X3 U291 ( .A(n523), .B(n97), .C(n123), .Z(n319) );
  HS65_LH_OAI21X3 U292 ( .A(n524), .B(n97), .C(n123), .Z(n308) );
  HS65_LH_OAI21X3 U293 ( .A(n525), .B(n97), .C(n123), .Z(n294) );
  HS65_LH_OAI21X3 U294 ( .A(n520), .B(n55), .C(n123), .Z(n345) );
  HS65_LH_OAI21X3 U295 ( .A(n521), .B(n55), .C(n123), .Z(n339) );
  HS65_LH_OAI21X3 U296 ( .A(n522), .B(n55), .C(n123), .Z(n329) );
  HS65_LH_MX41X7 U297 ( .D0(n16), .S0(n306), .D1(n301), .S1(n305), .D2(n304), 
        .S2(n302), .D3(n374), .S3(n303), .Z(n252) );
  HS65_LH_MX41X7 U298 ( .D0(n16), .S0(n292), .D1(n7), .S1(n337), .D2(n304), 
        .S2(n336), .D3(n374), .S3(n592), .Z(n227) );
  HS65_LH_MX41X7 U299 ( .D0(n16), .S0(n278), .D1(n301), .S1(n327), .D2(n304), 
        .S2(n326), .D3(n374), .S3(n188), .Z(n210) );
  HS65_LH_OAI21X3 U300 ( .A(n81), .B(n97), .C(n40), .Z(n122) );
  HS65_LH_OAI21X3 U301 ( .A(n300), .B(n97), .C(n123), .Z(n376) );
  HS65_LH_IVX9 U302 ( .A(\alu_i[SRC_A][31] ), .Z(n562) );
  HS65_LH_AO22X9 U303 ( .A(n302), .B(n16), .C(n303), .D(n301), .Z(n165) );
  HS65_LH_AO22X9 U304 ( .A(n326), .B(n16), .C(n188), .D(n301), .Z(n141) );
  HS65_LH_AO22X9 U305 ( .A(n336), .B(n16), .C(n592), .D(n7), .Z(n153) );
  HS65_LH_IVX9 U306 ( .A(\alu_i[SRC_A][28] ), .Z(n566) );
  HS65_LH_AO22X9 U307 ( .A(n299), .B(n16), .C(n247), .D(n301), .Z(n116) );
  HS65_LH_AO22X9 U308 ( .A(n313), .B(n16), .C(n263), .D(n7), .Z(n131) );
  HS65_LH_AO22X9 U309 ( .A(n334), .B(n16), .C(n222), .D(n7), .Z(n291) );
  HS65_LH_OAI212X5 U310 ( .A(\alu_i[SRC_A][24] ), .B(n54), .C(n14), .D(n569), 
        .E(n41), .Z(n318) );
  HS65_LH_IVX9 U311 ( .A(\alu_i[SRC_A][24] ), .Z(n569) );
  HS65_LH_OAI212X5 U312 ( .A(\alu_i[SRC_A][21] ), .B(n55), .C(n15), .D(n573), 
        .E(n41), .Z(n344) );
  HS65_LH_IVX9 U313 ( .A(\alu_i[SRC_A][21] ), .Z(n573) );
  HS65_LH_IVX9 U314 ( .A(n190), .Z(n563) );
  HS65_LH_OAI212X5 U315 ( .A(\alu_i[SRC_A][18] ), .B(n55), .C(n15), .D(n576), 
        .E(n40), .Z(n375) );
  HS65_LH_IVX9 U316 ( .A(\alu_i[SRC_A][18] ), .Z(n576) );
  HS65_LH_IVX9 U317 ( .A(n264), .Z(n583) );
  HS65_LH_OAI212X5 U318 ( .A(\alu_i[SRC_A][6] ), .B(n54), .C(n14), .D(n588), 
        .E(n41), .Z(n158) );
  HS65_LH_IVX9 U319 ( .A(\alu_i[SRC_A][6] ), .Z(n588) );
  HS65_LH_OAI212X5 U320 ( .A(\alu_i[SRC_A][0] ), .B(n97), .C(n14), .D(n594), 
        .E(n441), .Z(n439) );
  HS65_LH_AOI12X2 U321 ( .A(n599), .B(n196), .C(n42), .Z(n441) );
  HS65_LH_OAI212X5 U322 ( .A(\alu_i[SRC_A][30] ), .B(n54), .C(n14), .D(n565), 
        .E(n41), .Z(n223) );
  HS65_LH_OAI212X5 U323 ( .A(\alu_i[SRC_A][1] ), .B(n55), .C(n15), .D(n593), 
        .E(n41), .Z(n357) );
  HS65_LH_CBI4I6X5 U324 ( .A(n531), .B(n54), .C(n40), .D(n565), .Z(n224) );
  HS65_LH_CBI4I6X5 U325 ( .A(n69), .B(n54), .C(n40), .D(n594), .Z(n440) );
  HS65_LH_CBI4I6X5 U326 ( .A(n70), .B(n54), .C(n40), .D(n593), .Z(n358) );
  HS65_LH_IVX9 U327 ( .A(\alu_i[SRC_A][30] ), .Z(n565) );
  HS65_LH_OAI21X3 U328 ( .A(n78), .B(n97), .C(n40), .Z(n159) );
  HS65_LH_OAI21X3 U329 ( .A(n80), .B(n54), .C(n40), .Z(n135) );
  HS65_LH_OAI21X3 U330 ( .A(n82), .B(n97), .C(n40), .Z(n429) );
  HS65_LH_OAI21X3 U331 ( .A(n87), .B(n54), .C(n40), .Z(n404) );
  HS65_LH_OAI21X3 U332 ( .A(n89), .B(n97), .C(n123), .Z(n389) );
  HS65_LH_IVX9 U333 ( .A(\alu_i[SRC_A][0] ), .Z(n594) );
  HS65_LH_IVX9 U334 ( .A(\alu_i[SRC_A][1] ), .Z(n593) );
  HS65_LH_IVX9 U335 ( .A(\alu_i[SRC_A][3] ), .Z(n590) );
  HS65_LH_NOR3X4 U336 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][4] ), .C(n607), .Z(
        n434) );
  HS65_LH_BFX9 U337 ( .A(n104), .Z(n46) );
  HS65_LH_OAI21X3 U338 ( .A(\alu_i[OP][0] ), .B(n437), .C(n443), .Z(n104) );
  HS65_LH_OAI21X3 U339 ( .A(n436), .B(n435), .C(n390), .Z(n443) );
  HS65_LH_NOR2X6 U340 ( .A(n596), .B(n96), .Z(n275) );
  HS65_LH_NAND2X7 U341 ( .A(n7), .B(n596), .Z(n189) );
  HS65_LH_NOR2X6 U342 ( .A(n602), .B(n601), .Z(n374) );
  HS65_LH_NOR2X6 U343 ( .A(n596), .B(n98), .Z(n117) );
  HS65_LH_NOR2X6 U344 ( .A(n609), .B(\alu_i[OP][1] ), .Z(n391) );
  HS65_LH_NOR2X6 U345 ( .A(\alu_i[OP][1] ), .B(\alu_i[OP][0] ), .Z(n438) );
  HS65_LH_NOR2X6 U346 ( .A(n611), .B(\alu_i[OP][0] ), .Z(n436) );
  HS65_LH_AND2X4 U347 ( .A(n192), .B(n606), .Z(n277) );
  HS65_LH_NAND2X7 U348 ( .A(n193), .B(n605), .Z(n208) );
  HS65_LH_NAND2X7 U349 ( .A(n193), .B(n606), .Z(n186) );
  HS65_LH_NAND4ABX3 U350 ( .A(\alu_i[OP][4] ), .B(\alu_i[OP][2] ), .C(n611), 
        .D(n607), .Z(n437) );
  HS65_LH_IVX9 U351 ( .A(\alu_i[OP][0] ), .Z(n609) );
  HS65_LH_NOR2AX3 U352 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][4] ), .Z(n445) );
  HS65_LH_IVX9 U353 ( .A(\alu_i[OP][4] ), .Z(n612) );
  HS65_LH_AND2X4 U354 ( .A(n448), .B(n602), .Z(n195) );
  HS65_LH_IVX9 U355 ( .A(\alu_i[OP][3] ), .Z(n607) );
  HS65_LH_IVX9 U356 ( .A(\alu_i[OP][1] ), .Z(n611) );
  HS65_LH_AND2X4 U357 ( .A(n192), .B(n605), .Z(n118) );
  HS65_LH_AND2X4 U358 ( .A(n445), .B(\alu_i[OP][3] ), .Z(n390) );
  HS65_LH_IVX9 U359 ( .A(n35), .Z(n38) );
  HS65_LH_IVX9 U360 ( .A(n6), .Z(n16) );
  HS65_LH_BFX9 U361 ( .A(n199), .Z(n18) );
  HS65_LH_BFX9 U362 ( .A(n197), .Z(n30) );
  HS65_LH_BFX9 U363 ( .A(n197), .Z(n29) );
  HS65_LH_BFX9 U364 ( .A(n25), .Z(n26) );
  HS65_LH_BFX9 U365 ( .A(n25), .Z(n28) );
  HS65_LH_BFX9 U366 ( .A(n25), .Z(n27) );
  HS65_LH_BFX9 U367 ( .A(n199), .Z(n19) );
  HS65_LH_IVX9 U368 ( .A(n6), .Z(n17) );
  HS65_LH_AO22X9 U369 ( .A(N226), .B(n61), .C(\HI_LO_c[HI][31] ), .D(n57), .Z(
        n516) );
  HS65_LH_IVX9 U370 ( .A(\alu_i[SRC_A][2] ), .Z(n535) );
  HS65_LH_IVX9 U371 ( .A(\alu_i[SRC_A][5] ), .Z(n537) );
  HS65_LH_IVX9 U372 ( .A(\alu_i[SRC_A][8] ), .Z(n539) );
  HS65_LH_IVX9 U373 ( .A(\alu_i[SRC_B][2] ), .Z(n72) );
  HS65_LH_BFX9 U374 ( .A(\alu_i[SRC_B][0] ), .Z(n69) );
  HS65_LH_AO22X9 U375 ( .A(N224), .B(n63), .C(\HI_LO_c[HI][29] ), .D(n57), .Z(
        n514) );
  HS65_LH_AO22X9 U376 ( .A(N225), .B(n62), .C(\HI_LO_c[HI][30] ), .D(n57), .Z(
        n515) );
  HS65_LH_IVX9 U377 ( .A(\alu_i[SRC_B][4] ), .Z(n76) );
  HS65_LH_IVX9 U378 ( .A(\alu_i[SRC_A][11] ), .Z(n541) );
  HS65_LH_IVX9 U379 ( .A(\alu_i[SRC_A][14] ), .Z(n543) );
  HS65_LH_IVX9 U380 ( .A(\alu_i[SRC_A][17] ), .Z(n545) );
  HS65_LH_IVX9 U381 ( .A(\alu_i[SRC_A][20] ), .Z(n547) );
  HS65_LH_IVX9 U382 ( .A(\alu_i[SRC_B][3] ), .Z(n74) );
  HS65_LH_AO22X9 U383 ( .A(N217), .B(n63), .C(\HI_LO_c[HI][22] ), .D(n57), .Z(
        n507) );
  HS65_LH_AO22X9 U384 ( .A(N218), .B(n63), .C(\HI_LO_c[HI][23] ), .D(n57), .Z(
        n508) );
  HS65_LH_AO22X9 U385 ( .A(N219), .B(n63), .C(\HI_LO_c[HI][24] ), .D(n57), .Z(
        n509) );
  HS65_LH_AO22X9 U386 ( .A(N220), .B(n63), .C(\HI_LO_c[HI][25] ), .D(n57), .Z(
        n510) );
  HS65_LH_AO22X9 U387 ( .A(N221), .B(n63), .C(\HI_LO_c[HI][26] ), .D(n57), .Z(
        n511) );
  HS65_LH_AO22X9 U388 ( .A(N222), .B(n63), .C(\HI_LO_c[HI][27] ), .D(n57), .Z(
        n512) );
  HS65_LH_AO22X9 U389 ( .A(N223), .B(n63), .C(\HI_LO_c[HI][28] ), .D(n57), .Z(
        n513) );
  HS65_LH_IVX9 U390 ( .A(\alu_i[SRC_B][11] ), .Z(n84) );
  HS65_LH_IVX9 U391 ( .A(\alu_i[SRC_A][23] ), .Z(n549) );
  HS65_LH_IVX9 U392 ( .A(\alu_i[SRC_A][26] ), .Z(n551) );
  HS65_LH_IVX9 U393 ( .A(\alu_i[SRC_A][29] ), .Z(n553) );
  HS65_LH_AO22X9 U394 ( .A(N210), .B(n63), .C(\HI_LO_c[HI][15] ), .D(n58), .Z(
        n500) );
  HS65_LH_AO22X9 U395 ( .A(N211), .B(n63), .C(\HI_LO_c[HI][16] ), .D(n58), .Z(
        n501) );
  HS65_LH_AO22X9 U396 ( .A(N212), .B(n63), .C(\HI_LO_c[HI][17] ), .D(n58), .Z(
        n502) );
  HS65_LH_AO22X9 U397 ( .A(N213), .B(n63), .C(\HI_LO_c[HI][18] ), .D(n58), .Z(
        n503) );
  HS65_LH_AO22X9 U398 ( .A(N214), .B(n63), .C(\HI_LO_c[HI][19] ), .D(n58), .Z(
        n504) );
  HS65_LH_AO22X9 U399 ( .A(N215), .B(n63), .C(\HI_LO_c[HI][20] ), .D(n57), .Z(
        n505) );
  HS65_LH_AO22X9 U400 ( .A(N216), .B(n63), .C(\HI_LO_c[HI][21] ), .D(n57), .Z(
        n506) );
  HS65_LH_IVX9 U401 ( .A(\alu_i[SRC_B][20] ), .Z(n519) );
  HS65_LH_AO22X9 U402 ( .A(N204), .B(n64), .C(\HI_LO_c[HI][9] ), .D(n58), .Z(
        n494) );
  HS65_LH_AO22X9 U403 ( .A(N205), .B(n63), .C(\HI_LO_c[HI][10] ), .D(n58), .Z(
        n495) );
  HS65_LH_AO22X9 U404 ( .A(N206), .B(n63), .C(\HI_LO_c[HI][11] ), .D(n58), .Z(
        n496) );
  HS65_LH_AO22X9 U405 ( .A(N207), .B(n63), .C(\HI_LO_c[HI][12] ), .D(n58), .Z(
        n497) );
  HS65_LH_AO22X9 U406 ( .A(N208), .B(n63), .C(\HI_LO_c[HI][13] ), .D(n58), .Z(
        n498) );
  HS65_LH_AO22X9 U407 ( .A(N209), .B(n63), .C(\HI_LO_c[HI][14] ), .D(n58), .Z(
        n499) );
  HS65_LH_IVX9 U408 ( .A(\alu_i[SRC_B][28] ), .Z(n529) );
  HS65_LH_IVX9 U409 ( .A(\alu_i[SRC_B][27] ), .Z(n527) );
  HS65_LH_AO22X9 U410 ( .A(N199), .B(n64), .C(\HI_LO_c[HI][4] ), .D(n58), .Z(
        n489) );
  HS65_LH_AO22X9 U411 ( .A(N200), .B(n64), .C(\HI_LO_c[HI][5] ), .D(n57), .Z(
        n490) );
  HS65_LH_AO22X9 U412 ( .A(N201), .B(n64), .C(\HI_LO_c[HI][6] ), .D(n58), .Z(
        n491) );
  HS65_LH_AO22X9 U413 ( .A(N202), .B(n64), .C(\HI_LO_c[HI][7] ), .D(n57), .Z(
        n492) );
  HS65_LH_AO22X9 U414 ( .A(N203), .B(n64), .C(\HI_LO_c[HI][8] ), .D(n58), .Z(
        n493) );
  HS65_LH_AO22X9 U415 ( .A(N197), .B(n64), .C(\HI_LO_c[HI][2] ), .D(n58), .Z(
        n487) );
  HS65_LH_AO22X9 U416 ( .A(N198), .B(n64), .C(\HI_LO_c[HI][3] ), .D(n57), .Z(
        n488) );
  HS65_LH_IVX9 U417 ( .A(\alu_i[SRC_B][31] ), .Z(n533) );
  HS65_LH_AO22X9 U418 ( .A(N194), .B(n64), .C(\HI_LO_c[LO][31] ), .D(n58), .Z(
        n484) );
  HS65_LH_AO22X9 U419 ( .A(N196), .B(n64), .C(\HI_LO_c[HI][1] ), .D(n57), .Z(
        n486) );
  HS65_LH_AO22X9 U420 ( .A(N191), .B(n64), .C(\HI_LO_c[LO][28] ), .D(n59), .Z(
        n481) );
  HS65_LH_AO22X9 U421 ( .A(N192), .B(n64), .C(\HI_LO_c[LO][29] ), .D(n58), .Z(
        n482) );
  HS65_LH_AO22X9 U422 ( .A(N193), .B(n64), .C(\HI_LO_c[LO][30] ), .D(n57), .Z(
        n483) );
  HS65_LH_AO22X9 U423 ( .A(N195), .B(n64), .C(\HI_LO_c[HI][0] ), .D(n60), .Z(
        n485) );
  HS65_LH_AO22X9 U424 ( .A(N184), .B(n65), .C(\HI_LO_c[LO][21] ), .D(n59), .Z(
        n474) );
  HS65_LH_AO22X9 U425 ( .A(N185), .B(n64), .C(\HI_LO_c[LO][22] ), .D(n59), .Z(
        n475) );
  HS65_LH_AO22X9 U426 ( .A(N186), .B(n64), .C(\HI_LO_c[LO][23] ), .D(n59), .Z(
        n476) );
  HS65_LH_AO22X9 U427 ( .A(N187), .B(n64), .C(\HI_LO_c[LO][24] ), .D(n59), .Z(
        n477) );
  HS65_LH_AO22X9 U428 ( .A(N188), .B(n64), .C(\HI_LO_c[LO][25] ), .D(n59), .Z(
        n478) );
  HS65_LH_AO22X9 U429 ( .A(N189), .B(n64), .C(\HI_LO_c[LO][26] ), .D(n59), .Z(
        n479) );
  HS65_LH_AO22X9 U430 ( .A(N190), .B(n64), .C(\HI_LO_c[LO][27] ), .D(n59), .Z(
        n480) );
  HS65_LH_AOI222X2 U431 ( .A(N157), .B(n51), .C(n11), .D(\HI_LO_c[HI][26] ), 
        .E(n8), .F(n526), .Z(n288) );
  HS65_LH_AOI222X2 U432 ( .A(N158), .B(n51), .C(n11), .D(\HI_LO_c[HI][27] ), 
        .E(n8), .F(n528), .Z(n273) );
  HS65_LH_AOI22X6 U433 ( .A(N128), .B(n48), .C(n606), .D(n250), .Z(n243) );
  HS65_LH_AO212X4 U434 ( .A(n251), .B(n595), .C(n252), .D(\alu_i[SHAMT][4] ), 
        .E(n253), .Z(n250) );
  HS65_LH_AO222X4 U435 ( .A(n192), .B(n254), .C(n193), .D(n255), .E(n195), .F(
        n256), .Z(n253) );
  HS65_LH_MX41X7 U436 ( .D0(n530), .S0(n196), .D1(n528), .S1(n31), .D2(n526), 
        .S2(n26), .D3(n525), .S3(n20), .Z(n255) );
  HS65_LH_AOI22X6 U437 ( .A(N129), .B(n48), .C(n606), .D(n225), .Z(n218) );
  HS65_LH_AO212X4 U438 ( .A(n226), .B(n595), .C(n227), .D(\alu_i[SHAMT][4] ), 
        .E(n228), .Z(n225) );
  HS65_LH_AO222X4 U439 ( .A(n192), .B(n229), .C(n193), .D(n230), .E(n195), .F(
        n231), .Z(n228) );
  HS65_LH_MX41X7 U440 ( .D0(n531), .S0(n36), .D1(n530), .S1(n31), .D2(n528), 
        .S2(n26), .D3(n526), .S3(n20), .Z(n230) );
  HS65_LH_MX41X7 U441 ( .D0(n45), .S0(\HI_LO_c[LO][25] ), .D1(n106), .S1(n81), 
        .D2(N124), .S2(n48), .D3(n599), .S3(n251), .Z(n295) );
  HS65_LH_MX41X7 U442 ( .D0(n45), .S0(\HI_LO_c[LO][26] ), .D1(n106), .S1(n82), 
        .D2(N125), .S2(n48), .D3(n599), .S3(n226), .Z(n286) );
  HS65_LH_MX41X7 U443 ( .D0(n45), .S0(\HI_LO_c[LO][27] ), .D1(n106), .S1(n83), 
        .D2(N126), .S2(n48), .D3(n599), .S3(n209), .Z(n271) );
  HS65_LH_AO22X9 U444 ( .A(N177), .B(n65), .C(\HI_LO_c[LO][14] ), .D(n60), .Z(
        n467) );
  HS65_LH_AO22X9 U445 ( .A(N178), .B(n65), .C(\HI_LO_c[LO][15] ), .D(n60), .Z(
        n468) );
  HS65_LH_AO22X9 U446 ( .A(N179), .B(n65), .C(\HI_LO_c[LO][16] ), .D(n59), .Z(
        n469) );
  HS65_LH_AO22X9 U447 ( .A(N180), .B(n65), .C(\HI_LO_c[LO][17] ), .D(n59), .Z(
        n470) );
  HS65_LH_AO22X9 U448 ( .A(N181), .B(n65), .C(\HI_LO_c[LO][18] ), .D(n59), .Z(
        n471) );
  HS65_LH_AO22X9 U449 ( .A(N182), .B(n65), .C(\HI_LO_c[LO][19] ), .D(n59), .Z(
        n472) );
  HS65_LH_AO22X9 U450 ( .A(N183), .B(n65), .C(\HI_LO_c[LO][20] ), .D(n59), .Z(
        n473) );
  HS65_LH_NAND4ABX3 U451 ( .A(n295), .B(n296), .C(n297), .D(n298), .Z(
        \alu_o[RESULT][25] ) );
  HS65_LH_MX41X7 U452 ( .D0(n277), .S0(n306), .D1(n598), .S1(n254), .D2(n524), 
        .S2(n307), .D3(\alu_i[SRC_A][25] ), .S3(n308), .Z(n296) );
  HS65_LH_AOI222X2 U453 ( .A(n275), .B(n112), .C(n279), .D(n256), .E(n284), 
        .F(n116), .Z(n298) );
  HS65_LH_NAND4ABX3 U454 ( .A(n286), .B(n287), .C(n288), .D(n289), .Z(
        \alu_o[RESULT][26] ) );
  HS65_LH_MX41X7 U455 ( .D0(n277), .S0(n292), .D1(n598), .S1(n229), .D2(n525), 
        .S2(n293), .D3(n550), .S3(n294), .Z(n287) );
  HS65_LH_AOI222X2 U456 ( .A(n275), .B(n290), .C(n279), .D(n231), .E(n284), 
        .F(n291), .Z(n289) );
  HS65_LH_NAND4ABX3 U457 ( .A(n271), .B(n272), .C(n273), .D(n274), .Z(
        \alu_o[RESULT][27] ) );
  HS65_LH_AOI222X2 U458 ( .A(n275), .B(n276), .C(n277), .D(n278), .E(n279), 
        .F(n214), .Z(n274) );
  HS65_LH_OAI212X5 U459 ( .A(n280), .B(n527), .C(n575), .D(n281), .E(n282), 
        .Z(n272) );
  HS65_LH_NAND3X5 U460 ( .A(n243), .B(n244), .C(n245), .Z(\alu_o[RESULT][29] )
         );
  HS65_LH_AOI212X4 U461 ( .A(n600), .B(n247), .C(n530), .D(n248), .E(n249), 
        .Z(n244) );
  HS65_LH_AOI212X4 U462 ( .A(n10), .B(n531), .C(N160), .D(n53), .E(n246), .Z(
        n245) );
  HS65_LH_NAND3X5 U463 ( .A(n218), .B(n219), .C(n220), .Z(\alu_o[RESULT][30] )
         );
  HS65_LH_AOI212X4 U464 ( .A(n600), .B(n222), .C(n531), .D(n223), .E(n224), 
        .Z(n219) );
  HS65_LH_AOI212X4 U465 ( .A(n10), .B(n532), .C(N161), .D(n53), .E(n221), .Z(
        n220) );
  HS65_LH_NAND2X7 U466 ( .A(n257), .B(n258), .Z(\alu_o[RESULT][28] ) );
  HS65_LH_AOI212X4 U467 ( .A(n9), .B(n530), .C(N159), .D(n53), .E(n270), .Z(
        n257) );
  HS65_LH_AOI212X4 U468 ( .A(N127), .B(n48), .C(n606), .D(n259), .E(n260), .Z(
        n258) );
  HS65_LH_NAND2X7 U469 ( .A(n201), .B(n202), .Z(\alu_o[RESULT][31] ) );
  HS65_LH_AOI212X4 U470 ( .A(n13), .B(\HI_LO_c[HI][31] ), .C(N162), .D(n53), 
        .E(n217), .Z(n201) );
  HS65_LH_AOI212X4 U471 ( .A(N130), .B(n48), .C(n606), .D(n203), .E(n204), .Z(
        n202) );
  HS65_LH_AOI222X2 U472 ( .A(N152), .B(n52), .C(n11), .D(\HI_LO_c[HI][21] ), 
        .E(n8), .F(n521), .Z(n342) );
  HS65_LH_AOI222X2 U473 ( .A(N153), .B(n51), .C(n11), .D(\HI_LO_c[HI][22] ), 
        .E(n8), .F(n522), .Z(n332) );
  HS65_LH_AOI222X2 U474 ( .A(N154), .B(n51), .C(n11), .D(\HI_LO_c[HI][23] ), 
        .E(n8), .F(n523), .Z(n322) );
  HS65_LH_AOI222X2 U475 ( .A(N155), .B(n51), .C(n11), .D(\HI_LO_c[HI][24] ), 
        .E(n8), .F(n524), .Z(n311) );
  HS65_LH_AOI222X2 U476 ( .A(N156), .B(n51), .C(n11), .D(\HI_LO_c[HI][25] ), 
        .E(n8), .F(n525), .Z(n297) );
  HS65_LH_AOI222X2 U477 ( .A(N149), .B(n52), .C(n12), .D(\HI_LO_c[HI][18] ), 
        .E(n9), .F(n517), .Z(n372) );
  HS65_LH_AOI222X2 U478 ( .A(N150), .B(n52), .C(n12), .D(\HI_LO_c[HI][19] ), 
        .E(n9), .F(n518), .Z(n365) );
  HS65_LH_AOI222X2 U479 ( .A(N151), .B(n52), .C(n12), .D(\HI_LO_c[HI][20] ), 
        .E(n9), .F(n520), .Z(n348) );
  HS65_LH_AOI212X4 U480 ( .A(n10), .B(n70), .C(N131), .D(n53), .E(n433), .Z(
        n432) );
  HS65_LH_AO222X4 U481 ( .A(N649), .B(n103), .C(n13), .D(\HI_LO_c[HI][0] ), 
        .E(N648), .F(n102), .Z(n433) );
  HS65_LH_MX41X7 U482 ( .D0(n45), .S0(\HI_LO_c[LO][17] ), .D1(n106), .S1(n70), 
        .D2(N116), .S2(n49), .D3(n599), .S3(n254), .Z(n377) );
  HS65_LH_MX41X7 U483 ( .D0(n45), .S0(\HI_LO_c[LO][18] ), .D1(n106), .S1(n71), 
        .D2(N117), .S2(n49), .D3(n599), .S3(n229), .Z(n370) );
  HS65_LH_MX41X7 U484 ( .D0(n45), .S0(\HI_LO_c[LO][19] ), .D1(n106), .S1(n73), 
        .D2(N118), .S2(n48), .D3(n599), .S3(n212), .Z(n363) );
  HS65_LH_MX41X7 U485 ( .D0(n45), .S0(\HI_LO_c[LO][20] ), .D1(n106), .S1(n75), 
        .D2(N119), .S2(n48), .D3(n599), .S3(n268), .Z(n346) );
  HS65_LH_MX41X7 U486 ( .D0(n45), .S0(\HI_LO_c[LO][21] ), .D1(n106), .S1(n77), 
        .D2(N120), .S2(n48), .D3(n599), .S3(n256), .Z(n340) );
  HS65_LH_MX41X7 U487 ( .D0(n45), .S0(\HI_LO_c[LO][22] ), .D1(n106), .S1(n78), 
        .D2(N121), .S2(n48), .D3(n599), .S3(n231), .Z(n330) );
  HS65_LH_MX41X7 U488 ( .D0(n45), .S0(\HI_LO_c[LO][23] ), .D1(n106), .S1(n79), 
        .D2(N122), .S2(n48), .D3(n599), .S3(n214), .Z(n320) );
  HS65_LH_MX41X7 U489 ( .D0(n45), .S0(\HI_LO_c[LO][24] ), .D1(n106), .S1(n80), 
        .D2(N123), .S2(n48), .D3(n599), .S3(n269), .Z(n309) );
  HS65_LH_AO22X9 U490 ( .A(N171), .B(n65), .C(\HI_LO_c[LO][8] ), .D(n60), .Z(
        n461) );
  HS65_LH_AO22X9 U491 ( .A(N172), .B(n65), .C(\HI_LO_c[LO][9] ), .D(n60), .Z(
        n462) );
  HS65_LH_AO22X9 U492 ( .A(N173), .B(n65), .C(\HI_LO_c[LO][10] ), .D(n60), .Z(
        n463) );
  HS65_LH_AO22X9 U493 ( .A(N174), .B(n65), .C(\HI_LO_c[LO][11] ), .D(n60), .Z(
        n464) );
  HS65_LH_AO22X9 U494 ( .A(N175), .B(n65), .C(\HI_LO_c[LO][12] ), .D(n60), .Z(
        n465) );
  HS65_LH_AO22X9 U495 ( .A(N176), .B(n65), .C(\HI_LO_c[LO][13] ), .D(n60), .Z(
        n466) );
  HS65_LH_NAND4ABX3 U496 ( .A(n340), .B(n341), .C(n342), .D(n343), .Z(
        \alu_o[RESULT][21] ) );
  HS65_LH_MX41X7 U497 ( .D0(n277), .S0(n305), .D1(n598), .S1(n306), .D2(n520), 
        .S2(n344), .D3(\alu_i[SRC_A][21] ), .S3(n345), .Z(n341) );
  HS65_LH_AOI222X2 U498 ( .A(n275), .B(n165), .C(n279), .D(n254), .E(n284), 
        .F(n166), .Z(n343) );
  HS65_LH_NAND4ABX3 U499 ( .A(n330), .B(n331), .C(n332), .D(n333), .Z(
        \alu_o[RESULT][22] ) );
  HS65_LH_MX41X7 U500 ( .D0(n277), .S0(n337), .D1(n598), .S1(n292), .D2(n521), 
        .S2(n338), .D3(\alu_i[SRC_A][22] ), .S3(n339), .Z(n331) );
  HS65_LH_AOI222X2 U501 ( .A(n275), .B(n153), .C(n279), .D(n229), .E(n284), 
        .F(n155), .Z(n333) );
  HS65_LH_NAND4ABX3 U502 ( .A(n320), .B(n321), .C(n322), .D(n323), .Z(
        \alu_o[RESULT][23] ) );
  HS65_LH_MX41X7 U503 ( .D0(n277), .S0(n327), .D1(n598), .S1(n278), .D2(n522), 
        .S2(n328), .D3(n548), .S3(n329), .Z(n321) );
  HS65_LH_AOI222X2 U504 ( .A(n275), .B(n141), .C(n279), .D(n212), .E(n284), 
        .F(n143), .Z(n323) );
  HS65_LH_NAND4ABX3 U505 ( .A(n309), .B(n310), .C(n311), .D(n312), .Z(
        \alu_o[RESULT][24] ) );
  HS65_LH_MX41X7 U506 ( .D0(n277), .S0(n317), .D1(n598), .S1(n266), .D2(n523), 
        .S2(n318), .D3(\alu_i[SRC_A][24] ), .S3(n319), .Z(n310) );
  HS65_LH_AOI222X2 U507 ( .A(n275), .B(n129), .C(n279), .D(n268), .E(n284), 
        .F(n131), .Z(n312) );
  HS65_LH_NAND4ABX3 U508 ( .A(n377), .B(n378), .C(n379), .D(n380), .Z(
        \alu_o[RESULT][17] ) );
  HS65_LH_MX41X7 U509 ( .D0(n598), .S0(n305), .D1(n90), .S1(n381), .D2(n368), 
        .S2(n303), .D3(n544), .S3(n382), .Z(n378) );
  HS65_LH_AOI222X2 U510 ( .A(n284), .B(n360), .C(n277), .D(n302), .E(n279), 
        .F(n306), .Z(n380) );
  HS65_LH_NAND4ABX3 U511 ( .A(n370), .B(n371), .C(n372), .D(n373), .Z(
        \alu_o[RESULT][18] ) );
  HS65_LH_MX41X7 U512 ( .D0(n598), .S0(n337), .D1(n300), .S1(n375), .D2(n368), 
        .S2(n592), .D3(\alu_i[SRC_A][18] ), .S3(n376), .Z(n371) );
  HS65_LH_AOI222X2 U513 ( .A(n284), .B(n239), .C(n277), .D(n336), .E(n279), 
        .F(n292), .Z(n373) );
  HS65_LH_NAND4ABX3 U514 ( .A(n363), .B(n364), .C(n365), .D(n366), .Z(
        \alu_o[RESULT][19] ) );
  HS65_LH_MX41X7 U515 ( .D0(n598), .S0(n327), .D1(n517), .S1(n367), .D2(n368), 
        .S2(n188), .D3(\alu_i[SRC_A][19] ), .S3(n369), .Z(n364) );
  HS65_LH_AOI222X2 U516 ( .A(n284), .B(n563), .C(n277), .D(n326), .E(n279), 
        .F(n278), .Z(n366) );
  HS65_LH_NAND4ABX3 U517 ( .A(n346), .B(n347), .C(n348), .D(n349), .Z(
        \alu_o[RESULT][20] ) );
  HS65_LH_AOI222X2 U518 ( .A(n284), .B(n174), .C(n277), .D(n316), .E(n279), 
        .F(n266), .Z(n349) );
  HS65_LH_OAI212X5 U519 ( .A(n350), .B(n519), .C(n582), .D(n281), .E(n351), 
        .Z(n347) );
  HS65_LH_NAND3X5 U520 ( .A(n430), .B(n431), .C(n432), .Z(\alu_o[RESULT][0] )
         );
  HS65_LH_AOI212X4 U521 ( .A(N99), .B(n48), .C(n69), .D(n439), .E(n440), .Z(
        n431) );
  HS65_LH_AOI22X6 U522 ( .A(n605), .B(n444), .C(n45), .D(\HI_LO_c[LO][0] ), 
        .Z(n430) );
  HS65_LH_AOI222X2 U523 ( .A(n44), .B(\HI_LO_c[LO][9] ), .C(n600), .D(n111), 
        .E(N108), .F(n47), .Z(n110) );
  HS65_LH_AOI222X2 U524 ( .A(n44), .B(\HI_LO_c[LO][10] ), .C(n600), .D(n154), 
        .E(N109), .F(n47), .Z(n427) );
  HS65_LH_AOI222X2 U525 ( .A(n44), .B(\HI_LO_c[LO][11] ), .C(n600), .D(n142), 
        .E(N110), .F(n47), .Z(n420) );
  HS65_LH_AOI222X2 U526 ( .A(n44), .B(\HI_LO_c[LO][12] ), .C(n600), .D(n130), 
        .E(N111), .F(n47), .Z(n414) );
  HS65_LH_AOI222X2 U527 ( .A(n44), .B(\HI_LO_c[LO][13] ), .C(n600), .D(n114), 
        .E(N112), .F(n47), .Z(n408) );
  HS65_LH_AOI222X2 U528 ( .A(n44), .B(\HI_LO_c[LO][14] ), .C(n600), .D(n157), 
        .E(N113), .F(n47), .Z(n402) );
  HS65_LH_AOI222X2 U529 ( .A(n44), .B(\HI_LO_c[LO][15] ), .C(n600), .D(n145), 
        .E(N114), .F(n47), .Z(n395) );
  HS65_LH_AOI222X2 U530 ( .A(N140), .B(n51), .C(n11), .D(\HI_LO_c[HI][9] ), 
        .E(n8), .F(n82), .Z(n109) );
  HS65_LH_AOI222X2 U531 ( .A(N141), .B(n52), .C(n12), .D(\HI_LO_c[HI][10] ), 
        .E(n9), .F(n83), .Z(n426) );
  HS65_LH_AOI222X2 U532 ( .A(N142), .B(n52), .C(n12), .D(\HI_LO_c[HI][11] ), 
        .E(n9), .F(n85), .Z(n419) );
  HS65_LH_AOI222X2 U533 ( .A(N143), .B(n52), .C(n12), .D(\HI_LO_c[HI][12] ), 
        .E(n9), .F(n86), .Z(n413) );
  HS65_LH_AOI222X2 U534 ( .A(N144), .B(n52), .C(n12), .D(\HI_LO_c[HI][13] ), 
        .E(n9), .F(n87), .Z(n407) );
  HS65_LH_AOI222X2 U535 ( .A(N145), .B(n52), .C(n12), .D(\HI_LO_c[HI][14] ), 
        .E(n9), .F(n88), .Z(n401) );
  HS65_LH_AOI222X2 U536 ( .A(N146), .B(n52), .C(n12), .D(\HI_LO_c[HI][15] ), 
        .E(n9), .F(n89), .Z(n394) );
  HS65_LH_AOI222X2 U537 ( .A(N147), .B(n52), .C(n12), .D(\HI_LO_c[HI][16] ), 
        .E(n9), .F(n90), .Z(n385) );
  HS65_LH_AOI222X2 U538 ( .A(N148), .B(n52), .C(n12), .D(\HI_LO_c[HI][17] ), 
        .E(n9), .F(n300), .Z(n379) );
  HS65_LH_MX41X7 U539 ( .D0(n45), .S0(\HI_LO_c[LO][16] ), .D1(n106), .S1(n69), 
        .D2(N115), .S2(n49), .D3(n599), .S3(n266), .Z(n383) );
  HS65_LH_AO22X9 U540 ( .A(N167), .B(n65), .C(\HI_LO_c[LO][4] ), .D(n60), .Z(
        n457) );
  HS65_LH_AO22X9 U541 ( .A(N168), .B(n65), .C(\HI_LO_c[LO][5] ), .D(n60), .Z(
        n458) );
  HS65_LH_AO22X9 U542 ( .A(N169), .B(n65), .C(\HI_LO_c[LO][6] ), .D(n60), .Z(
        n459) );
  HS65_LH_AO22X9 U543 ( .A(N170), .B(n65), .C(\HI_LO_c[LO][7] ), .D(n60), .Z(
        n460) );
  HS65_LH_AO22X9 U544 ( .A(N163), .B(n66), .C(\HI_LO_c[LO][0] ), .D(n60), .Z(
        n453) );
  HS65_LH_AO22X9 U545 ( .A(N164), .B(n66), .C(\HI_LO_c[LO][1] ), .D(n59), .Z(
        n454) );
  HS65_LH_AO22X9 U546 ( .A(N165), .B(n65), .C(\HI_LO_c[LO][2] ), .D(n60), .Z(
        n455) );
  HS65_LH_AO22X9 U547 ( .A(N166), .B(n65), .C(\HI_LO_c[LO][3] ), .D(n59), .Z(
        n456) );
  HS65_LH_NAND4ABX3 U548 ( .A(n383), .B(n384), .C(n385), .D(n386), .Z(
        \alu_o[RESULT][16] ) );
  HS65_LH_MX41X7 U549 ( .D0(n598), .S0(n316), .D1(n89), .S1(n388), .D2(n368), 
        .S2(n315), .D3(\alu_i[SRC_A][16] ), .S3(n389), .Z(n384) );
  HS65_LH_AOI222X2 U550 ( .A(n284), .B(n387), .C(n277), .D(n314), .E(n279), 
        .F(n317), .Z(n386) );
  HS65_LH_NAND4ABX3 U551 ( .A(n107), .B(n108), .C(n109), .D(n110), .Z(
        \alu_o[RESULT][9] ) );
  HS65_LH_MX41X7 U552 ( .D0(n118), .S0(n119), .D1(n597), .S1(n120), .D2(n81), 
        .S2(n121), .D3(\alu_i[SRC_A][9] ), .S3(n122), .Z(n107) );
  HS65_LH_AO222X4 U553 ( .A(n112), .B(n113), .C(n114), .D(n115), .E(n116), .F(
        n117), .Z(n108) );
  HS65_LH_NAND4ABX3 U554 ( .A(n424), .B(n425), .C(n426), .D(n427), .Z(
        \alu_o[RESULT][10] ) );
  HS65_LH_MX41X7 U555 ( .D0(n118), .S0(n335), .D1(n597), .S1(n156), .D2(n82), 
        .S2(n428), .D3(\alu_i[SRC_A][10] ), .S3(n429), .Z(n424) );
  HS65_LH_AO222X4 U556 ( .A(n290), .B(n113), .C(n157), .D(n115), .E(n291), .F(
        n117), .Z(n425) );
  HS65_LH_NAND4ABX3 U557 ( .A(n417), .B(n418), .C(n419), .D(n420), .Z(
        \alu_o[RESULT][11] ) );
  HS65_LH_OAI212X5 U558 ( .A(n421), .B(n84), .C(n572), .D(n176), .E(n422), .Z(
        n417) );
  HS65_LH_AO222X4 U559 ( .A(n145), .B(n115), .C(n325), .D(n118), .E(n276), .F(
        n113), .Z(n418) );
  HS65_LH_NAND4ABX3 U560 ( .A(n411), .B(n412), .C(n413), .D(n414), .Z(
        \alu_o[RESULT][12] ) );
  HS65_LH_MX41X7 U561 ( .D0(n597), .S0(n132), .D1(n85), .S1(n415), .D2(n397), 
        .S2(n263), .D3(\alu_i[SRC_A][12] ), .S3(n416), .Z(n411) );
  HS65_LH_AO222X4 U562 ( .A(n133), .B(n115), .C(n313), .D(n118), .E(n583), .F(
        n113), .Z(n412) );
  HS65_LH_NAND4ABX3 U563 ( .A(n405), .B(n406), .C(n407), .D(n408), .Z(
        \alu_o[RESULT][13] ) );
  HS65_LH_MX41X7 U564 ( .D0(n597), .S0(n119), .D1(n86), .S1(n409), .D2(n397), 
        .S2(n247), .D3(\alu_i[SRC_A][13] ), .S3(n410), .Z(n405) );
  HS65_LH_AO222X4 U565 ( .A(n120), .B(n115), .C(n299), .D(n118), .E(n252), .F(
        n113), .Z(n406) );
  HS65_LH_NAND4ABX3 U566 ( .A(n399), .B(n400), .C(n401), .D(n402), .Z(
        \alu_o[RESULT][14] ) );
  HS65_LH_MX41X7 U567 ( .D0(n597), .S0(n335), .D1(n87), .S1(n403), .D2(n397), 
        .S2(n222), .D3(n542), .S3(n404), .Z(n399) );
  HS65_LH_AO222X4 U568 ( .A(n156), .B(n115), .C(n334), .D(n118), .E(n227), .F(
        n113), .Z(n400) );
  HS65_LH_NAND4ABX3 U569 ( .A(n392), .B(n393), .C(n394), .D(n395), .Z(
        \alu_o[RESULT][15] ) );
  HS65_LH_MX41X7 U570 ( .D0(n597), .S0(n325), .D1(n88), .S1(n396), .D2(n397), 
        .S2(n216), .D3(\alu_i[SRC_A][15] ), .S3(n398), .Z(n392) );
  HS65_LH_AO222X4 U571 ( .A(n144), .B(n115), .C(n324), .D(n118), .E(n210), .F(
        n113), .Z(n393) );
  HS65_LH_AOI222X2 U572 ( .A(n317), .B(n16), .C(n316), .D(n301), .E(n178), .F(
        \alu_i[SHAMT][3] ), .Z(n264) );
  HS65_LH_AOI222X2 U573 ( .A(n144), .B(n16), .C(n325), .D(n7), .E(n283), .F(
        \alu_i[SHAMT][3] ), .Z(n190) );
  HS65_LH_AOI222X2 U574 ( .A(n44), .B(\HI_LO_c[LO][5] ), .C(n600), .D(n164), 
        .E(N104), .F(n47), .Z(n163) );
  HS65_LH_AOI222X2 U575 ( .A(n44), .B(\HI_LO_c[LO][6] ), .C(n600), .D(n152), 
        .E(N105), .F(n47), .Z(n151) );
  HS65_LH_AOI222X2 U576 ( .A(n44), .B(\HI_LO_c[LO][7] ), .C(n600), .D(n140), 
        .E(N106), .F(n47), .Z(n139) );
  HS65_LH_AOI222X2 U577 ( .A(n44), .B(\HI_LO_c[LO][8] ), .C(n600), .D(n128), 
        .E(N107), .F(n47), .Z(n127) );
  HS65_LH_AOI222X2 U578 ( .A(N135), .B(n51), .C(n11), .D(\HI_LO_c[HI][4] ), 
        .E(n8), .F(n77), .Z(n171) );
  HS65_LH_AOI222X2 U579 ( .A(N136), .B(n51), .C(n12), .D(\HI_LO_c[HI][5] ), 
        .E(n8), .F(n78), .Z(n162) );
  HS65_LH_AOI222X2 U580 ( .A(N137), .B(n51), .C(n11), .D(\HI_LO_c[HI][6] ), 
        .E(n8), .F(n79), .Z(n150) );
  HS65_LH_AOI222X2 U581 ( .A(N138), .B(n51), .C(n11), .D(\HI_LO_c[HI][7] ), 
        .E(n8), .F(n80), .Z(n138) );
  HS65_LH_AOI222X2 U582 ( .A(N139), .B(n51), .C(n11), .D(\HI_LO_c[HI][8] ), 
        .E(n8), .F(n81), .Z(n126) );
  HS65_LH_AOI22X6 U583 ( .A(N100), .B(n48), .C(n605), .D(n359), .Z(n353) );
  HS65_LH_AO212X4 U584 ( .A(n164), .B(n595), .C(n360), .D(\alu_i[SHAMT][4] ), 
        .E(n361), .Z(n359) );
  HS65_LH_AO222X4 U585 ( .A(n192), .B(n114), .C(n193), .D(n362), .E(n195), .F(
        n111), .Z(n361) );
  HS65_LH_MX41X7 U586 ( .D0(n70), .S0(n36), .D1(n71), .S1(n32), .D2(n73), .S2(
        n27), .D3(n75), .S3(n21), .Z(n362) );
  HS65_LH_AO22X9 U587 ( .A(n602), .B(n314), .C(\alu_i[SHAMT][2] ), .D(n315), 
        .Z(n178) );
  HS65_LH_AO22X9 U588 ( .A(n602), .B(n324), .C(\alu_i[SHAMT][2] ), .D(n216), 
        .Z(n283) );
  HS65_LH_NAND3X5 U589 ( .A(n353), .B(n354), .C(n355), .Z(\alu_o[RESULT][1] )
         );
  HS65_LH_AOI212X4 U590 ( .A(n599), .B(n303), .C(n70), .D(n357), .E(n358), .Z(
        n354) );
  HS65_LH_AOI212X4 U591 ( .A(n9), .B(n71), .C(N132), .D(n53), .E(n356), .Z(
        n355) );
  HS65_LH_AO212X4 U592 ( .A(n152), .B(n595), .C(n239), .D(\alu_i[SHAMT][4] ), 
        .E(n240), .Z(n234) );
  HS65_LH_AO222X4 U593 ( .A(n192), .B(n157), .C(n193), .D(n241), .E(n195), .F(
        n154), .Z(n240) );
  HS65_LH_MX41X7 U594 ( .D0(n71), .S0(n196), .D1(n73), .S1(n31), .D2(n75), 
        .S2(n26), .D3(n77), .S3(n20), .Z(n241) );
  HS65_LH_AO222X4 U595 ( .A(\HI_LO_c[LO][28] ), .B(n45), .C(n85), .D(n106), 
        .E(\HI_LO_c[HI][28] ), .F(n13), .Z(n270) );
  HS65_LH_AO222X4 U596 ( .A(\HI_LO_c[LO][29] ), .B(n45), .C(n86), .D(n106), 
        .E(\HI_LO_c[HI][29] ), .F(n13), .Z(n246) );
  HS65_LH_AO222X4 U597 ( .A(\HI_LO_c[LO][30] ), .B(n44), .C(n87), .D(n106), 
        .E(\HI_LO_c[HI][30] ), .F(n13), .Z(n221) );
  HS65_LH_AO212X4 U598 ( .A(n173), .B(n595), .C(n387), .D(\alu_i[SHAMT][4] ), 
        .E(n446), .Z(n444) );
  HS65_LH_AO222X4 U599 ( .A(n192), .B(n130), .C(n193), .D(n447), .E(n195), .F(
        n128), .Z(n446) );
  HS65_LH_AO212X4 U600 ( .A(n26), .B(n71), .C(n34), .D(n70), .E(n449), .Z(n447) );
  HS65_LH_AO12X9 U601 ( .A(n73), .B(n20), .C(n315), .Z(n449) );
  HS65_LH_AO22X9 U602 ( .A(\HI_LO_c[LO][31] ), .B(n45), .C(n88), .D(n106), .Z(
        n217) );
  HS65_LH_AO212X4 U603 ( .A(n209), .B(n595), .C(n210), .D(\alu_i[SHAMT][4] ), 
        .E(n211), .Z(n203) );
  HS65_LH_AO222X4 U604 ( .A(n192), .B(n212), .C(n193), .D(n213), .E(n195), .F(
        n214), .Z(n211) );
  HS65_LH_AO212X4 U605 ( .A(n26), .B(n530), .C(n34), .D(n531), .E(n215), .Z(
        n213) );
  HS65_LH_AO12X9 U606 ( .A(n528), .B(n20), .C(n216), .Z(n215) );
  HS65_LH_NAND4ABX3 U607 ( .A(n169), .B(n170), .C(n171), .D(n172), .Z(
        \alu_o[RESULT][4] ) );
  HS65_LH_OAI212X5 U608 ( .A(n175), .B(n76), .C(n579), .D(n176), .E(n177), .Z(
        n169) );
  HS65_LH_AOI222X2 U609 ( .A(n44), .B(\HI_LO_c[LO][4] ), .C(n600), .D(n173), 
        .E(N103), .F(n47), .Z(n172) );
  HS65_LH_NAND4ABX3 U610 ( .A(n160), .B(n161), .C(n162), .D(n163), .Z(
        \alu_o[RESULT][5] ) );
  HS65_LH_MX41X7 U611 ( .D0(n118), .S0(n120), .D1(n597), .S1(n114), .D2(n77), 
        .S2(n167), .D3(n536), .S3(n168), .Z(n160) );
  HS65_LH_AO222X4 U612 ( .A(n165), .B(n113), .C(n111), .D(n115), .E(n166), .F(
        n117), .Z(n161) );
  HS65_LH_NAND4ABX3 U613 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(
        \alu_o[RESULT][6] ) );
  HS65_LH_MX41X7 U614 ( .D0(n118), .S0(n156), .D1(n597), .S1(n157), .D2(n78), 
        .S2(n158), .D3(\alu_i[SRC_A][6] ), .S3(n159), .Z(n148) );
  HS65_LH_AO222X4 U615 ( .A(n153), .B(n113), .C(n154), .D(n115), .E(n155), .F(
        n117), .Z(n149) );
  HS65_LH_NAND4ABX3 U616 ( .A(n136), .B(n137), .C(n138), .D(n139), .Z(
        \alu_o[RESULT][7] ) );
  HS65_LH_MX41X7 U617 ( .D0(n118), .S0(n144), .D1(n597), .S1(n145), .D2(n79), 
        .S2(n146), .D3(\alu_i[SRC_A][7] ), .S3(n147), .Z(n136) );
  HS65_LH_AO222X4 U618 ( .A(n141), .B(n113), .C(n142), .D(n115), .E(n143), .F(
        n117), .Z(n137) );
  HS65_LH_NAND4ABX3 U619 ( .A(n124), .B(n125), .C(n126), .D(n127), .Z(
        \alu_o[RESULT][8] ) );
  HS65_LH_MX41X7 U620 ( .D0(n118), .S0(n132), .D1(n597), .S1(n133), .D2(n80), 
        .S2(n134), .D3(n538), .S3(n135), .Z(n124) );
  HS65_LH_AO222X4 U621 ( .A(n129), .B(n113), .C(n130), .D(n115), .E(n131), .F(
        n117), .Z(n125) );
  HS65_LH_NAND2X7 U622 ( .A(n232), .B(n233), .Z(\alu_o[RESULT][2] ) );
  HS65_LH_AOI212X4 U623 ( .A(n10), .B(n73), .C(N133), .D(n53), .E(n242), .Z(
        n232) );
  HS65_LH_AOI212X4 U624 ( .A(N101), .B(n48), .C(n605), .D(n234), .E(n235), .Z(
        n233) );
  HS65_LH_NAND2X7 U625 ( .A(n181), .B(n182), .Z(\alu_o[RESULT][3] ) );
  HS65_LH_AOI212X4 U626 ( .A(n10), .B(n75), .C(N134), .D(n53), .E(n200), .Z(
        n181) );
  HS65_LH_AOI212X4 U627 ( .A(N102), .B(n48), .C(n605), .D(n183), .E(n184), .Z(
        n182) );
  HS65_LH_OR2X9 U628 ( .A(\alu_i[SHAMT][2] ), .B(\alu_i[SHAMT][3] ), .Z(n6) );
  HS65_LH_NOR2X6 U629 ( .A(n602), .B(\alu_i[SHAMT][3] ), .Z(n301) );
  HS65_LH_NOR2X6 U630 ( .A(n602), .B(\alu_i[SHAMT][3] ), .Z(n7) );
  HS65_LH_IVX9 U631 ( .A(\alu_i[SHAMT][4] ), .Z(n596) );
  HS65_LH_AND2X4 U632 ( .A(\alu_i[SHAMT][1] ), .B(\alu_i[SHAMT][0] ), .Z(n199)
         );
  HS65_LH_NOR2X6 U633 ( .A(n6), .B(\alu_i[SHAMT][4] ), .Z(n193) );
  HS65_LH_NOR2X6 U634 ( .A(n601), .B(\alu_i[SHAMT][2] ), .Z(n304) );
  HS65_LH_NOR2X6 U635 ( .A(n96), .B(\alu_i[SHAMT][4] ), .Z(n113) );
  HS65_LH_NOR2AX3 U636 ( .A(\alu_i[SHAMT][0] ), .B(\alu_i[SHAMT][1] ), .Z(n197) );
  HS65_LH_IVX9 U637 ( .A(\alu_i[SHAMT][3] ), .Z(n601) );
  HS65_LH_NOR2X6 U638 ( .A(n601), .B(\alu_i[SHAMT][4] ), .Z(n448) );
  HS65_LH_IVX9 U639 ( .A(\alu_i[SHAMT][2] ), .Z(n602) );
  HS65_LH_AND2X4 U640 ( .A(n448), .B(\alu_i[SHAMT][2] ), .Z(n192) );
  HS65_LH_BFX9 U641 ( .A(n196), .Z(n35) );
  HS65_LH_NOR2X6 U642 ( .A(\alu_i[SHAMT][0] ), .B(\alu_i[SHAMT][1] ), .Z(n196)
         );
  HS65_LH_BFX9 U643 ( .A(n198), .Z(n25) );
  HS65_LH_NOR2AX3 U644 ( .A(\alu_i[SHAMT][1] ), .B(\alu_i[SHAMT][0] ), .Z(n198) );
  HS65_LH_AO22X9 U645 ( .A(\HI_LO_c[HI][1] ), .B(n13), .C(\HI_LO_c[LO][1] ), 
        .D(n45), .Z(n356) );
  HS65_LH_AO22X9 U646 ( .A(\HI_LO_c[HI][2] ), .B(n13), .C(\HI_LO_c[LO][2] ), 
        .D(n45), .Z(n242) );
  HS65_LH_AO22X9 U647 ( .A(\HI_LO_c[HI][3] ), .B(n13), .C(\HI_LO_c[LO][3] ), 
        .D(n45), .Z(n200) );
endmodule


module alu_ctrl ( .alu_ctrl_i({\alu_ctrl_i[OP][3] , \alu_ctrl_i[OP][2] , 
        \alu_ctrl_i[OP][1] , \alu_ctrl_i[OP][0] , \alu_ctrl_i[FUNCT][5] , 
        \alu_ctrl_i[FUNCT][4] , \alu_ctrl_i[FUNCT][3] , \alu_ctrl_i[FUNCT][2] , 
        \alu_ctrl_i[FUNCT][1] , \alu_ctrl_i[FUNCT][0] }), .alu_ctrl_o({
        \alu_ctrl_o[OP][4] , \alu_ctrl_o[OP][3] , \alu_ctrl_o[OP][2] , 
        \alu_ctrl_o[OP][1] , \alu_ctrl_o[OP][0] , \alu_ctrl_o[BRANCH_SRC][1] , 
        \alu_ctrl_o[BRANCH_SRC][0] }) );
  input \alu_ctrl_i[OP][3] , \alu_ctrl_i[OP][2] , \alu_ctrl_i[OP][1] ,
         \alu_ctrl_i[OP][0] , \alu_ctrl_i[FUNCT][5] , \alu_ctrl_i[FUNCT][4] ,
         \alu_ctrl_i[FUNCT][3] , \alu_ctrl_i[FUNCT][2] ,
         \alu_ctrl_i[FUNCT][1] , \alu_ctrl_i[FUNCT][0] ;
  output \alu_ctrl_o[OP][4] , \alu_ctrl_o[OP][3] , \alu_ctrl_o[OP][2] ,
         \alu_ctrl_o[OP][1] , \alu_ctrl_o[OP][0] , \alu_ctrl_o[BRANCH_SRC][1] ,
         \alu_ctrl_o[BRANCH_SRC][0] ;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17;

  HS65_LH_AOI12X2 U3 ( .A(n38), .B(n39), .C(\alu_ctrl_i[OP][3] ), .Z(
        \alu_ctrl_o[OP][0] ) );
  HS65_LH_OAI32X5 U4 ( .A(n41), .B(\alu_ctrl_i[OP][3] ), .C(
        \alu_ctrl_i[OP][1] ), .D(n17), .E(n28), .Z(\alu_ctrl_o[BRANCH_SRC][1] ) );
  HS65_LH_IVX9 U5 ( .A(n30), .Z(n13) );
  HS65_LH_NAND3X5 U6 ( .A(n16), .B(n14), .C(n17), .Z(n30) );
  HS65_LH_AO312X9 U7 ( .A(n11), .B(n7), .C(n1), .D(n25), .E(n12), .F(n23), .Z(
        \alu_ctrl_o[OP][2] ) );
  HS65_LH_OAI33X3 U8 ( .A(n29), .B(n9), .C(n30), .D(n14), .E(n17), .F(n16), 
        .Z(n25) );
  HS65_LH_IVX9 U9 ( .A(n31), .Z(n9) );
  HS65_LH_NAND2X7 U10 ( .A(n13), .B(n12), .Z(n20) );
  HS65_LH_IVX9 U11 ( .A(n35), .Z(n5) );
  HS65_LH_IVX9 U12 ( .A(n27), .Z(n1) );
  HS65_LH_IVX9 U13 ( .A(n41), .Z(n15) );
  HS65_LH_NOR2AX3 U14 ( .A(n19), .B(n20), .Z(\alu_ctrl_o[BRANCH_SRC][0] ) );
  HS65_LH_AOI311X4 U15 ( .A(\alu_ctrl_i[FUNCT][0] ), .B(n8), .C(n40), .D(n3), 
        .E(n15), .Z(n39) );
  HS65_LH_AOI12X2 U16 ( .A(\alu_ctrl_i[OP][1] ), .B(n17), .C(n44), .Z(n38) );
  HS65_LH_IVX9 U17 ( .A(n33), .Z(n3) );
  HS65_LH_OAI32X5 U18 ( .A(n26), .B(n7), .C(n27), .D(\alu_ctrl_i[OP][0] ), .E(
        n28), .Z(n23) );
  HS65_LH_NAND2X7 U19 ( .A(\alu_ctrl_i[FUNCT][1] ), .B(n11), .Z(n26) );
  HS65_LH_OAI211X5 U20 ( .A(n20), .B(n4), .C(n2), .D(n21), .Z(
        \alu_ctrl_o[OP][3] ) );
  HS65_LH_IVX9 U21 ( .A(n24), .Z(n4) );
  HS65_LH_AOI32X5 U22 ( .A(n1), .B(\alu_ctrl_i[FUNCT][0] ), .C(n22), .D(n5), 
        .E(n12), .Z(n21) );
  HS65_LH_IVX9 U23 ( .A(n23), .Z(n2) );
  HS65_LH_NOR3AX2 U24 ( .A(n45), .B(n30), .C(n6), .Z(n40) );
  HS65_LH_NOR3X4 U25 ( .A(n10), .B(\alu_ctrl_i[FUNCT][4] ), .C(
        \alu_ctrl_i[FUNCT][2] ), .Z(n45) );
  HS65_LH_IVX9 U26 ( .A(\alu_ctrl_i[FUNCT][0] ), .Z(n11) );
  HS65_LH_AOI32X5 U27 ( .A(\alu_ctrl_i[FUNCT][4] ), .B(\alu_ctrl_i[FUNCT][0] ), 
        .C(\alu_ctrl_i[FUNCT][3] ), .D(n11), .E(n7), .Z(n37) );
  HS65_LH_NOR3X4 U28 ( .A(n7), .B(\alu_ctrl_i[FUNCT][1] ), .C(n43), .Z(n24) );
  HS65_LHS_XNOR2X6 U29 ( .A(\alu_ctrl_i[FUNCT][0] ), .B(n10), .Z(n31) );
  HS65_LH_CBI4I6X5 U30 ( .A(n30), .B(n29), .C(n35), .D(\alu_ctrl_i[FUNCT][0] ), 
        .Z(n44) );
  HS65_LH_IVX9 U31 ( .A(\alu_ctrl_i[OP][0] ), .Z(n17) );
  HS65_LH_IVX9 U32 ( .A(\alu_ctrl_i[FUNCT][1] ), .Z(n10) );
  HS65_LH_IVX9 U33 ( .A(\alu_ctrl_i[FUNCT][4] ), .Z(n7) );
  HS65_LH_OAI21X3 U34 ( .A(n42), .B(n24), .C(n13), .Z(n33) );
  HS65_LH_NOR3X4 U35 ( .A(n43), .B(\alu_ctrl_i[FUNCT][4] ), .C(n10), .Z(n42)
         );
  HS65_LH_IVX9 U36 ( .A(\alu_ctrl_i[OP][3] ), .Z(n12) );
  HS65_LH_IVX9 U37 ( .A(\alu_ctrl_i[OP][1] ), .Z(n16) );
  HS65_LH_NAND4ABX3 U38 ( .A(\alu_ctrl_i[FUNCT][3] ), .B(
        \alu_ctrl_i[FUNCT][2] ), .C(n6), .D(n11), .Z(n43) );
  HS65_LH_NAND4ABX3 U39 ( .A(\alu_ctrl_i[FUNCT][2] ), .B(n20), .C(n8), .D(n6), 
        .Z(n27) );
  HS65_LH_NAND2X7 U40 ( .A(n40), .B(\alu_ctrl_i[FUNCT][3] ), .Z(n35) );
  HS65_LH_IVX9 U41 ( .A(\alu_ctrl_i[OP][2] ), .Z(n14) );
  HS65_LH_AOI13X5 U42 ( .A(n32), .B(n33), .C(n34), .D(\alu_ctrl_i[OP][3] ), 
        .Z(\alu_ctrl_o[OP][1] ) );
  HS65_LH_AOI22X6 U43 ( .A(n5), .B(\alu_ctrl_i[FUNCT][0] ), .C(n15), .D(
        \alu_ctrl_i[OP][1] ), .Z(n34) );
  HS65_LH_NAND3X5 U44 ( .A(n36), .B(n10), .C(n13), .Z(n32) );
  HS65_LH_OAI32X5 U45 ( .A(n37), .B(\alu_ctrl_i[FUNCT][5] ), .C(
        \alu_ctrl_i[FUNCT][2] ), .D(\alu_ctrl_i[FUNCT][0] ), .E(n29), .Z(n36)
         );
  HS65_LH_NOR2X6 U46 ( .A(\alu_ctrl_i[OP][3] ), .B(n18), .Z(
        \alu_ctrl_o[OP][4] ) );
  HS65_LH_AOI312X4 U47 ( .A(n17), .B(n16), .C(n19), .D(\alu_ctrl_i[OP][1] ), 
        .E(\alu_ctrl_i[OP][0] ), .F(n15), .Z(n18) );
  HS65_LH_NAND4ABX3 U48 ( .A(\alu_ctrl_i[FUNCT][4] ), .B(
        \alu_ctrl_i[FUNCT][3] ), .C(\alu_ctrl_i[FUNCT][5] ), .D(
        \alu_ctrl_i[FUNCT][2] ), .Z(n29) );
  HS65_LH_NAND3X5 U49 ( .A(n14), .B(n12), .C(\alu_ctrl_i[OP][1] ), .Z(n28) );
  HS65_LH_NOR4ABX2 U50 ( .A(n11), .B(n46), .C(n8), .D(n31), .Z(n19) );
  HS65_LH_NOR3X4 U51 ( .A(\alu_ctrl_i[FUNCT][2] ), .B(\alu_ctrl_i[FUNCT][5] ), 
        .C(\alu_ctrl_i[FUNCT][4] ), .Z(n46) );
  HS65_LH_IVX9 U52 ( .A(\alu_ctrl_i[FUNCT][3] ), .Z(n8) );
  HS65_LH_NOR2X6 U53 ( .A(\alu_ctrl_i[FUNCT][4] ), .B(n10), .Z(n22) );
  HS65_LH_IVX9 U54 ( .A(\alu_ctrl_i[FUNCT][5] ), .Z(n6) );
  HS65_LH_NAND2X7 U55 ( .A(\alu_ctrl_i[OP][2] ), .B(n17), .Z(n41) );
endmodule


module exe_top_DW01_add_0 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [11:1] carry;

  HS65_LH_FA1X4 U1_1 ( .A0(A[1]), .B0(B[1]), .CI(n1), .CO(carry[2]), .S0(
        SUM[1]) );
  HS65_LH_FA1X4 U1_10 ( .A0(A[10]), .B0(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S0(SUM[10]) );
  HS65_LH_FA1X4 U1_9 ( .A0(A[9]), .B0(B[9]), .CI(carry[9]), .CO(carry[10]), 
        .S0(SUM[9]) );
  HS65_LH_FA1X4 U1_8 ( .A0(A[8]), .B0(B[8]), .CI(carry[8]), .CO(carry[9]), 
        .S0(SUM[8]) );
  HS65_LH_FA1X4 U1_7 ( .A0(A[7]), .B0(B[7]), .CI(carry[7]), .CO(carry[8]), 
        .S0(SUM[7]) );
  HS65_LH_FA1X4 U1_6 ( .A0(A[6]), .B0(B[6]), .CI(carry[6]), .CO(carry[7]), 
        .S0(SUM[6]) );
  HS65_LH_FA1X4 U1_5 ( .A0(A[5]), .B0(B[5]), .CI(carry[5]), .CO(carry[6]), 
        .S0(SUM[5]) );
  HS65_LH_FA1X4 U1_4 ( .A0(A[4]), .B0(B[4]), .CI(carry[4]), .CO(carry[5]), 
        .S0(SUM[4]) );
  HS65_LH_FA1X4 U1_3 ( .A0(A[3]), .B0(B[3]), .CI(carry[3]), .CO(carry[4]), 
        .S0(SUM[3]) );
  HS65_LH_FA1X4 U1_2 ( .A0(A[2]), .B0(B[2]), .CI(carry[2]), .CO(carry[3]), 
        .S0(SUM[2]) );
  HS65_LHS_XOR3X2 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Z(SUM[11]) );
  HS65_LH_AND2X4 U1 ( .A(A[0]), .B(B[0]), .Z(n1) );
  HS65_LHS_XOR2X6 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module exe_top ( clk, rst_n, .exe_top_i({\exe_top_i[SHAMT][4] , 
        \exe_top_i[SHAMT][3] , \exe_top_i[SHAMT][2] , \exe_top_i[SHAMT][1] , 
        \exe_top_i[SHAMT][0] , \exe_top_i[REGS_A][31] , 
        \exe_top_i[REGS_A][30] , \exe_top_i[REGS_A][29] , 
        \exe_top_i[REGS_A][28] , \exe_top_i[REGS_A][27] , 
        \exe_top_i[REGS_A][26] , \exe_top_i[REGS_A][25] , 
        \exe_top_i[REGS_A][24] , \exe_top_i[REGS_A][23] , 
        \exe_top_i[REGS_A][22] , \exe_top_i[REGS_A][21] , 
        \exe_top_i[REGS_A][20] , \exe_top_i[REGS_A][19] , 
        \exe_top_i[REGS_A][18] , \exe_top_i[REGS_A][17] , 
        \exe_top_i[REGS_A][16] , \exe_top_i[REGS_A][15] , 
        \exe_top_i[REGS_A][14] , \exe_top_i[REGS_A][13] , 
        \exe_top_i[REGS_A][12] , \exe_top_i[REGS_A][11] , 
        \exe_top_i[REGS_A][10] , \exe_top_i[REGS_A][9] , 
        \exe_top_i[REGS_A][8] , \exe_top_i[REGS_A][7] , \exe_top_i[REGS_A][6] , 
        \exe_top_i[REGS_A][5] , \exe_top_i[REGS_A][4] , \exe_top_i[REGS_A][3] , 
        \exe_top_i[REGS_A][2] , \exe_top_i[REGS_A][1] , \exe_top_i[REGS_A][0] , 
        \exe_top_i[REGS_B][31] , \exe_top_i[REGS_B][30] , 
        \exe_top_i[REGS_B][29] , \exe_top_i[REGS_B][28] , 
        \exe_top_i[REGS_B][27] , \exe_top_i[REGS_B][26] , 
        \exe_top_i[REGS_B][25] , \exe_top_i[REGS_B][24] , 
        \exe_top_i[REGS_B][23] , \exe_top_i[REGS_B][22] , 
        \exe_top_i[REGS_B][21] , \exe_top_i[REGS_B][20] , 
        \exe_top_i[REGS_B][19] , \exe_top_i[REGS_B][18] , 
        \exe_top_i[REGS_B][17] , \exe_top_i[REGS_B][16] , 
        \exe_top_i[REGS_B][15] , \exe_top_i[REGS_B][14] , 
        \exe_top_i[REGS_B][13] , \exe_top_i[REGS_B][12] , 
        \exe_top_i[REGS_B][11] , \exe_top_i[REGS_B][10] , 
        \exe_top_i[REGS_B][9] , \exe_top_i[REGS_B][8] , \exe_top_i[REGS_B][7] , 
        \exe_top_i[REGS_B][6] , \exe_top_i[REGS_B][5] , \exe_top_i[REGS_B][4] , 
        \exe_top_i[REGS_B][3] , \exe_top_i[REGS_B][2] , \exe_top_i[REGS_B][1] , 
        \exe_top_i[REGS_B][0] , \exe_top_i[ALU_SRC_B] , 
        \exe_top_i[IMMIDIATE][31] , \exe_top_i[IMMIDIATE][30] , 
        \exe_top_i[IMMIDIATE][29] , \exe_top_i[IMMIDIATE][28] , 
        \exe_top_i[IMMIDIATE][27] , \exe_top_i[IMMIDIATE][26] , 
        \exe_top_i[IMMIDIATE][25] , \exe_top_i[IMMIDIATE][24] , 
        \exe_top_i[IMMIDIATE][23] , \exe_top_i[IMMIDIATE][22] , 
        \exe_top_i[IMMIDIATE][21] , \exe_top_i[IMMIDIATE][20] , 
        \exe_top_i[IMMIDIATE][19] , \exe_top_i[IMMIDIATE][18] , 
        \exe_top_i[IMMIDIATE][17] , \exe_top_i[IMMIDIATE][16] , 
        \exe_top_i[IMMIDIATE][15] , \exe_top_i[IMMIDIATE][14] , 
        \exe_top_i[IMMIDIATE][13] , \exe_top_i[IMMIDIATE][12] , 
        \exe_top_i[IMMIDIATE][11] , \exe_top_i[IMMIDIATE][10] , 
        \exe_top_i[IMMIDIATE][9] , \exe_top_i[IMMIDIATE][8] , 
        \exe_top_i[IMMIDIATE][7] , \exe_top_i[IMMIDIATE][6] , 
        \exe_top_i[IMMIDIATE][5] , \exe_top_i[IMMIDIATE][4] , 
        \exe_top_i[IMMIDIATE][3] , \exe_top_i[IMMIDIATE][2] , 
        \exe_top_i[IMMIDIATE][1] , \exe_top_i[IMMIDIATE][0] , 
        \exe_top_i[OP][3] , \exe_top_i[OP][2] , \exe_top_i[OP][1] , 
        \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] , \exe_top_i[FUNCT][4] , 
        \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] , \exe_top_i[FUNCT][1] , 
        \exe_top_i[FUNCT][0] , \exe_top_i[PC_PLUS1][11] , 
        \exe_top_i[PC_PLUS1][10] , \exe_top_i[PC_PLUS1][9] , 
        \exe_top_i[PC_PLUS1][8] , \exe_top_i[PC_PLUS1][7] , 
        \exe_top_i[PC_PLUS1][6] , \exe_top_i[PC_PLUS1][5] , 
        \exe_top_i[PC_PLUS1][4] , \exe_top_i[PC_PLUS1][3] , 
        \exe_top_i[PC_PLUS1][2] , \exe_top_i[PC_PLUS1][1] , 
        \exe_top_i[PC_PLUS1][0] , \exe_top_i[REGDST] , \exe_top_i[RT][4] , 
        \exe_top_i[RT][3] , \exe_top_i[RT][2] , \exe_top_i[RT][1] , 
        \exe_top_i[RT][0] , \exe_top_i[RD][4] , \exe_top_i[RD][3] , 
        \exe_top_i[RD][2] , \exe_top_i[RD][1] , \exe_top_i[RD][0] }), 
    .exe_top_o({\exe_top_o[BRANCH] , \exe_top_o[BRANCH_PC][11] , 
        \exe_top_o[BRANCH_PC][10] , \exe_top_o[BRANCH_PC][9] , 
        \exe_top_o[BRANCH_PC][8] , \exe_top_o[BRANCH_PC][7] , 
        \exe_top_o[BRANCH_PC][6] , \exe_top_o[BRANCH_PC][5] , 
        \exe_top_o[BRANCH_PC][4] , \exe_top_o[BRANCH_PC][3] , 
        \exe_top_o[BRANCH_PC][2] , \exe_top_o[BRANCH_PC][1] , 
        \exe_top_o[BRANCH_PC][0] , \exe_top_o[RESULT][31] , 
        \exe_top_o[RESULT][30] , \exe_top_o[RESULT][29] , 
        \exe_top_o[RESULT][28] , \exe_top_o[RESULT][27] , 
        \exe_top_o[RESULT][26] , \exe_top_o[RESULT][25] , 
        \exe_top_o[RESULT][24] , \exe_top_o[RESULT][23] , 
        \exe_top_o[RESULT][22] , \exe_top_o[RESULT][21] , 
        \exe_top_o[RESULT][20] , \exe_top_o[RESULT][19] , 
        \exe_top_o[RESULT][18] , \exe_top_o[RESULT][17] , 
        \exe_top_o[RESULT][16] , \exe_top_o[RESULT][15] , 
        \exe_top_o[RESULT][14] , \exe_top_o[RESULT][13] , 
        \exe_top_o[RESULT][12] , \exe_top_o[RESULT][11] , 
        \exe_top_o[RESULT][10] , \exe_top_o[RESULT][9] , 
        \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] , \exe_top_o[RESULT][6] , 
        \exe_top_o[RESULT][5] , \exe_top_o[RESULT][4] , \exe_top_o[RESULT][3] , 
        \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] , \exe_top_o[RESULT][0] , 
        \exe_top_o[WRITE_REG][4] , \exe_top_o[WRITE_REG][3] , 
        \exe_top_o[WRITE_REG][2] , \exe_top_o[WRITE_REG][1] , 
        \exe_top_o[WRITE_REG][0] , \exe_top_o[DMEM_DATA][31] , 
        \exe_top_o[DMEM_DATA][30] , \exe_top_o[DMEM_DATA][29] , 
        \exe_top_o[DMEM_DATA][28] , \exe_top_o[DMEM_DATA][27] , 
        \exe_top_o[DMEM_DATA][26] , \exe_top_o[DMEM_DATA][25] , 
        \exe_top_o[DMEM_DATA][24] , \exe_top_o[DMEM_DATA][23] , 
        \exe_top_o[DMEM_DATA][22] , \exe_top_o[DMEM_DATA][21] , 
        \exe_top_o[DMEM_DATA][20] , \exe_top_o[DMEM_DATA][19] , 
        \exe_top_o[DMEM_DATA][18] , \exe_top_o[DMEM_DATA][17] , 
        \exe_top_o[DMEM_DATA][16] , \exe_top_o[DMEM_DATA][15] , 
        \exe_top_o[DMEM_DATA][14] , \exe_top_o[DMEM_DATA][13] , 
        \exe_top_o[DMEM_DATA][12] , \exe_top_o[DMEM_DATA][11] , 
        \exe_top_o[DMEM_DATA][10] , \exe_top_o[DMEM_DATA][9] , 
        \exe_top_o[DMEM_DATA][8] , \exe_top_o[DMEM_DATA][7] , 
        \exe_top_o[DMEM_DATA][6] , \exe_top_o[DMEM_DATA][5] , 
        \exe_top_o[DMEM_DATA][4] , \exe_top_o[DMEM_DATA][3] , 
        \exe_top_o[DMEM_DATA][2] , \exe_top_o[DMEM_DATA][1] , 
        \exe_top_o[DMEM_DATA][0] }) );
  input clk, rst_n, \exe_top_i[SHAMT][4] , \exe_top_i[SHAMT][3] ,
         \exe_top_i[SHAMT][2] , \exe_top_i[SHAMT][1] , \exe_top_i[SHAMT][0] ,
         \exe_top_i[REGS_A][31] , \exe_top_i[REGS_A][30] ,
         \exe_top_i[REGS_A][29] , \exe_top_i[REGS_A][28] ,
         \exe_top_i[REGS_A][27] , \exe_top_i[REGS_A][26] ,
         \exe_top_i[REGS_A][25] , \exe_top_i[REGS_A][24] ,
         \exe_top_i[REGS_A][23] , \exe_top_i[REGS_A][22] ,
         \exe_top_i[REGS_A][21] , \exe_top_i[REGS_A][20] ,
         \exe_top_i[REGS_A][19] , \exe_top_i[REGS_A][18] ,
         \exe_top_i[REGS_A][17] , \exe_top_i[REGS_A][16] ,
         \exe_top_i[REGS_A][15] , \exe_top_i[REGS_A][14] ,
         \exe_top_i[REGS_A][13] , \exe_top_i[REGS_A][12] ,
         \exe_top_i[REGS_A][11] , \exe_top_i[REGS_A][10] ,
         \exe_top_i[REGS_A][9] , \exe_top_i[REGS_A][8] ,
         \exe_top_i[REGS_A][7] , \exe_top_i[REGS_A][6] ,
         \exe_top_i[REGS_A][5] , \exe_top_i[REGS_A][4] ,
         \exe_top_i[REGS_A][3] , \exe_top_i[REGS_A][2] ,
         \exe_top_i[REGS_A][1] , \exe_top_i[REGS_A][0] ,
         \exe_top_i[REGS_B][31] , \exe_top_i[REGS_B][30] ,
         \exe_top_i[REGS_B][29] , \exe_top_i[REGS_B][28] ,
         \exe_top_i[REGS_B][27] , \exe_top_i[REGS_B][26] ,
         \exe_top_i[REGS_B][25] , \exe_top_i[REGS_B][24] ,
         \exe_top_i[REGS_B][23] , \exe_top_i[REGS_B][22] ,
         \exe_top_i[REGS_B][21] , \exe_top_i[REGS_B][20] ,
         \exe_top_i[REGS_B][19] , \exe_top_i[REGS_B][18] ,
         \exe_top_i[REGS_B][17] , \exe_top_i[REGS_B][16] ,
         \exe_top_i[REGS_B][15] , \exe_top_i[REGS_B][14] ,
         \exe_top_i[REGS_B][13] , \exe_top_i[REGS_B][12] ,
         \exe_top_i[REGS_B][11] , \exe_top_i[REGS_B][10] ,
         \exe_top_i[REGS_B][9] , \exe_top_i[REGS_B][8] ,
         \exe_top_i[REGS_B][7] , \exe_top_i[REGS_B][6] ,
         \exe_top_i[REGS_B][5] , \exe_top_i[REGS_B][4] ,
         \exe_top_i[REGS_B][3] , \exe_top_i[REGS_B][2] ,
         \exe_top_i[REGS_B][1] , \exe_top_i[REGS_B][0] ,
         \exe_top_i[ALU_SRC_B] , \exe_top_i[IMMIDIATE][31] ,
         \exe_top_i[IMMIDIATE][30] , \exe_top_i[IMMIDIATE][29] ,
         \exe_top_i[IMMIDIATE][28] , \exe_top_i[IMMIDIATE][27] ,
         \exe_top_i[IMMIDIATE][26] , \exe_top_i[IMMIDIATE][25] ,
         \exe_top_i[IMMIDIATE][24] , \exe_top_i[IMMIDIATE][23] ,
         \exe_top_i[IMMIDIATE][22] , \exe_top_i[IMMIDIATE][21] ,
         \exe_top_i[IMMIDIATE][20] , \exe_top_i[IMMIDIATE][19] ,
         \exe_top_i[IMMIDIATE][18] , \exe_top_i[IMMIDIATE][17] ,
         \exe_top_i[IMMIDIATE][16] , \exe_top_i[IMMIDIATE][15] ,
         \exe_top_i[IMMIDIATE][14] , \exe_top_i[IMMIDIATE][13] ,
         \exe_top_i[IMMIDIATE][12] , \exe_top_i[IMMIDIATE][11] ,
         \exe_top_i[IMMIDIATE][10] , \exe_top_i[IMMIDIATE][9] ,
         \exe_top_i[IMMIDIATE][8] , \exe_top_i[IMMIDIATE][7] ,
         \exe_top_i[IMMIDIATE][6] , \exe_top_i[IMMIDIATE][5] ,
         \exe_top_i[IMMIDIATE][4] , \exe_top_i[IMMIDIATE][3] ,
         \exe_top_i[IMMIDIATE][2] , \exe_top_i[IMMIDIATE][1] ,
         \exe_top_i[IMMIDIATE][0] , \exe_top_i[OP][3] , \exe_top_i[OP][2] ,
         \exe_top_i[OP][1] , \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] ,
         \exe_top_i[FUNCT][4] , \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] ,
         \exe_top_i[FUNCT][1] , \exe_top_i[FUNCT][0] ,
         \exe_top_i[PC_PLUS1][11] , \exe_top_i[PC_PLUS1][10] ,
         \exe_top_i[PC_PLUS1][9] , \exe_top_i[PC_PLUS1][8] ,
         \exe_top_i[PC_PLUS1][7] , \exe_top_i[PC_PLUS1][6] ,
         \exe_top_i[PC_PLUS1][5] , \exe_top_i[PC_PLUS1][4] ,
         \exe_top_i[PC_PLUS1][3] , \exe_top_i[PC_PLUS1][2] ,
         \exe_top_i[PC_PLUS1][1] , \exe_top_i[PC_PLUS1][0] ,
         \exe_top_i[REGDST] , \exe_top_i[RT][4] , \exe_top_i[RT][3] ,
         \exe_top_i[RT][2] , \exe_top_i[RT][1] , \exe_top_i[RT][0] ,
         \exe_top_i[RD][4] , \exe_top_i[RD][3] , \exe_top_i[RD][2] ,
         \exe_top_i[RD][1] , \exe_top_i[RD][0] ;
  output \exe_top_o[BRANCH] , \exe_top_o[BRANCH_PC][11] ,
         \exe_top_o[BRANCH_PC][10] , \exe_top_o[BRANCH_PC][9] ,
         \exe_top_o[BRANCH_PC][8] , \exe_top_o[BRANCH_PC][7] ,
         \exe_top_o[BRANCH_PC][6] , \exe_top_o[BRANCH_PC][5] ,
         \exe_top_o[BRANCH_PC][4] , \exe_top_o[BRANCH_PC][3] ,
         \exe_top_o[BRANCH_PC][2] , \exe_top_o[BRANCH_PC][1] ,
         \exe_top_o[BRANCH_PC][0] , \exe_top_o[RESULT][31] ,
         \exe_top_o[RESULT][30] , \exe_top_o[RESULT][29] ,
         \exe_top_o[RESULT][28] , \exe_top_o[RESULT][27] ,
         \exe_top_o[RESULT][26] , \exe_top_o[RESULT][25] ,
         \exe_top_o[RESULT][24] , \exe_top_o[RESULT][23] ,
         \exe_top_o[RESULT][22] , \exe_top_o[RESULT][21] ,
         \exe_top_o[RESULT][20] , \exe_top_o[RESULT][19] ,
         \exe_top_o[RESULT][18] , \exe_top_o[RESULT][17] ,
         \exe_top_o[RESULT][16] , \exe_top_o[RESULT][15] ,
         \exe_top_o[RESULT][14] , \exe_top_o[RESULT][13] ,
         \exe_top_o[RESULT][12] , \exe_top_o[RESULT][11] ,
         \exe_top_o[RESULT][10] , \exe_top_o[RESULT][9] ,
         \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] ,
         \exe_top_o[RESULT][6] , \exe_top_o[RESULT][5] ,
         \exe_top_o[RESULT][4] , \exe_top_o[RESULT][3] ,
         \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] ,
         \exe_top_o[RESULT][0] , \exe_top_o[WRITE_REG][4] ,
         \exe_top_o[WRITE_REG][3] , \exe_top_o[WRITE_REG][2] ,
         \exe_top_o[WRITE_REG][1] , \exe_top_o[WRITE_REG][0] ,
         \exe_top_o[DMEM_DATA][31] , \exe_top_o[DMEM_DATA][30] ,
         \exe_top_o[DMEM_DATA][29] , \exe_top_o[DMEM_DATA][28] ,
         \exe_top_o[DMEM_DATA][27] , \exe_top_o[DMEM_DATA][26] ,
         \exe_top_o[DMEM_DATA][25] , \exe_top_o[DMEM_DATA][24] ,
         \exe_top_o[DMEM_DATA][23] , \exe_top_o[DMEM_DATA][22] ,
         \exe_top_o[DMEM_DATA][21] , \exe_top_o[DMEM_DATA][20] ,
         \exe_top_o[DMEM_DATA][19] , \exe_top_o[DMEM_DATA][18] ,
         \exe_top_o[DMEM_DATA][17] , \exe_top_o[DMEM_DATA][16] ,
         \exe_top_o[DMEM_DATA][15] , \exe_top_o[DMEM_DATA][14] ,
         \exe_top_o[DMEM_DATA][13] , \exe_top_o[DMEM_DATA][12] ,
         \exe_top_o[DMEM_DATA][11] , \exe_top_o[DMEM_DATA][10] ,
         \exe_top_o[DMEM_DATA][9] , \exe_top_o[DMEM_DATA][8] ,
         \exe_top_o[DMEM_DATA][7] , \exe_top_o[DMEM_DATA][6] ,
         \exe_top_o[DMEM_DATA][5] , \exe_top_o[DMEM_DATA][4] ,
         \exe_top_o[DMEM_DATA][3] , \exe_top_o[DMEM_DATA][2] ,
         \exe_top_o[DMEM_DATA][1] , \exe_top_o[DMEM_DATA][0] ;
  wire   N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, n7, n8,
         n9, n10, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49;
  wire   [4:0] op_aluCtrl_alu;
  wire   [31:0] src_a;
  wire   [31:0] src_b;
  wire   [1:0] s_branch_src;

  alu alu_inst ( .clk(clk), .rst_n(n47), .alu_i({src_a, src_b, op_aluCtrl_alu, 
        \exe_top_i[SHAMT][4] , \exe_top_i[SHAMT][3] , \exe_top_i[SHAMT][2] , 
        \exe_top_i[SHAMT][1] , \exe_top_i[SHAMT][0] }), .alu_o({
        \exe_top_o[BRANCH] , \exe_top_o[RESULT][31] , \exe_top_o[RESULT][30] , 
        \exe_top_o[RESULT][29] , \exe_top_o[RESULT][28] , 
        \exe_top_o[RESULT][27] , \exe_top_o[RESULT][26] , 
        \exe_top_o[RESULT][25] , \exe_top_o[RESULT][24] , 
        \exe_top_o[RESULT][23] , \exe_top_o[RESULT][22] , 
        \exe_top_o[RESULT][21] , \exe_top_o[RESULT][20] , 
        \exe_top_o[RESULT][19] , \exe_top_o[RESULT][18] , 
        \exe_top_o[RESULT][17] , \exe_top_o[RESULT][16] , 
        \exe_top_o[RESULT][15] , \exe_top_o[RESULT][14] , 
        \exe_top_o[RESULT][13] , \exe_top_o[RESULT][12] , 
        \exe_top_o[RESULT][11] , \exe_top_o[RESULT][10] , 
        \exe_top_o[RESULT][9] , \exe_top_o[RESULT][8] , \exe_top_o[RESULT][7] , 
        \exe_top_o[RESULT][6] , \exe_top_o[RESULT][5] , \exe_top_o[RESULT][4] , 
        \exe_top_o[RESULT][3] , \exe_top_o[RESULT][2] , \exe_top_o[RESULT][1] , 
        \exe_top_o[RESULT][0] }) );
  alu_ctrl alu_ctrl_inst ( .alu_ctrl_i({\exe_top_i[OP][3] , \exe_top_i[OP][2] , 
        \exe_top_i[OP][1] , \exe_top_i[OP][0] , \exe_top_i[FUNCT][5] , 
        \exe_top_i[FUNCT][4] , \exe_top_i[FUNCT][3] , \exe_top_i[FUNCT][2] , 
        \exe_top_i[FUNCT][1] , \exe_top_i[FUNCT][0] }), .alu_ctrl_o({
        op_aluCtrl_alu, s_branch_src}) );
  exe_top_DW01_add_0 add_53 ( .A({\exe_top_i[PC_PLUS1][11] , 
        \exe_top_i[PC_PLUS1][10] , \exe_top_i[PC_PLUS1][9] , 
        \exe_top_i[PC_PLUS1][8] , \exe_top_i[PC_PLUS1][7] , 
        \exe_top_i[PC_PLUS1][6] , \exe_top_i[PC_PLUS1][5] , 
        \exe_top_i[PC_PLUS1][4] , \exe_top_i[PC_PLUS1][3] , 
        \exe_top_i[PC_PLUS1][2] , \exe_top_i[PC_PLUS1][1] , 
        \exe_top_i[PC_PLUS1][0] }), .B({\exe_top_i[IMMIDIATE][11] , 
        \exe_top_i[IMMIDIATE][10] , \exe_top_i[IMMIDIATE][9] , 
        \exe_top_i[IMMIDIATE][8] , \exe_top_i[IMMIDIATE][7] , 
        \exe_top_i[IMMIDIATE][6] , \exe_top_i[IMMIDIATE][5] , 
        \exe_top_i[IMMIDIATE][4] , \exe_top_i[IMMIDIATE][3] , 
        \exe_top_i[IMMIDIATE][2] , \exe_top_i[IMMIDIATE][1] , 
        \exe_top_i[IMMIDIATE][0] }), .CI(1'b0), .SUM({N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22}) );
  HS65_LH_NOR2AX3 U4 ( .A(\exe_top_i[REGS_A][12] ), .B(n38), .Z(src_a[12]) );
  HS65_LH_NOR2AX3 U5 ( .A(\exe_top_i[REGS_A][13] ), .B(n38), .Z(src_a[13]) );
  HS65_LH_NOR2AX3 U6 ( .A(\exe_top_i[REGS_A][15] ), .B(n38), .Z(src_a[15]) );
  HS65_LH_NOR2AX3 U7 ( .A(\exe_top_i[REGS_A][22] ), .B(n39), .Z(src_a[22]) );
  HS65_LH_NOR2AX3 U8 ( .A(\exe_top_i[REGS_A][27] ), .B(n39), .Z(src_a[27]) );
  HS65_LH_NOR2AX3 U9 ( .A(\exe_top_i[REGS_A][28] ), .B(n39), .Z(src_a[28]) );
  HS65_LH_NOR2AX3 U10 ( .A(\exe_top_i[REGS_A][16] ), .B(n38), .Z(src_a[16]) );
  HS65_LH_NOR2AX3 U11 ( .A(\exe_top_i[REGS_A][18] ), .B(n38), .Z(src_a[18]) );
  HS65_LH_NOR2AX3 U12 ( .A(\exe_top_i[REGS_A][21] ), .B(n38), .Z(src_a[21]) );
  HS65_LH_NOR2AX3 U13 ( .A(\exe_top_i[REGS_A][24] ), .B(n38), .Z(src_a[24]) );
  HS65_LH_NOR2AX3 U14 ( .A(\exe_top_i[REGS_A][30] ), .B(n38), .Z(src_a[30]) );
  HS65_LH_NOR2AX3 U15 ( .A(\exe_top_i[REGS_A][31] ), .B(n38), .Z(src_a[31]) );
  HS65_LH_BFX9 U16 ( .A(n48), .Z(n39) );
  HS65_LH_BFX9 U17 ( .A(n48), .Z(n38) );
  HS65_LH_BFX9 U18 ( .A(n48), .Z(n40) );
  HS65_LH_IVX9 U19 ( .A(n7), .Z(n48) );
  HS65_LH_IVX9 U20 ( .A(n44), .Z(n42) );
  HS65_LH_IVX9 U21 ( .A(n44), .Z(n43) );
  HS65_LH_BFX9 U22 ( .A(rst_n), .Z(n47) );
  HS65_LH_NAND3X5 U23 ( .A(op_aluCtrl_alu[4]), .B(op_aluCtrl_alu[0]), .C(n8), 
        .Z(n7) );
  HS65_LH_NOR3X4 U24 ( .A(op_aluCtrl_alu[1]), .B(op_aluCtrl_alu[3]), .C(
        op_aluCtrl_alu[2]), .Z(n8) );
  HS65_LH_BFX9 U25 ( .A(n41), .Z(n44) );
  HS65_LH_BFX9 U26 ( .A(n41), .Z(n45) );
  HS65_LH_BFX9 U27 ( .A(n41), .Z(n46) );
  HS65_LH_NOR2AX3 U28 ( .A(s_branch_src[0]), .B(s_branch_src[1]), .Z(n9) );
  HS65_LH_NOR2X6 U29 ( .A(s_branch_src[0]), .B(s_branch_src[1]), .Z(n10) );
  HS65_LH_AO22X9 U30 ( .A(\exe_top_i[REGS_A][2] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][2] ), .D(n39), .Z(src_a[2]) );
  HS65_LH_AO22X9 U31 ( .A(\exe_top_i[REGS_A][5] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][5] ), .D(n39), .Z(src_a[5]) );
  HS65_LH_AO22X9 U32 ( .A(\exe_top_i[REGS_A][8] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][8] ), .D(n39), .Z(src_a[8]) );
  HS65_LH_AO22X9 U33 ( .A(\exe_top_i[REGS_A][0] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][0] ), .D(n40), .Z(src_a[0]) );
  HS65_LH_AO22X9 U34 ( .A(\exe_top_i[REGS_A][4] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][4] ), .D(n39), .Z(src_a[4]) );
  HS65_LH_AO22X9 U35 ( .A(\exe_top_i[REGS_A][1] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][1] ), .D(n40), .Z(src_a[1]) );
  HS65_LH_AO22X9 U36 ( .A(\exe_top_i[REGS_A][3] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][3] ), .D(n39), .Z(src_a[3]) );
  HS65_LH_AO22X9 U37 ( .A(\exe_top_i[IMMIDIATE][2] ), .B(n46), .C(
        \exe_top_i[REGS_B][2] ), .D(n43), .Z(src_b[2]) );
  HS65_LH_AO22X9 U38 ( .A(\exe_top_i[IMMIDIATE][0] ), .B(n44), .C(
        \exe_top_i[REGS_B][0] ), .D(n42), .Z(src_b[0]) );
  HS65_LH_AO22X9 U39 ( .A(\exe_top_i[IMMIDIATE][4] ), .B(n46), .C(
        \exe_top_i[REGS_B][4] ), .D(n43), .Z(src_b[4]) );
  HS65_LH_AO22X9 U40 ( .A(\exe_top_i[REGS_A][11] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][11] ), .D(n40), .Z(src_a[11]) );
  HS65_LH_NOR2AX3 U41 ( .A(\exe_top_i[REGS_A][14] ), .B(n38), .Z(src_a[14]) );
  HS65_LH_NOR2AX3 U42 ( .A(\exe_top_i[REGS_A][17] ), .B(n38), .Z(src_a[17]) );
  HS65_LH_NOR2AX3 U43 ( .A(\exe_top_i[REGS_A][20] ), .B(n39), .Z(src_a[20]) );
  HS65_LH_AO22X9 U44 ( .A(\exe_top_i[REGS_A][10] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][10] ), .D(n40), .Z(src_a[10]) );
  HS65_LH_AO22X9 U45 ( .A(\exe_top_i[REGS_A][6] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][6] ), .D(n39), .Z(src_a[6]) );
  HS65_LH_AO22X9 U46 ( .A(\exe_top_i[REGS_A][7] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][7] ), .D(n39), .Z(src_a[7]) );
  HS65_LH_AO22X9 U47 ( .A(\exe_top_i[REGS_A][9] ), .B(n7), .C(
        \exe_top_i[PC_PLUS1][9] ), .D(n39), .Z(src_a[9]) );
  HS65_LH_AO22X9 U48 ( .A(\exe_top_i[IMMIDIATE][7] ), .B(n46), .C(
        \exe_top_i[REGS_B][7] ), .D(n43), .Z(src_b[7]) );
  HS65_LH_AO22X9 U49 ( .A(\exe_top_i[IMMIDIATE][5] ), .B(n46), .C(
        \exe_top_i[REGS_B][5] ), .D(n43), .Z(src_b[5]) );
  HS65_LH_AO22X9 U50 ( .A(\exe_top_i[IMMIDIATE][1] ), .B(n45), .C(
        \exe_top_i[REGS_B][1] ), .D(n42), .Z(src_b[1]) );
  HS65_LH_AO22X9 U51 ( .A(\exe_top_i[IMMIDIATE][3] ), .B(n46), .C(
        \exe_top_i[REGS_B][3] ), .D(n43), .Z(src_b[3]) );
  HS65_LH_AO22X9 U52 ( .A(\exe_top_i[IMMIDIATE][6] ), .B(n46), .C(
        \exe_top_i[REGS_B][6] ), .D(n43), .Z(src_b[6]) );
  HS65_LH_AO22X9 U53 ( .A(\exe_top_i[IMMIDIATE][8] ), .B(n46), .C(
        \exe_top_i[REGS_B][8] ), .D(n43), .Z(src_b[8]) );
  HS65_LH_AO22X9 U54 ( .A(\exe_top_i[IMMIDIATE][11] ), .B(n45), .C(
        \exe_top_i[REGS_B][11] ), .D(n42), .Z(src_b[11]) );
  HS65_LH_NOR2AX3 U55 ( .A(\exe_top_i[REGS_A][25] ), .B(n39), .Z(src_a[25]) );
  HS65_LH_NOR2AX3 U56 ( .A(\exe_top_i[REGS_A][19] ), .B(n38), .Z(src_a[19]) );
  HS65_LH_NOR2AX3 U57 ( .A(\exe_top_i[REGS_A][23] ), .B(n38), .Z(src_a[23]) );
  HS65_LH_NOR2AX3 U58 ( .A(\exe_top_i[REGS_A][26] ), .B(n39), .Z(src_a[26]) );
  HS65_LH_AO22X9 U59 ( .A(\exe_top_i[IMMIDIATE][13] ), .B(n45), .C(
        \exe_top_i[REGS_B][13] ), .D(n42), .Z(src_b[13]) );
  HS65_LH_AO22X9 U60 ( .A(\exe_top_i[IMMIDIATE][12] ), .B(n45), .C(
        \exe_top_i[REGS_B][12] ), .D(n42), .Z(src_b[12]) );
  HS65_LH_AO22X9 U61 ( .A(\exe_top_i[IMMIDIATE][9] ), .B(n46), .C(
        \exe_top_i[REGS_B][9] ), .D(n43), .Z(src_b[9]) );
  HS65_LH_AO22X9 U62 ( .A(\exe_top_i[IMMIDIATE][14] ), .B(n45), .C(
        \exe_top_i[REGS_B][14] ), .D(n42), .Z(src_b[14]) );
  HS65_LH_AO22X9 U63 ( .A(\exe_top_i[IMMIDIATE][10] ), .B(n45), .C(
        \exe_top_i[REGS_B][10] ), .D(n42), .Z(src_b[10]) );
  HS65_LH_NOR2AX3 U64 ( .A(\exe_top_i[REGS_A][29] ), .B(n39), .Z(src_a[29]) );
  HS65_LH_AO22X9 U65 ( .A(\exe_top_i[IMMIDIATE][19] ), .B(n45), .C(
        \exe_top_i[REGS_B][19] ), .D(n42), .Z(src_b[19]) );
  HS65_LH_AO22X9 U66 ( .A(\exe_top_i[IMMIDIATE][15] ), .B(n45), .C(
        \exe_top_i[REGS_B][15] ), .D(n42), .Z(src_b[15]) );
  HS65_LH_AO22X9 U67 ( .A(\exe_top_i[IMMIDIATE][21] ), .B(n45), .C(
        \exe_top_i[REGS_B][21] ), .D(n43), .Z(src_b[21]) );
  HS65_LH_AO22X9 U68 ( .A(\exe_top_i[IMMIDIATE][17] ), .B(n45), .C(
        \exe_top_i[REGS_B][17] ), .D(n42), .Z(src_b[17]) );
  HS65_LH_AO22X9 U69 ( .A(\exe_top_i[IMMIDIATE][18] ), .B(n45), .C(
        \exe_top_i[REGS_B][18] ), .D(n42), .Z(src_b[18]) );
  HS65_LH_AO22X9 U70 ( .A(\exe_top_i[IMMIDIATE][20] ), .B(n45), .C(
        \exe_top_i[REGS_B][20] ), .D(n43), .Z(src_b[20]) );
  HS65_LH_AO22X9 U71 ( .A(\exe_top_i[IMMIDIATE][16] ), .B(n45), .C(
        \exe_top_i[REGS_B][16] ), .D(n42), .Z(src_b[16]) );
  HS65_LH_BFX9 U72 ( .A(\exe_top_i[ALU_SRC_B] ), .Z(n41) );
  HS65_LH_AO22X9 U73 ( .A(\exe_top_i[IMMIDIATE][23] ), .B(n45), .C(
        \exe_top_i[REGS_B][23] ), .D(n43), .Z(src_b[23]) );
  HS65_LH_AO22X9 U74 ( .A(\exe_top_i[IMMIDIATE][25] ), .B(n45), .C(
        \exe_top_i[REGS_B][25] ), .D(n43), .Z(src_b[25]) );
  HS65_LH_AO22X9 U75 ( .A(\exe_top_i[IMMIDIATE][22] ), .B(n45), .C(
        \exe_top_i[REGS_B][22] ), .D(n43), .Z(src_b[22]) );
  HS65_LH_AO22X9 U76 ( .A(\exe_top_i[IMMIDIATE][26] ), .B(n45), .C(
        \exe_top_i[REGS_B][26] ), .D(n43), .Z(src_b[26]) );
  HS65_LH_AO22X9 U77 ( .A(\exe_top_i[IMMIDIATE][24] ), .B(n45), .C(
        \exe_top_i[REGS_B][24] ), .D(n43), .Z(src_b[24]) );
  HS65_LH_AO22X9 U78 ( .A(\exe_top_i[IMMIDIATE][28] ), .B(n45), .C(
        \exe_top_i[REGS_B][28] ), .D(n43), .Z(src_b[28]) );
  HS65_LH_AO22X9 U79 ( .A(\exe_top_i[IMMIDIATE][27] ), .B(n45), .C(
        \exe_top_i[REGS_B][27] ), .D(n43), .Z(src_b[27]) );
  HS65_LH_AO22X9 U80 ( .A(\exe_top_i[IMMIDIATE][29] ), .B(n46), .C(
        \exe_top_i[REGS_B][29] ), .D(n43), .Z(src_b[29]) );
  HS65_LH_AO22X9 U81 ( .A(\exe_top_i[IMMIDIATE][30] ), .B(n46), .C(
        \exe_top_i[REGS_B][30] ), .D(n43), .Z(src_b[30]) );
  HS65_LH_AO22X9 U82 ( .A(\exe_top_i[IMMIDIATE][31] ), .B(n46), .C(
        \exe_top_i[REGS_B][31] ), .D(n43), .Z(src_b[31]) );
  HS65_LH_AO222X4 U83 ( .A(n9), .B(\exe_top_i[REGS_A][9] ), .C(N31), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][9] ), .Z(
        \exe_top_o[BRANCH_PC][9] ) );
  HS65_LH_AO222X4 U84 ( .A(n9), .B(\exe_top_i[REGS_A][0] ), .C(N22), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][0] ), .Z(
        \exe_top_o[BRANCH_PC][0] ) );
  HS65_LH_AO222X4 U85 ( .A(n9), .B(\exe_top_i[REGS_A][1] ), .C(N23), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][1] ), .Z(
        \exe_top_o[BRANCH_PC][1] ) );
  HS65_LH_AO222X4 U86 ( .A(n9), .B(\exe_top_i[REGS_A][2] ), .C(N24), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][2] ), .Z(
        \exe_top_o[BRANCH_PC][2] ) );
  HS65_LH_AO222X4 U87 ( .A(n9), .B(\exe_top_i[REGS_A][3] ), .C(N25), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][3] ), .Z(
        \exe_top_o[BRANCH_PC][3] ) );
  HS65_LH_AO222X4 U88 ( .A(n9), .B(\exe_top_i[REGS_A][4] ), .C(N26), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][4] ), .Z(
        \exe_top_o[BRANCH_PC][4] ) );
  HS65_LH_AO222X4 U89 ( .A(n9), .B(\exe_top_i[REGS_A][5] ), .C(N27), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][5] ), .Z(
        \exe_top_o[BRANCH_PC][5] ) );
  HS65_LH_AO222X4 U90 ( .A(n9), .B(\exe_top_i[REGS_A][6] ), .C(N28), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][6] ), .Z(
        \exe_top_o[BRANCH_PC][6] ) );
  HS65_LH_AO222X4 U91 ( .A(n9), .B(\exe_top_i[REGS_A][7] ), .C(N29), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][7] ), .Z(
        \exe_top_o[BRANCH_PC][7] ) );
  HS65_LH_AO222X4 U92 ( .A(n9), .B(\exe_top_i[REGS_A][8] ), .C(N30), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][8] ), .Z(
        \exe_top_o[BRANCH_PC][8] ) );
  HS65_LH_AO222X4 U93 ( .A(n9), .B(\exe_top_i[REGS_A][10] ), .C(N32), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][10] ), .Z(
        \exe_top_o[BRANCH_PC][10] ) );
  HS65_LH_AO222X4 U94 ( .A(n9), .B(\exe_top_i[REGS_A][11] ), .C(N33), .D(n10), 
        .E(s_branch_src[1]), .F(\exe_top_i[IMMIDIATE][11] ), .Z(
        \exe_top_o[BRANCH_PC][11] ) );
  HS65_LH_BFX9 U95 ( .A(\exe_top_i[REGS_B][9] ), .Z(\exe_top_o[DMEM_DATA][9] )
         );
  HS65_LH_BFX9 U96 ( .A(\exe_top_i[REGS_B][12] ), .Z(
        \exe_top_o[DMEM_DATA][12] ) );
  HS65_LH_BFX9 U97 ( .A(\exe_top_i[REGS_B][13] ), .Z(
        \exe_top_o[DMEM_DATA][13] ) );
  HS65_LH_BFX9 U98 ( .A(\exe_top_i[REGS_B][14] ), .Z(
        \exe_top_o[DMEM_DATA][14] ) );
  HS65_LH_BFX9 U99 ( .A(\exe_top_i[REGS_B][15] ), .Z(
        \exe_top_o[DMEM_DATA][15] ) );
  HS65_LH_BFX9 U100 ( .A(\exe_top_i[REGS_B][16] ), .Z(
        \exe_top_o[DMEM_DATA][16] ) );
  HS65_LH_BFX9 U101 ( .A(\exe_top_i[REGS_B][17] ), .Z(
        \exe_top_o[DMEM_DATA][17] ) );
  HS65_LH_BFX9 U102 ( .A(\exe_top_i[REGS_B][18] ), .Z(
        \exe_top_o[DMEM_DATA][18] ) );
  HS65_LH_BFX9 U103 ( .A(\exe_top_i[REGS_B][19] ), .Z(
        \exe_top_o[DMEM_DATA][19] ) );
  HS65_LH_BFX9 U104 ( .A(\exe_top_i[REGS_B][20] ), .Z(
        \exe_top_o[DMEM_DATA][20] ) );
  HS65_LH_BFX9 U105 ( .A(\exe_top_i[REGS_B][21] ), .Z(
        \exe_top_o[DMEM_DATA][21] ) );
  HS65_LH_BFX9 U106 ( .A(\exe_top_i[REGS_B][22] ), .Z(
        \exe_top_o[DMEM_DATA][22] ) );
  HS65_LH_BFX9 U107 ( .A(\exe_top_i[REGS_B][23] ), .Z(
        \exe_top_o[DMEM_DATA][23] ) );
  HS65_LH_BFX9 U108 ( .A(\exe_top_i[REGS_B][24] ), .Z(
        \exe_top_o[DMEM_DATA][24] ) );
  HS65_LH_BFX9 U109 ( .A(\exe_top_i[REGS_B][25] ), .Z(
        \exe_top_o[DMEM_DATA][25] ) );
  HS65_LH_BFX9 U110 ( .A(\exe_top_i[REGS_B][26] ), .Z(
        \exe_top_o[DMEM_DATA][26] ) );
  HS65_LH_BFX9 U111 ( .A(\exe_top_i[REGS_B][27] ), .Z(
        \exe_top_o[DMEM_DATA][27] ) );
  HS65_LH_BFX9 U112 ( .A(\exe_top_i[REGS_B][28] ), .Z(
        \exe_top_o[DMEM_DATA][28] ) );
  HS65_LH_BFX9 U113 ( .A(\exe_top_i[REGS_B][29] ), .Z(
        \exe_top_o[DMEM_DATA][29] ) );
  HS65_LH_BFX9 U114 ( .A(\exe_top_i[REGS_B][30] ), .Z(
        \exe_top_o[DMEM_DATA][30] ) );
  HS65_LH_BFX9 U115 ( .A(\exe_top_i[REGS_B][31] ), .Z(
        \exe_top_o[DMEM_DATA][31] ) );
  HS65_LH_BFX9 U116 ( .A(\exe_top_i[REGS_B][0] ), .Z(\exe_top_o[DMEM_DATA][0] ) );
  HS65_LH_BFX9 U117 ( .A(\exe_top_i[REGS_B][1] ), .Z(\exe_top_o[DMEM_DATA][1] ) );
  HS65_LH_BFX9 U118 ( .A(\exe_top_i[REGS_B][2] ), .Z(\exe_top_o[DMEM_DATA][2] ) );
  HS65_LH_BFX9 U119 ( .A(\exe_top_i[REGS_B][3] ), .Z(\exe_top_o[DMEM_DATA][3] ) );
  HS65_LH_BFX9 U120 ( .A(\exe_top_i[REGS_B][4] ), .Z(\exe_top_o[DMEM_DATA][4] ) );
  HS65_LH_BFX9 U121 ( .A(\exe_top_i[REGS_B][5] ), .Z(\exe_top_o[DMEM_DATA][5] ) );
  HS65_LH_BFX9 U122 ( .A(\exe_top_i[REGS_B][6] ), .Z(\exe_top_o[DMEM_DATA][6] ) );
  HS65_LH_BFX9 U123 ( .A(\exe_top_i[REGS_B][7] ), .Z(\exe_top_o[DMEM_DATA][7] ) );
  HS65_LH_BFX9 U124 ( .A(\exe_top_i[REGS_B][8] ), .Z(\exe_top_o[DMEM_DATA][8] ) );
  HS65_LH_BFX9 U125 ( .A(\exe_top_i[REGS_B][10] ), .Z(
        \exe_top_o[DMEM_DATA][10] ) );
  HS65_LH_BFX9 U126 ( .A(\exe_top_i[REGS_B][11] ), .Z(
        \exe_top_o[DMEM_DATA][11] ) );
  HS65_LH_AO212X4 U127 ( .A(\exe_top_i[RD][0] ), .B(\exe_top_i[REGDST] ), .C(
        \exe_top_i[RT][0] ), .D(n49), .E(n40), .Z(\exe_top_o[WRITE_REG][0] )
         );
  HS65_LH_AO212X4 U128 ( .A(\exe_top_i[RD][1] ), .B(\exe_top_i[REGDST] ), .C(
        \exe_top_i[RT][1] ), .D(n49), .E(n40), .Z(\exe_top_o[WRITE_REG][1] )
         );
  HS65_LH_AO212X4 U129 ( .A(\exe_top_i[RD][2] ), .B(\exe_top_i[REGDST] ), .C(
        \exe_top_i[RT][2] ), .D(n49), .E(n40), .Z(\exe_top_o[WRITE_REG][2] )
         );
  HS65_LH_AO212X4 U130 ( .A(\exe_top_i[RD][3] ), .B(\exe_top_i[REGDST] ), .C(
        \exe_top_i[RT][3] ), .D(n49), .E(n40), .Z(\exe_top_o[WRITE_REG][3] )
         );
  HS65_LH_AO212X4 U131 ( .A(\exe_top_i[REGDST] ), .B(\exe_top_i[RD][4] ), .C(
        \exe_top_i[RT][4] ), .D(n49), .E(n40), .Z(\exe_top_o[WRITE_REG][4] )
         );
  HS65_LH_IVX9 U132 ( .A(\exe_top_i[REGDST] ), .Z(n49) );
endmodule


module forwarding_unit ( .forwarding_unit_i({\forwarding_unit_i[EXE_IN_RS][4] , 
        \forwarding_unit_i[EXE_IN_RS][3] , \forwarding_unit_i[EXE_IN_RS][2] , 
        \forwarding_unit_i[EXE_IN_RS][1] , \forwarding_unit_i[EXE_IN_RS][0] , 
        \forwarding_unit_i[EXE_IN_RT][4] , \forwarding_unit_i[EXE_IN_RT][3] , 
        \forwarding_unit_i[EXE_IN_RT][2] , \forwarding_unit_i[EXE_IN_RT][1] , 
        \forwarding_unit_i[EXE_IN_RT][0] , \forwarding_unit_i[ID_OUT_RS][4] , 
        \forwarding_unit_i[ID_OUT_RS][3] , \forwarding_unit_i[ID_OUT_RS][2] , 
        \forwarding_unit_i[ID_OUT_RS][1] , \forwarding_unit_i[ID_OUT_RS][0] , 
        \forwarding_unit_i[ID_OUT_RT][4] , \forwarding_unit_i[ID_OUT_RT][3] , 
        \forwarding_unit_i[ID_OUT_RT][2] , \forwarding_unit_i[ID_OUT_RT][1] , 
        \forwarding_unit_i[ID_OUT_RT][0] , 
        \forwarding_unit_i[MEM_IN_WRITE_REG][4] , 
        \forwarding_unit_i[MEM_IN_WRITE_REG][3] , 
        \forwarding_unit_i[MEM_IN_WRITE_REG][2] , 
        \forwarding_unit_i[MEM_IN_WRITE_REG][1] , 
        \forwarding_unit_i[MEM_IN_WRITE_REG][0] , 
        \forwarding_unit_i[WB_IN_WRITE_REG][4] , 
        \forwarding_unit_i[WB_IN_WRITE_REG][3] , 
        \forwarding_unit_i[WB_IN_WRITE_REG][2] , 
        \forwarding_unit_i[WB_IN_WRITE_REG][1] , 
        \forwarding_unit_i[WB_IN_WRITE_REG][0] , 
        \forwarding_unit_i[MEM_IN_REGWRITE] , 
        \forwarding_unit_i[WB_IN_REGWRITE] }), .forwarding_unit_o({
        \forwarding_unit_o[FORWARD_A][1] , \forwarding_unit_o[FORWARD_A][0] , 
        \forwarding_unit_o[FORWARD_B][1] , \forwarding_unit_o[FORWARD_B][0] , 
        \forwarding_unit_o[REGFILE_FORWARD_A] , 
        \forwarding_unit_o[REGFILE_FORWARD_B] }) );
  input \forwarding_unit_i[EXE_IN_RS][4] , \forwarding_unit_i[EXE_IN_RS][3] ,
         \forwarding_unit_i[EXE_IN_RS][2] , \forwarding_unit_i[EXE_IN_RS][1] ,
         \forwarding_unit_i[EXE_IN_RS][0] , \forwarding_unit_i[EXE_IN_RT][4] ,
         \forwarding_unit_i[EXE_IN_RT][3] , \forwarding_unit_i[EXE_IN_RT][2] ,
         \forwarding_unit_i[EXE_IN_RT][1] , \forwarding_unit_i[EXE_IN_RT][0] ,
         \forwarding_unit_i[ID_OUT_RS][4] , \forwarding_unit_i[ID_OUT_RS][3] ,
         \forwarding_unit_i[ID_OUT_RS][2] , \forwarding_unit_i[ID_OUT_RS][1] ,
         \forwarding_unit_i[ID_OUT_RS][0] , \forwarding_unit_i[ID_OUT_RT][4] ,
         \forwarding_unit_i[ID_OUT_RT][3] , \forwarding_unit_i[ID_OUT_RT][2] ,
         \forwarding_unit_i[ID_OUT_RT][1] , \forwarding_unit_i[ID_OUT_RT][0] ,
         \forwarding_unit_i[MEM_IN_WRITE_REG][4] ,
         \forwarding_unit_i[MEM_IN_WRITE_REG][3] ,
         \forwarding_unit_i[MEM_IN_WRITE_REG][2] ,
         \forwarding_unit_i[MEM_IN_WRITE_REG][1] ,
         \forwarding_unit_i[MEM_IN_WRITE_REG][0] ,
         \forwarding_unit_i[WB_IN_WRITE_REG][4] ,
         \forwarding_unit_i[WB_IN_WRITE_REG][3] ,
         \forwarding_unit_i[WB_IN_WRITE_REG][2] ,
         \forwarding_unit_i[WB_IN_WRITE_REG][1] ,
         \forwarding_unit_i[WB_IN_WRITE_REG][0] ,
         \forwarding_unit_i[MEM_IN_REGWRITE] ,
         \forwarding_unit_i[WB_IN_REGWRITE] ;
  output \forwarding_unit_o[FORWARD_A][1] , \forwarding_unit_o[FORWARD_A][0] ,
         \forwarding_unit_o[FORWARD_B][1] , \forwarding_unit_o[FORWARD_B][0] ,
         \forwarding_unit_o[REGFILE_FORWARD_A] ,
         \forwarding_unit_o[REGFILE_FORWARD_B] ;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n1;

  HS65_LH_NOR4ABX2 U2 ( .A(n58), .B(n59), .C(n60), .D(n61), .Z(
        \forwarding_unit_o[FORWARD_A][1] ) );
  HS65_LH_NOR4ABX2 U3 ( .A(n45), .B(n46), .C(n47), .D(n48), .Z(
        \forwarding_unit_o[FORWARD_B][1] ) );
  HS65_LHS_XOR2X6 U4 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][0] ), .B(
        \forwarding_unit_i[EXE_IN_RS][0] ), .Z(n60) );
  HS65_LHS_XNOR2X6 U5 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][3] ), .B(
        \forwarding_unit_i[EXE_IN_RS][3] ), .Z(n59) );
  HS65_LHS_XNOR2X6 U6 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][1] ), .B(
        \forwarding_unit_i[EXE_IN_RS][1] ), .Z(n58) );
  HS65_LH_NOR4ABX2 U7 ( .A(n51), .B(n52), .C(n53), .D(n54), .Z(
        \forwarding_unit_o[FORWARD_A][0] ) );
  HS65_LHS_XNOR2X6 U8 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][3] ), .B(
        \forwarding_unit_i[EXE_IN_RS][3] ), .Z(n51) );
  HS65_LHS_XOR2X6 U9 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][0] ), .B(
        \forwarding_unit_i[EXE_IN_RS][0] ), .Z(n54) );
  HS65_LHS_XNOR2X6 U10 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][1] ), .B(
        \forwarding_unit_i[EXE_IN_RS][1] ), .Z(n52) );
  HS65_LH_OA31X9 U11 ( .A(n57), .B(\forwarding_unit_i[WB_IN_WRITE_REG][1] ), 
        .C(\forwarding_unit_i[WB_IN_WRITE_REG][0] ), .D(
        \forwarding_unit_i[WB_IN_REGWRITE] ), .Z(n27) );
  HS65_LH_OR3X9 U12 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][3] ), .C(
        \forwarding_unit_i[WB_IN_WRITE_REG][2] ), .Z(n57) );
  HS65_LH_NAND4ABX3 U13 ( .A(n62), .B(n63), .C(
        \forwarding_unit_i[MEM_IN_REGWRITE] ), .D(n1), .Z(n61) );
  HS65_LHS_XOR2X6 U14 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][2] ), .B(
        \forwarding_unit_i[EXE_IN_RS][2] ), .Z(n63) );
  HS65_LHS_XOR2X6 U15 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[EXE_IN_RS][4] ), .Z(n62) );
  HS65_LH_NAND4ABX3 U16 ( .A(n55), .B(\forwarding_unit_o[FORWARD_A][1] ), .C(
        n56), .D(n27), .Z(n53) );
  HS65_LHS_XNOR2X6 U17 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][2] ), .B(
        \forwarding_unit_i[EXE_IN_RS][2] ), .Z(n56) );
  HS65_LHS_XOR2X6 U18 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[EXE_IN_RS][4] ), .Z(n55) );
  HS65_LH_IVX9 U19 ( .A(n64), .Z(n1) );
  HS65_LH_NOR3AX2 U20 ( .A(n65), .B(\forwarding_unit_i[MEM_IN_WRITE_REG][0] ), 
        .C(\forwarding_unit_i[MEM_IN_WRITE_REG][1] ), .Z(n64) );
  HS65_LH_NOR3X4 U21 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][2] ), .B(
        \forwarding_unit_i[MEM_IN_WRITE_REG][4] ), .C(
        \forwarding_unit_i[MEM_IN_WRITE_REG][3] ), .Z(n65) );
  HS65_LHS_XOR2X6 U22 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][3] ), .B(
        \forwarding_unit_i[EXE_IN_RT][3] ), .Z(n47) );
  HS65_LHS_XNOR2X6 U23 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][0] ), .B(
        \forwarding_unit_i[EXE_IN_RT][0] ), .Z(n46) );
  HS65_LHS_XNOR2X6 U24 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][1] ), .B(
        \forwarding_unit_i[EXE_IN_RT][1] ), .Z(n45) );
  HS65_LH_NOR4ABX2 U25 ( .A(n39), .B(n40), .C(n41), .D(n42), .Z(
        \forwarding_unit_o[FORWARD_B][0] ) );
  HS65_LHS_XNOR2X6 U26 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][3] ), .B(
        \forwarding_unit_i[EXE_IN_RT][3] ), .Z(n39) );
  HS65_LHS_XOR2X6 U27 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][0] ), .B(
        \forwarding_unit_i[EXE_IN_RT][0] ), .Z(n42) );
  HS65_LHS_XNOR2X6 U28 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][1] ), .B(
        \forwarding_unit_i[EXE_IN_RT][1] ), .Z(n40) );
  HS65_LH_NAND4ABX3 U29 ( .A(n49), .B(n50), .C(
        \forwarding_unit_i[MEM_IN_REGWRITE] ), .D(n1), .Z(n48) );
  HS65_LHS_XOR2X6 U30 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][2] ), .B(
        \forwarding_unit_i[EXE_IN_RT][2] ), .Z(n50) );
  HS65_LHS_XOR2X6 U31 ( .A(\forwarding_unit_i[MEM_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[EXE_IN_RT][4] ), .Z(n49) );
  HS65_LH_NAND4ABX3 U32 ( .A(n43), .B(\forwarding_unit_o[FORWARD_B][1] ), .C(
        n44), .D(n27), .Z(n41) );
  HS65_LHS_XNOR2X6 U33 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][2] ), .B(
        \forwarding_unit_i[EXE_IN_RT][2] ), .Z(n44) );
  HS65_LHS_XOR2X6 U34 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[EXE_IN_RT][4] ), .Z(n43) );
  HS65_LH_NOR4ABX2 U35 ( .A(n33), .B(n27), .C(n34), .D(n35), .Z(
        \forwarding_unit_o[REGFILE_FORWARD_A] ) );
  HS65_LHS_XOR2X6 U36 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[ID_OUT_RS][4] ), .Z(n35) );
  HS65_LHS_XNOR2X6 U37 ( .A(\forwarding_unit_i[ID_OUT_RS][2] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][2] ), .Z(n33) );
  HS65_LH_NOR4ABX2 U38 ( .A(n26), .B(n27), .C(n28), .D(n29), .Z(
        \forwarding_unit_o[REGFILE_FORWARD_B] ) );
  HS65_LHS_XOR2X6 U39 ( .A(\forwarding_unit_i[WB_IN_WRITE_REG][4] ), .B(
        \forwarding_unit_i[ID_OUT_RT][4] ), .Z(n29) );
  HS65_LHS_XNOR2X6 U40 ( .A(\forwarding_unit_i[ID_OUT_RT][3] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][3] ), .Z(n26) );
  HS65_LH_NAND3X5 U41 ( .A(n30), .B(n31), .C(n32), .Z(n28) );
  HS65_LHS_XNOR2X6 U42 ( .A(\forwarding_unit_i[ID_OUT_RT][1] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][1] ), .Z(n32) );
  HS65_LHS_XNOR2X6 U43 ( .A(\forwarding_unit_i[ID_OUT_RT][2] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][2] ), .Z(n31) );
  HS65_LHS_XNOR2X6 U44 ( .A(\forwarding_unit_i[ID_OUT_RT][0] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][0] ), .Z(n30) );
  HS65_LH_NAND3X5 U45 ( .A(n36), .B(n37), .C(n38), .Z(n34) );
  HS65_LHS_XNOR2X6 U46 ( .A(\forwarding_unit_i[ID_OUT_RS][1] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][1] ), .Z(n38) );
  HS65_LHS_XNOR2X6 U47 ( .A(\forwarding_unit_i[ID_OUT_RS][3] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][3] ), .Z(n36) );
  HS65_LHS_XNOR2X6 U48 ( .A(\forwarding_unit_i[ID_OUT_RS][0] ), .B(
        \forwarding_unit_i[WB_IN_WRITE_REG][0] ), .Z(n37) );
endmodule


module exe_mem ( clk, rst_n, halt_i, .EXE_MEM_i({\EXE_MEM_i[ALU_RES][31] , 
        \EXE_MEM_i[ALU_RES][30] , \EXE_MEM_i[ALU_RES][29] , 
        \EXE_MEM_i[ALU_RES][28] , \EXE_MEM_i[ALU_RES][27] , 
        \EXE_MEM_i[ALU_RES][26] , \EXE_MEM_i[ALU_RES][25] , 
        \EXE_MEM_i[ALU_RES][24] , \EXE_MEM_i[ALU_RES][23] , 
        \EXE_MEM_i[ALU_RES][22] , \EXE_MEM_i[ALU_RES][21] , 
        \EXE_MEM_i[ALU_RES][20] , \EXE_MEM_i[ALU_RES][19] , 
        \EXE_MEM_i[ALU_RES][18] , \EXE_MEM_i[ALU_RES][17] , 
        \EXE_MEM_i[ALU_RES][16] , \EXE_MEM_i[ALU_RES][15] , 
        \EXE_MEM_i[ALU_RES][14] , \EXE_MEM_i[ALU_RES][13] , 
        \EXE_MEM_i[ALU_RES][12] , \EXE_MEM_i[ALU_RES][11] , 
        \EXE_MEM_i[ALU_RES][10] , \EXE_MEM_i[ALU_RES][9] , 
        \EXE_MEM_i[ALU_RES][8] , \EXE_MEM_i[ALU_RES][7] , 
        \EXE_MEM_i[ALU_RES][6] , \EXE_MEM_i[ALU_RES][5] , 
        \EXE_MEM_i[ALU_RES][4] , \EXE_MEM_i[ALU_RES][3] , 
        \EXE_MEM_i[ALU_RES][2] , \EXE_MEM_i[ALU_RES][1] , 
        \EXE_MEM_i[ALU_RES][0] , \EXE_MEM_i[DMEM_DATA][31] , 
        \EXE_MEM_i[DMEM_DATA][30] , \EXE_MEM_i[DMEM_DATA][29] , 
        \EXE_MEM_i[DMEM_DATA][28] , \EXE_MEM_i[DMEM_DATA][27] , 
        \EXE_MEM_i[DMEM_DATA][26] , \EXE_MEM_i[DMEM_DATA][25] , 
        \EXE_MEM_i[DMEM_DATA][24] , \EXE_MEM_i[DMEM_DATA][23] , 
        \EXE_MEM_i[DMEM_DATA][22] , \EXE_MEM_i[DMEM_DATA][21] , 
        \EXE_MEM_i[DMEM_DATA][20] , \EXE_MEM_i[DMEM_DATA][19] , 
        \EXE_MEM_i[DMEM_DATA][18] , \EXE_MEM_i[DMEM_DATA][17] , 
        \EXE_MEM_i[DMEM_DATA][16] , \EXE_MEM_i[DMEM_DATA][15] , 
        \EXE_MEM_i[DMEM_DATA][14] , \EXE_MEM_i[DMEM_DATA][13] , 
        \EXE_MEM_i[DMEM_DATA][12] , \EXE_MEM_i[DMEM_DATA][11] , 
        \EXE_MEM_i[DMEM_DATA][10] , \EXE_MEM_i[DMEM_DATA][9] , 
        \EXE_MEM_i[DMEM_DATA][8] , \EXE_MEM_i[DMEM_DATA][7] , 
        \EXE_MEM_i[DMEM_DATA][6] , \EXE_MEM_i[DMEM_DATA][5] , 
        \EXE_MEM_i[DMEM_DATA][4] , \EXE_MEM_i[DMEM_DATA][3] , 
        \EXE_MEM_i[DMEM_DATA][2] , \EXE_MEM_i[DMEM_DATA][1] , 
        \EXE_MEM_i[DMEM_DATA][0] , \EXE_MEM_i[WRITE_REG][4] , 
        \EXE_MEM_i[WRITE_REG][3] , \EXE_MEM_i[WRITE_REG][2] , 
        \EXE_MEM_i[WRITE_REG][1] , \EXE_MEM_i[WRITE_REG][0] , 
        \EXE_MEM_i[MEMTOREG] , \EXE_MEM_i[REGWRITE] , \EXE_MEM_i[MEMWEN_N] }), 
    .EXE_MEM_o({\EXE_MEM_o[ALU_RES][31] , \EXE_MEM_o[ALU_RES][30] , 
        \EXE_MEM_o[ALU_RES][29] , \EXE_MEM_o[ALU_RES][28] , 
        \EXE_MEM_o[ALU_RES][27] , \EXE_MEM_o[ALU_RES][26] , 
        \EXE_MEM_o[ALU_RES][25] , \EXE_MEM_o[ALU_RES][24] , 
        \EXE_MEM_o[ALU_RES][23] , \EXE_MEM_o[ALU_RES][22] , 
        \EXE_MEM_o[ALU_RES][21] , \EXE_MEM_o[ALU_RES][20] , 
        \EXE_MEM_o[ALU_RES][19] , \EXE_MEM_o[ALU_RES][18] , 
        \EXE_MEM_o[ALU_RES][17] , \EXE_MEM_o[ALU_RES][16] , 
        \EXE_MEM_o[ALU_RES][15] , \EXE_MEM_o[ALU_RES][14] , 
        \EXE_MEM_o[ALU_RES][13] , \EXE_MEM_o[ALU_RES][12] , 
        \EXE_MEM_o[ALU_RES][11] , \EXE_MEM_o[ALU_RES][10] , 
        \EXE_MEM_o[ALU_RES][9] , \EXE_MEM_o[ALU_RES][8] , 
        \EXE_MEM_o[ALU_RES][7] , \EXE_MEM_o[ALU_RES][6] , 
        \EXE_MEM_o[ALU_RES][5] , \EXE_MEM_o[ALU_RES][4] , 
        \EXE_MEM_o[ALU_RES][3] , \EXE_MEM_o[ALU_RES][2] , 
        \EXE_MEM_o[ALU_RES][1] , \EXE_MEM_o[ALU_RES][0] , 
        \EXE_MEM_o[DMEM_DATA][31] , \EXE_MEM_o[DMEM_DATA][30] , 
        \EXE_MEM_o[DMEM_DATA][29] , \EXE_MEM_o[DMEM_DATA][28] , 
        \EXE_MEM_o[DMEM_DATA][27] , \EXE_MEM_o[DMEM_DATA][26] , 
        \EXE_MEM_o[DMEM_DATA][25] , \EXE_MEM_o[DMEM_DATA][24] , 
        \EXE_MEM_o[DMEM_DATA][23] , \EXE_MEM_o[DMEM_DATA][22] , 
        \EXE_MEM_o[DMEM_DATA][21] , \EXE_MEM_o[DMEM_DATA][20] , 
        \EXE_MEM_o[DMEM_DATA][19] , \EXE_MEM_o[DMEM_DATA][18] , 
        \EXE_MEM_o[DMEM_DATA][17] , \EXE_MEM_o[DMEM_DATA][16] , 
        \EXE_MEM_o[DMEM_DATA][15] , \EXE_MEM_o[DMEM_DATA][14] , 
        \EXE_MEM_o[DMEM_DATA][13] , \EXE_MEM_o[DMEM_DATA][12] , 
        \EXE_MEM_o[DMEM_DATA][11] , \EXE_MEM_o[DMEM_DATA][10] , 
        \EXE_MEM_o[DMEM_DATA][9] , \EXE_MEM_o[DMEM_DATA][8] , 
        \EXE_MEM_o[DMEM_DATA][7] , \EXE_MEM_o[DMEM_DATA][6] , 
        \EXE_MEM_o[DMEM_DATA][5] , \EXE_MEM_o[DMEM_DATA][4] , 
        \EXE_MEM_o[DMEM_DATA][3] , \EXE_MEM_o[DMEM_DATA][2] , 
        \EXE_MEM_o[DMEM_DATA][1] , \EXE_MEM_o[DMEM_DATA][0] , 
        \EXE_MEM_o[WRITE_REG][4] , \EXE_MEM_o[WRITE_REG][3] , 
        \EXE_MEM_o[WRITE_REG][2] , \EXE_MEM_o[WRITE_REG][1] , 
        \EXE_MEM_o[WRITE_REG][0] , \EXE_MEM_o[MEMTOREG] , 
        \EXE_MEM_o[REGWRITE] , \EXE_MEM_o[MEMWEN_N] }) );
  input clk, rst_n, halt_i, \EXE_MEM_i[ALU_RES][31] , \EXE_MEM_i[ALU_RES][30] ,
         \EXE_MEM_i[ALU_RES][29] , \EXE_MEM_i[ALU_RES][28] ,
         \EXE_MEM_i[ALU_RES][27] , \EXE_MEM_i[ALU_RES][26] ,
         \EXE_MEM_i[ALU_RES][25] , \EXE_MEM_i[ALU_RES][24] ,
         \EXE_MEM_i[ALU_RES][23] , \EXE_MEM_i[ALU_RES][22] ,
         \EXE_MEM_i[ALU_RES][21] , \EXE_MEM_i[ALU_RES][20] ,
         \EXE_MEM_i[ALU_RES][19] , \EXE_MEM_i[ALU_RES][18] ,
         \EXE_MEM_i[ALU_RES][17] , \EXE_MEM_i[ALU_RES][16] ,
         \EXE_MEM_i[ALU_RES][15] , \EXE_MEM_i[ALU_RES][14] ,
         \EXE_MEM_i[ALU_RES][13] , \EXE_MEM_i[ALU_RES][12] ,
         \EXE_MEM_i[ALU_RES][11] , \EXE_MEM_i[ALU_RES][10] ,
         \EXE_MEM_i[ALU_RES][9] , \EXE_MEM_i[ALU_RES][8] ,
         \EXE_MEM_i[ALU_RES][7] , \EXE_MEM_i[ALU_RES][6] ,
         \EXE_MEM_i[ALU_RES][5] , \EXE_MEM_i[ALU_RES][4] ,
         \EXE_MEM_i[ALU_RES][3] , \EXE_MEM_i[ALU_RES][2] ,
         \EXE_MEM_i[ALU_RES][1] , \EXE_MEM_i[ALU_RES][0] ,
         \EXE_MEM_i[DMEM_DATA][31] , \EXE_MEM_i[DMEM_DATA][30] ,
         \EXE_MEM_i[DMEM_DATA][29] , \EXE_MEM_i[DMEM_DATA][28] ,
         \EXE_MEM_i[DMEM_DATA][27] , \EXE_MEM_i[DMEM_DATA][26] ,
         \EXE_MEM_i[DMEM_DATA][25] , \EXE_MEM_i[DMEM_DATA][24] ,
         \EXE_MEM_i[DMEM_DATA][23] , \EXE_MEM_i[DMEM_DATA][22] ,
         \EXE_MEM_i[DMEM_DATA][21] , \EXE_MEM_i[DMEM_DATA][20] ,
         \EXE_MEM_i[DMEM_DATA][19] , \EXE_MEM_i[DMEM_DATA][18] ,
         \EXE_MEM_i[DMEM_DATA][17] , \EXE_MEM_i[DMEM_DATA][16] ,
         \EXE_MEM_i[DMEM_DATA][15] , \EXE_MEM_i[DMEM_DATA][14] ,
         \EXE_MEM_i[DMEM_DATA][13] , \EXE_MEM_i[DMEM_DATA][12] ,
         \EXE_MEM_i[DMEM_DATA][11] , \EXE_MEM_i[DMEM_DATA][10] ,
         \EXE_MEM_i[DMEM_DATA][9] , \EXE_MEM_i[DMEM_DATA][8] ,
         \EXE_MEM_i[DMEM_DATA][7] , \EXE_MEM_i[DMEM_DATA][6] ,
         \EXE_MEM_i[DMEM_DATA][5] , \EXE_MEM_i[DMEM_DATA][4] ,
         \EXE_MEM_i[DMEM_DATA][3] , \EXE_MEM_i[DMEM_DATA][2] ,
         \EXE_MEM_i[DMEM_DATA][1] , \EXE_MEM_i[DMEM_DATA][0] ,
         \EXE_MEM_i[WRITE_REG][4] , \EXE_MEM_i[WRITE_REG][3] ,
         \EXE_MEM_i[WRITE_REG][2] , \EXE_MEM_i[WRITE_REG][1] ,
         \EXE_MEM_i[WRITE_REG][0] , \EXE_MEM_i[MEMTOREG] ,
         \EXE_MEM_i[REGWRITE] , \EXE_MEM_i[MEMWEN_N] ;
  output \EXE_MEM_o[ALU_RES][31] , \EXE_MEM_o[ALU_RES][30] ,
         \EXE_MEM_o[ALU_RES][29] , \EXE_MEM_o[ALU_RES][28] ,
         \EXE_MEM_o[ALU_RES][27] , \EXE_MEM_o[ALU_RES][26] ,
         \EXE_MEM_o[ALU_RES][25] , \EXE_MEM_o[ALU_RES][24] ,
         \EXE_MEM_o[ALU_RES][23] , \EXE_MEM_o[ALU_RES][22] ,
         \EXE_MEM_o[ALU_RES][21] , \EXE_MEM_o[ALU_RES][20] ,
         \EXE_MEM_o[ALU_RES][19] , \EXE_MEM_o[ALU_RES][18] ,
         \EXE_MEM_o[ALU_RES][17] , \EXE_MEM_o[ALU_RES][16] ,
         \EXE_MEM_o[ALU_RES][15] , \EXE_MEM_o[ALU_RES][14] ,
         \EXE_MEM_o[ALU_RES][13] , \EXE_MEM_o[ALU_RES][12] ,
         \EXE_MEM_o[ALU_RES][11] , \EXE_MEM_o[ALU_RES][10] ,
         \EXE_MEM_o[ALU_RES][9] , \EXE_MEM_o[ALU_RES][8] ,
         \EXE_MEM_o[ALU_RES][7] , \EXE_MEM_o[ALU_RES][6] ,
         \EXE_MEM_o[ALU_RES][5] , \EXE_MEM_o[ALU_RES][4] ,
         \EXE_MEM_o[ALU_RES][3] , \EXE_MEM_o[ALU_RES][2] ,
         \EXE_MEM_o[ALU_RES][1] , \EXE_MEM_o[ALU_RES][0] ,
         \EXE_MEM_o[DMEM_DATA][31] , \EXE_MEM_o[DMEM_DATA][30] ,
         \EXE_MEM_o[DMEM_DATA][29] , \EXE_MEM_o[DMEM_DATA][28] ,
         \EXE_MEM_o[DMEM_DATA][27] , \EXE_MEM_o[DMEM_DATA][26] ,
         \EXE_MEM_o[DMEM_DATA][25] , \EXE_MEM_o[DMEM_DATA][24] ,
         \EXE_MEM_o[DMEM_DATA][23] , \EXE_MEM_o[DMEM_DATA][22] ,
         \EXE_MEM_o[DMEM_DATA][21] , \EXE_MEM_o[DMEM_DATA][20] ,
         \EXE_MEM_o[DMEM_DATA][19] , \EXE_MEM_o[DMEM_DATA][18] ,
         \EXE_MEM_o[DMEM_DATA][17] , \EXE_MEM_o[DMEM_DATA][16] ,
         \EXE_MEM_o[DMEM_DATA][15] , \EXE_MEM_o[DMEM_DATA][14] ,
         \EXE_MEM_o[DMEM_DATA][13] , \EXE_MEM_o[DMEM_DATA][12] ,
         \EXE_MEM_o[DMEM_DATA][11] , \EXE_MEM_o[DMEM_DATA][10] ,
         \EXE_MEM_o[DMEM_DATA][9] , \EXE_MEM_o[DMEM_DATA][8] ,
         \EXE_MEM_o[DMEM_DATA][7] , \EXE_MEM_o[DMEM_DATA][6] ,
         \EXE_MEM_o[DMEM_DATA][5] , \EXE_MEM_o[DMEM_DATA][4] ,
         \EXE_MEM_o[DMEM_DATA][3] , \EXE_MEM_o[DMEM_DATA][2] ,
         \EXE_MEM_o[DMEM_DATA][1] , \EXE_MEM_o[DMEM_DATA][0] ,
         \EXE_MEM_o[WRITE_REG][4] , \EXE_MEM_o[WRITE_REG][3] ,
         \EXE_MEM_o[WRITE_REG][2] , \EXE_MEM_o[WRITE_REG][1] ,
         \EXE_MEM_o[WRITE_REG][0] , \EXE_MEM_o[MEMTOREG] ,
         \EXE_MEM_o[REGWRITE] , \EXE_MEM_o[MEMWEN_N] ;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n1, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89;

  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][31]  ( .D(n73), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][31] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][30]  ( .D(n72), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][30] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][29]  ( .D(n71), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][29] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][28]  ( .D(n70), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][28] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][27]  ( .D(n69), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][27] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][26]  ( .D(n68), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][26] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][25]  ( .D(n67), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][25] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][24]  ( .D(n66), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][24] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][23]  ( .D(n65), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][23] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][22]  ( .D(n64), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][22] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][21]  ( .D(n63), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][21] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][20]  ( .D(n62), .CP(clk), .RN(n83), 
        .Q(\EXE_MEM_o[ALU_RES][20] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][19]  ( .D(n61), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][19] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][18]  ( .D(n60), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][18] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][17]  ( .D(n59), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][17] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][16]  ( .D(n58), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][16] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][15]  ( .D(n57), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][15] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][14]  ( .D(n56), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][14] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][13]  ( .D(n55), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][13] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][12]  ( .D(n54), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][12] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][11]  ( .D(n53), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][11] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][10]  ( .D(n52), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][10] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][9]  ( .D(n51), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][9] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][8]  ( .D(n50), .CP(clk), .RN(n84), 
        .Q(\EXE_MEM_o[ALU_RES][8] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][7]  ( .D(n49), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][7] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][6]  ( .D(n48), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][6] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][5]  ( .D(n47), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][5] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][4]  ( .D(n46), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][4] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][3]  ( .D(n45), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][3] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][2]  ( .D(n44), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][2] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][1]  ( .D(n43), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][1] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[ALU_RES][0]  ( .D(n42), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[ALU_RES][0] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][31]  ( .D(n41), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[DMEM_DATA][31] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][30]  ( .D(n40), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[DMEM_DATA][30] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][29]  ( .D(n39), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[DMEM_DATA][29] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][28]  ( .D(n38), .CP(clk), .RN(n85), 
        .Q(\EXE_MEM_o[DMEM_DATA][28] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][27]  ( .D(n37), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][27] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][26]  ( .D(n36), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][26] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][25]  ( .D(n35), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][25] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][24]  ( .D(n34), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][24] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][23]  ( .D(n33), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][23] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][22]  ( .D(n32), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][22] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][21]  ( .D(n31), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][21] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][20]  ( .D(n30), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][20] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][19]  ( .D(n29), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][19] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][18]  ( .D(n28), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][18] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][17]  ( .D(n27), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][17] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][16]  ( .D(n26), .CP(clk), .RN(n86), 
        .Q(\EXE_MEM_o[DMEM_DATA][16] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][15]  ( .D(n25), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][15] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][14]  ( .D(n24), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][14] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][13]  ( .D(n23), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][13] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][12]  ( .D(n22), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][12] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][11]  ( .D(n21), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][11] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][10]  ( .D(n20), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][10] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][9]  ( .D(n19), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][9] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][8]  ( .D(n18), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][8] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][7]  ( .D(n17), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][7] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][6]  ( .D(n16), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][6] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][5]  ( .D(n15), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][5] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][4]  ( .D(n14), .CP(clk), .RN(n87), 
        .Q(\EXE_MEM_o[DMEM_DATA][4] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][3]  ( .D(n13), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[DMEM_DATA][3] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][2]  ( .D(n12), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[DMEM_DATA][2] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][1]  ( .D(n11), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[DMEM_DATA][1] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[DMEM_DATA][0]  ( .D(n10), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[DMEM_DATA][0] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[WRITE_REG][4]  ( .D(n9), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[WRITE_REG][4] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[WRITE_REG][3]  ( .D(n8), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[WRITE_REG][3] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[WRITE_REG][2]  ( .D(n7), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[WRITE_REG][2] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[WRITE_REG][1]  ( .D(n6), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[WRITE_REG][1] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[WRITE_REG][0]  ( .D(n5), .CP(clk), .RN(n88), 
        .Q(\EXE_MEM_o[WRITE_REG][0] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[MEMTOREG]  ( .D(n4), .CP(clk), .RN(n88), .Q(
        \EXE_MEM_o[MEMTOREG] ) );
  HS65_LH_DFPRQX9 \exe_mem_c_reg[REGWRITE]  ( .D(n3), .CP(clk), .RN(n88), .Q(
        \EXE_MEM_o[REGWRITE] ) );
  HS65_LH_DFPSQX9 \exe_mem_c_reg[MEMWEN_N]  ( .D(n2), .CP(clk), .SN(n88), .Q(
        \EXE_MEM_o[MEMWEN_N] ) );
  HS65_LH_BFX9 U2 ( .A(n82), .Z(n87) );
  HS65_LH_BFX9 U3 ( .A(n82), .Z(n86) );
  HS65_LH_BFX9 U4 ( .A(n81), .Z(n85) );
  HS65_LH_BFX9 U5 ( .A(n81), .Z(n84) );
  HS65_LH_BFX9 U6 ( .A(n81), .Z(n83) );
  HS65_LH_BFX9 U7 ( .A(n82), .Z(n88) );
  HS65_LH_BFX9 U8 ( .A(rst_n), .Z(n82) );
  HS65_LH_BFX9 U9 ( .A(rst_n), .Z(n81) );
  HS65_LH_BFX9 U10 ( .A(n1), .Z(n75) );
  HS65_LH_BFX9 U11 ( .A(n1), .Z(n76) );
  HS65_LH_BFX9 U12 ( .A(n1), .Z(n77) );
  HS65_LH_BFX9 U13 ( .A(n74), .Z(n78) );
  HS65_LH_BFX9 U14 ( .A(n74), .Z(n79) );
  HS65_LH_BFX9 U15 ( .A(n74), .Z(n80) );
  HS65_LH_BFX9 U16 ( .A(n89), .Z(n1) );
  HS65_LH_BFX9 U17 ( .A(n89), .Z(n74) );
  HS65_LH_AO22X9 U18 ( .A(\EXE_MEM_o[ALU_RES][25] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][25] ), .D(n80), .Z(n67) );
  HS65_LH_AO22X9 U19 ( .A(\EXE_MEM_o[ALU_RES][26] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][26] ), .D(n80), .Z(n68) );
  HS65_LH_AO22X9 U20 ( .A(\EXE_MEM_o[ALU_RES][27] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][27] ), .D(n80), .Z(n69) );
  HS65_LH_AO22X9 U21 ( .A(\EXE_MEM_o[ALU_RES][29] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][29] ), .D(n80), .Z(n71) );
  HS65_LH_AO22X9 U22 ( .A(\EXE_MEM_o[ALU_RES][30] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][30] ), .D(n80), .Z(n72) );
  HS65_LH_AO22X9 U23 ( .A(\EXE_MEM_o[ALU_RES][28] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][28] ), .D(n80), .Z(n70) );
  HS65_LH_AO22X9 U24 ( .A(\EXE_MEM_o[ALU_RES][31] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][31] ), .D(n80), .Z(n73) );
  HS65_LH_AO22X9 U25 ( .A(\EXE_MEM_o[ALU_RES][21] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][21] ), .D(n80), .Z(n63) );
  HS65_LH_AO22X9 U26 ( .A(\EXE_MEM_o[ALU_RES][22] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][22] ), .D(n80), .Z(n64) );
  HS65_LH_AO22X9 U27 ( .A(\EXE_MEM_o[ALU_RES][23] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][23] ), .D(n80), .Z(n65) );
  HS65_LH_AO22X9 U28 ( .A(\EXE_MEM_o[ALU_RES][24] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][24] ), .D(n80), .Z(n66) );
  HS65_LH_AO22X9 U29 ( .A(\EXE_MEM_o[ALU_RES][17] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][17] ), .D(n79), .Z(n59) );
  HS65_LH_AO22X9 U30 ( .A(\EXE_MEM_o[ALU_RES][18] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][18] ), .D(n79), .Z(n60) );
  HS65_LH_AO22X9 U31 ( .A(\EXE_MEM_o[ALU_RES][19] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][19] ), .D(n79), .Z(n61) );
  HS65_LH_AO22X9 U32 ( .A(\EXE_MEM_o[ALU_RES][20] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][20] ), .D(n80), .Z(n62) );
  HS65_LH_AO22X9 U33 ( .A(\EXE_MEM_o[ALU_RES][0] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][0] ), .D(n78), .Z(n42) );
  HS65_LH_AO22X9 U34 ( .A(\EXE_MEM_o[ALU_RES][16] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][16] ), .D(n79), .Z(n58) );
  HS65_LH_AO22X9 U35 ( .A(\EXE_MEM_o[ALU_RES][9] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][9] ), .D(n79), .Z(n51) );
  HS65_LH_AO22X9 U36 ( .A(\EXE_MEM_o[ALU_RES][10] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][10] ), .D(n79), .Z(n52) );
  HS65_LH_AO22X9 U37 ( .A(\EXE_MEM_o[ALU_RES][11] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][11] ), .D(n79), .Z(n53) );
  HS65_LH_AO22X9 U38 ( .A(\EXE_MEM_o[ALU_RES][12] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][12] ), .D(n79), .Z(n54) );
  HS65_LH_AO22X9 U39 ( .A(\EXE_MEM_o[ALU_RES][13] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][13] ), .D(n79), .Z(n55) );
  HS65_LH_AO22X9 U40 ( .A(\EXE_MEM_o[ALU_RES][14] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][14] ), .D(n79), .Z(n56) );
  HS65_LH_AO22X9 U41 ( .A(\EXE_MEM_o[ALU_RES][15] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][15] ), .D(n79), .Z(n57) );
  HS65_LH_AO22X9 U42 ( .A(\EXE_MEM_o[ALU_RES][1] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][1] ), .D(n78), .Z(n43) );
  HS65_LH_AO22X9 U43 ( .A(\EXE_MEM_o[ALU_RES][4] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][4] ), .D(n78), .Z(n46) );
  HS65_LH_AO22X9 U44 ( .A(\EXE_MEM_o[ALU_RES][5] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][5] ), .D(n78), .Z(n47) );
  HS65_LH_AO22X9 U45 ( .A(\EXE_MEM_o[ALU_RES][6] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][6] ), .D(n78), .Z(n48) );
  HS65_LH_AO22X9 U46 ( .A(\EXE_MEM_o[ALU_RES][7] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][7] ), .D(n78), .Z(n49) );
  HS65_LH_AO22X9 U47 ( .A(\EXE_MEM_o[ALU_RES][8] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][8] ), .D(n79), .Z(n50) );
  HS65_LH_AO22X9 U48 ( .A(\EXE_MEM_o[ALU_RES][2] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][2] ), .D(n78), .Z(n44) );
  HS65_LH_AO22X9 U49 ( .A(\EXE_MEM_o[ALU_RES][3] ), .B(halt_i), .C(
        \EXE_MEM_i[ALU_RES][3] ), .D(n78), .Z(n45) );
  HS65_LH_AO22X9 U50 ( .A(\EXE_MEM_o[DMEM_DATA][9] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][9] ), .D(n76), .Z(n19) );
  HS65_LH_AO22X9 U51 ( .A(\EXE_MEM_o[DMEM_DATA][12] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][12] ), .D(n76), .Z(n22) );
  HS65_LH_AO22X9 U52 ( .A(\EXE_MEM_o[DMEM_DATA][13] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][13] ), .D(n76), .Z(n23) );
  HS65_LH_AO22X9 U53 ( .A(\EXE_MEM_o[DMEM_DATA][14] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][14] ), .D(n76), .Z(n24) );
  HS65_LH_AO22X9 U54 ( .A(\EXE_MEM_o[DMEM_DATA][15] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][15] ), .D(n76), .Z(n25) );
  HS65_LH_AO22X9 U55 ( .A(\EXE_MEM_o[DMEM_DATA][16] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][16] ), .D(n77), .Z(n26) );
  HS65_LH_AO22X9 U56 ( .A(\EXE_MEM_o[DMEM_DATA][17] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][17] ), .D(n77), .Z(n27) );
  HS65_LH_AO22X9 U57 ( .A(\EXE_MEM_o[DMEM_DATA][18] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][18] ), .D(n77), .Z(n28) );
  HS65_LH_AO22X9 U58 ( .A(\EXE_MEM_o[DMEM_DATA][19] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][19] ), .D(n77), .Z(n29) );
  HS65_LH_AO22X9 U59 ( .A(\EXE_MEM_o[DMEM_DATA][20] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][20] ), .D(n77), .Z(n30) );
  HS65_LH_AO22X9 U60 ( .A(\EXE_MEM_o[DMEM_DATA][21] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][21] ), .D(n77), .Z(n31) );
  HS65_LH_AO22X9 U61 ( .A(\EXE_MEM_o[DMEM_DATA][22] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][22] ), .D(n77), .Z(n32) );
  HS65_LH_AO22X9 U62 ( .A(\EXE_MEM_o[DMEM_DATA][23] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][23] ), .D(n77), .Z(n33) );
  HS65_LH_AO22X9 U63 ( .A(\EXE_MEM_o[DMEM_DATA][24] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][24] ), .D(n77), .Z(n34) );
  HS65_LH_AO22X9 U64 ( .A(\EXE_MEM_o[DMEM_DATA][25] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][25] ), .D(n77), .Z(n35) );
  HS65_LH_AO22X9 U65 ( .A(\EXE_MEM_o[DMEM_DATA][26] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][26] ), .D(n77), .Z(n36) );
  HS65_LH_AO22X9 U66 ( .A(\EXE_MEM_o[DMEM_DATA][27] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][27] ), .D(n77), .Z(n37) );
  HS65_LH_AO22X9 U67 ( .A(\EXE_MEM_o[DMEM_DATA][28] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][28] ), .D(n78), .Z(n38) );
  HS65_LH_AO22X9 U68 ( .A(\EXE_MEM_o[DMEM_DATA][29] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][29] ), .D(n78), .Z(n39) );
  HS65_LH_AO22X9 U69 ( .A(\EXE_MEM_o[DMEM_DATA][30] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][30] ), .D(n78), .Z(n40) );
  HS65_LH_AO22X9 U70 ( .A(\EXE_MEM_o[DMEM_DATA][31] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][31] ), .D(n78), .Z(n41) );
  HS65_LH_AO22X9 U71 ( .A(\EXE_MEM_o[DMEM_DATA][0] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][0] ), .D(n75), .Z(n10) );
  HS65_LH_AO22X9 U72 ( .A(\EXE_MEM_o[DMEM_DATA][1] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][1] ), .D(n75), .Z(n11) );
  HS65_LH_AO22X9 U73 ( .A(\EXE_MEM_o[DMEM_DATA][2] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][2] ), .D(n75), .Z(n12) );
  HS65_LH_AO22X9 U74 ( .A(\EXE_MEM_o[DMEM_DATA][3] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][3] ), .D(n75), .Z(n13) );
  HS65_LH_AO22X9 U75 ( .A(\EXE_MEM_o[DMEM_DATA][4] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][4] ), .D(n76), .Z(n14) );
  HS65_LH_AO22X9 U76 ( .A(\EXE_MEM_o[DMEM_DATA][5] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][5] ), .D(n76), .Z(n15) );
  HS65_LH_AO22X9 U77 ( .A(\EXE_MEM_o[DMEM_DATA][6] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][6] ), .D(n76), .Z(n16) );
  HS65_LH_AO22X9 U78 ( .A(\EXE_MEM_o[DMEM_DATA][7] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][7] ), .D(n76), .Z(n17) );
  HS65_LH_AO22X9 U79 ( .A(\EXE_MEM_o[DMEM_DATA][8] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][8] ), .D(n76), .Z(n18) );
  HS65_LH_AO22X9 U80 ( .A(\EXE_MEM_o[DMEM_DATA][10] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][10] ), .D(n76), .Z(n20) );
  HS65_LH_AO22X9 U81 ( .A(\EXE_MEM_o[DMEM_DATA][11] ), .B(halt_i), .C(
        \EXE_MEM_i[DMEM_DATA][11] ), .D(n76), .Z(n21) );
  HS65_LH_AO22X9 U82 ( .A(\EXE_MEM_o[WRITE_REG][0] ), .B(halt_i), .C(
        \EXE_MEM_i[WRITE_REG][0] ), .D(n75), .Z(n5) );
  HS65_LH_AO22X9 U83 ( .A(\EXE_MEM_o[WRITE_REG][1] ), .B(halt_i), .C(
        \EXE_MEM_i[WRITE_REG][1] ), .D(n75), .Z(n6) );
  HS65_LH_AO22X9 U84 ( .A(\EXE_MEM_o[WRITE_REG][2] ), .B(halt_i), .C(
        \EXE_MEM_i[WRITE_REG][2] ), .D(n75), .Z(n7) );
  HS65_LH_AO22X9 U85 ( .A(\EXE_MEM_o[WRITE_REG][3] ), .B(halt_i), .C(
        \EXE_MEM_i[WRITE_REG][3] ), .D(n75), .Z(n8) );
  HS65_LH_AO22X9 U86 ( .A(\EXE_MEM_o[WRITE_REG][4] ), .B(halt_i), .C(
        \EXE_MEM_i[WRITE_REG][4] ), .D(n75), .Z(n9) );
  HS65_LH_AO22X9 U87 ( .A(halt_i), .B(\EXE_MEM_o[MEMWEN_N] ), .C(
        \EXE_MEM_i[MEMWEN_N] ), .D(n75), .Z(n2) );
  HS65_LH_AO22X9 U88 ( .A(\EXE_MEM_o[REGWRITE] ), .B(halt_i), .C(
        \EXE_MEM_i[REGWRITE] ), .D(n75), .Z(n3) );
  HS65_LH_AO22X9 U89 ( .A(\EXE_MEM_o[MEMTOREG] ), .B(halt_i), .C(
        \EXE_MEM_i[MEMTOREG] ), .D(n75), .Z(n4) );
  HS65_LH_IVX9 U90 ( .A(halt_i), .Z(n89) );
endmodule


module mem_wb ( clk, rst_n, halt_i, .MEM_WB_i({\MEM_WB_i[ALU_RES][31] , 
        \MEM_WB_i[ALU_RES][30] , \MEM_WB_i[ALU_RES][29] , 
        \MEM_WB_i[ALU_RES][28] , \MEM_WB_i[ALU_RES][27] , 
        \MEM_WB_i[ALU_RES][26] , \MEM_WB_i[ALU_RES][25] , 
        \MEM_WB_i[ALU_RES][24] , \MEM_WB_i[ALU_RES][23] , 
        \MEM_WB_i[ALU_RES][22] , \MEM_WB_i[ALU_RES][21] , 
        \MEM_WB_i[ALU_RES][20] , \MEM_WB_i[ALU_RES][19] , 
        \MEM_WB_i[ALU_RES][18] , \MEM_WB_i[ALU_RES][17] , 
        \MEM_WB_i[ALU_RES][16] , \MEM_WB_i[ALU_RES][15] , 
        \MEM_WB_i[ALU_RES][14] , \MEM_WB_i[ALU_RES][13] , 
        \MEM_WB_i[ALU_RES][12] , \MEM_WB_i[ALU_RES][11] , 
        \MEM_WB_i[ALU_RES][10] , \MEM_WB_i[ALU_RES][9] , 
        \MEM_WB_i[ALU_RES][8] , \MEM_WB_i[ALU_RES][7] , \MEM_WB_i[ALU_RES][6] , 
        \MEM_WB_i[ALU_RES][5] , \MEM_WB_i[ALU_RES][4] , \MEM_WB_i[ALU_RES][3] , 
        \MEM_WB_i[ALU_RES][2] , \MEM_WB_i[ALU_RES][1] , \MEM_WB_i[ALU_RES][0] , 
        \MEM_WB_i[WRITE_REG][4] , \MEM_WB_i[WRITE_REG][3] , 
        \MEM_WB_i[WRITE_REG][2] , \MEM_WB_i[WRITE_REG][1] , 
        \MEM_WB_i[WRITE_REG][0] , \MEM_WB_i[MEMTOREG] , \MEM_WB_i[REGWRITE] }), 
    .MEM_WB_o({\MEM_WB_o[ALU_RES][31] , \MEM_WB_o[ALU_RES][30] , 
        \MEM_WB_o[ALU_RES][29] , \MEM_WB_o[ALU_RES][28] , 
        \MEM_WB_o[ALU_RES][27] , \MEM_WB_o[ALU_RES][26] , 
        \MEM_WB_o[ALU_RES][25] , \MEM_WB_o[ALU_RES][24] , 
        \MEM_WB_o[ALU_RES][23] , \MEM_WB_o[ALU_RES][22] , 
        \MEM_WB_o[ALU_RES][21] , \MEM_WB_o[ALU_RES][20] , 
        \MEM_WB_o[ALU_RES][19] , \MEM_WB_o[ALU_RES][18] , 
        \MEM_WB_o[ALU_RES][17] , \MEM_WB_o[ALU_RES][16] , 
        \MEM_WB_o[ALU_RES][15] , \MEM_WB_o[ALU_RES][14] , 
        \MEM_WB_o[ALU_RES][13] , \MEM_WB_o[ALU_RES][12] , 
        \MEM_WB_o[ALU_RES][11] , \MEM_WB_o[ALU_RES][10] , 
        \MEM_WB_o[ALU_RES][9] , \MEM_WB_o[ALU_RES][8] , \MEM_WB_o[ALU_RES][7] , 
        \MEM_WB_o[ALU_RES][6] , \MEM_WB_o[ALU_RES][5] , \MEM_WB_o[ALU_RES][4] , 
        \MEM_WB_o[ALU_RES][3] , \MEM_WB_o[ALU_RES][2] , \MEM_WB_o[ALU_RES][1] , 
        \MEM_WB_o[ALU_RES][0] , \MEM_WB_o[WRITE_REG][4] , 
        \MEM_WB_o[WRITE_REG][3] , \MEM_WB_o[WRITE_REG][2] , 
        \MEM_WB_o[WRITE_REG][1] , \MEM_WB_o[WRITE_REG][0] , 
        \MEM_WB_o[MEMTOREG] , \MEM_WB_o[REGWRITE] }) );
  input clk, rst_n, halt_i, \MEM_WB_i[ALU_RES][31] , \MEM_WB_i[ALU_RES][30] ,
         \MEM_WB_i[ALU_RES][29] , \MEM_WB_i[ALU_RES][28] ,
         \MEM_WB_i[ALU_RES][27] , \MEM_WB_i[ALU_RES][26] ,
         \MEM_WB_i[ALU_RES][25] , \MEM_WB_i[ALU_RES][24] ,
         \MEM_WB_i[ALU_RES][23] , \MEM_WB_i[ALU_RES][22] ,
         \MEM_WB_i[ALU_RES][21] , \MEM_WB_i[ALU_RES][20] ,
         \MEM_WB_i[ALU_RES][19] , \MEM_WB_i[ALU_RES][18] ,
         \MEM_WB_i[ALU_RES][17] , \MEM_WB_i[ALU_RES][16] ,
         \MEM_WB_i[ALU_RES][15] , \MEM_WB_i[ALU_RES][14] ,
         \MEM_WB_i[ALU_RES][13] , \MEM_WB_i[ALU_RES][12] ,
         \MEM_WB_i[ALU_RES][11] , \MEM_WB_i[ALU_RES][10] ,
         \MEM_WB_i[ALU_RES][9] , \MEM_WB_i[ALU_RES][8] ,
         \MEM_WB_i[ALU_RES][7] , \MEM_WB_i[ALU_RES][6] ,
         \MEM_WB_i[ALU_RES][5] , \MEM_WB_i[ALU_RES][4] ,
         \MEM_WB_i[ALU_RES][3] , \MEM_WB_i[ALU_RES][2] ,
         \MEM_WB_i[ALU_RES][1] , \MEM_WB_i[ALU_RES][0] ,
         \MEM_WB_i[WRITE_REG][4] , \MEM_WB_i[WRITE_REG][3] ,
         \MEM_WB_i[WRITE_REG][2] , \MEM_WB_i[WRITE_REG][1] ,
         \MEM_WB_i[WRITE_REG][0] , \MEM_WB_i[MEMTOREG] , \MEM_WB_i[REGWRITE] ;
  output \MEM_WB_o[ALU_RES][31] , \MEM_WB_o[ALU_RES][30] ,
         \MEM_WB_o[ALU_RES][29] , \MEM_WB_o[ALU_RES][28] ,
         \MEM_WB_o[ALU_RES][27] , \MEM_WB_o[ALU_RES][26] ,
         \MEM_WB_o[ALU_RES][25] , \MEM_WB_o[ALU_RES][24] ,
         \MEM_WB_o[ALU_RES][23] , \MEM_WB_o[ALU_RES][22] ,
         \MEM_WB_o[ALU_RES][21] , \MEM_WB_o[ALU_RES][20] ,
         \MEM_WB_o[ALU_RES][19] , \MEM_WB_o[ALU_RES][18] ,
         \MEM_WB_o[ALU_RES][17] , \MEM_WB_o[ALU_RES][16] ,
         \MEM_WB_o[ALU_RES][15] , \MEM_WB_o[ALU_RES][14] ,
         \MEM_WB_o[ALU_RES][13] , \MEM_WB_o[ALU_RES][12] ,
         \MEM_WB_o[ALU_RES][11] , \MEM_WB_o[ALU_RES][10] ,
         \MEM_WB_o[ALU_RES][9] , \MEM_WB_o[ALU_RES][8] ,
         \MEM_WB_o[ALU_RES][7] , \MEM_WB_o[ALU_RES][6] ,
         \MEM_WB_o[ALU_RES][5] , \MEM_WB_o[ALU_RES][4] ,
         \MEM_WB_o[ALU_RES][3] , \MEM_WB_o[ALU_RES][2] ,
         \MEM_WB_o[ALU_RES][1] , \MEM_WB_o[ALU_RES][0] ,
         \MEM_WB_o[WRITE_REG][4] , \MEM_WB_o[WRITE_REG][3] ,
         \MEM_WB_o[WRITE_REG][2] , \MEM_WB_o[WRITE_REG][1] ,
         \MEM_WB_o[WRITE_REG][0] , \MEM_WB_o[MEMTOREG] , \MEM_WB_o[REGWRITE] ;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n1, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52;

  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][31]  ( .D(n40), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][31] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][30]  ( .D(n39), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][30] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][29]  ( .D(n38), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][29] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][28]  ( .D(n37), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][28] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][27]  ( .D(n36), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][27] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][26]  ( .D(n35), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][26] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][25]  ( .D(n34), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][25] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][24]  ( .D(n33), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][24] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][23]  ( .D(n32), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][23] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][22]  ( .D(n31), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][22] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][21]  ( .D(n30), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][21] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][20]  ( .D(n29), .CP(clk), .RN(n48), 
        .Q(\MEM_WB_o[ALU_RES][20] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][19]  ( .D(n28), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][19] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][18]  ( .D(n27), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][18] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][17]  ( .D(n26), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][17] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][16]  ( .D(n25), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][16] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][15]  ( .D(n24), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][15] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][14]  ( .D(n23), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][14] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][13]  ( .D(n22), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][13] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][12]  ( .D(n21), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][12] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][11]  ( .D(n20), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][11] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][10]  ( .D(n19), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][10] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][9]  ( .D(n18), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][9] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][8]  ( .D(n17), .CP(clk), .RN(n49), 
        .Q(\MEM_WB_o[ALU_RES][8] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][7]  ( .D(n16), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][7] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][6]  ( .D(n15), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][6] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][5]  ( .D(n14), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][5] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][4]  ( .D(n13), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][4] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][3]  ( .D(n12), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][3] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][2]  ( .D(n11), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][2] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][1]  ( .D(n10), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[ALU_RES][1] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[ALU_RES][0]  ( .D(n9), .CP(clk), .RN(n50), .Q(
        \MEM_WB_o[ALU_RES][0] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[WRITE_REG][4]  ( .D(n8), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[WRITE_REG][4] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[WRITE_REG][3]  ( .D(n7), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[WRITE_REG][3] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[WRITE_REG][2]  ( .D(n6), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[WRITE_REG][2] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[WRITE_REG][1]  ( .D(n5), .CP(clk), .RN(n50), 
        .Q(\MEM_WB_o[WRITE_REG][1] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[WRITE_REG][0]  ( .D(n4), .CP(clk), .RN(n51), 
        .Q(\MEM_WB_o[WRITE_REG][0] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[MEMTOREG]  ( .D(n3), .CP(clk), .RN(n51), .Q(
        \MEM_WB_o[MEMTOREG] ) );
  HS65_LH_DFPRQX9 \mem_wb_c_reg[REGWRITE]  ( .D(n2), .CP(clk), .RN(n51), .Q(
        \MEM_WB_o[REGWRITE] ) );
  HS65_LH_BFX9 U2 ( .A(n47), .Z(n50) );
  HS65_LH_BFX9 U3 ( .A(n46), .Z(n49) );
  HS65_LH_BFX9 U4 ( .A(n46), .Z(n48) );
  HS65_LH_BFX9 U5 ( .A(n47), .Z(n51) );
  HS65_LH_BFX9 U6 ( .A(rst_n), .Z(n47) );
  HS65_LH_BFX9 U7 ( .A(rst_n), .Z(n46) );
  HS65_LH_BFX9 U8 ( .A(n1), .Z(n42) );
  HS65_LH_BFX9 U9 ( .A(n1), .Z(n43) );
  HS65_LH_BFX9 U10 ( .A(n41), .Z(n44) );
  HS65_LH_BFX9 U11 ( .A(n41), .Z(n45) );
  HS65_LH_BFX9 U12 ( .A(n52), .Z(n1) );
  HS65_LH_BFX9 U13 ( .A(n52), .Z(n41) );
  HS65_LH_AO22X9 U14 ( .A(\MEM_WB_o[WRITE_REG][2] ), .B(halt_i), .C(
        \MEM_WB_i[WRITE_REG][2] ), .D(n42), .Z(n6) );
  HS65_LH_AO22X9 U15 ( .A(\MEM_WB_o[WRITE_REG][4] ), .B(halt_i), .C(
        \MEM_WB_i[WRITE_REG][4] ), .D(n42), .Z(n8) );
  HS65_LH_AO22X9 U16 ( .A(\MEM_WB_o[WRITE_REG][0] ), .B(halt_i), .C(
        \MEM_WB_i[WRITE_REG][0] ), .D(n42), .Z(n4) );
  HS65_LH_AO22X9 U17 ( .A(\MEM_WB_o[WRITE_REG][3] ), .B(halt_i), .C(
        \MEM_WB_i[WRITE_REG][3] ), .D(n42), .Z(n7) );
  HS65_LH_AO22X9 U18 ( .A(\MEM_WB_o[WRITE_REG][1] ), .B(halt_i), .C(
        \MEM_WB_i[WRITE_REG][1] ), .D(n42), .Z(n5) );
  HS65_LH_AO22X9 U19 ( .A(\MEM_WB_o[ALU_RES][0] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][0] ), .D(n42), .Z(n9) );
  HS65_LH_AO22X9 U20 ( .A(\MEM_WB_o[ALU_RES][1] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][1] ), .D(n42), .Z(n10) );
  HS65_LH_AO22X9 U21 ( .A(\MEM_WB_o[ALU_RES][2] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][2] ), .D(n42), .Z(n11) );
  HS65_LH_AO22X9 U22 ( .A(\MEM_WB_o[ALU_RES][3] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][3] ), .D(n42), .Z(n12) );
  HS65_LH_AO22X9 U23 ( .A(\MEM_WB_o[ALU_RES][4] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][4] ), .D(n42), .Z(n13) );
  HS65_LH_AO22X9 U24 ( .A(\MEM_WB_o[ALU_RES][5] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][5] ), .D(n43), .Z(n14) );
  HS65_LH_AO22X9 U25 ( .A(\MEM_WB_o[ALU_RES][6] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][6] ), .D(n43), .Z(n15) );
  HS65_LH_AO22X9 U26 ( .A(\MEM_WB_o[ALU_RES][7] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][7] ), .D(n43), .Z(n16) );
  HS65_LH_AO22X9 U27 ( .A(\MEM_WB_o[ALU_RES][8] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][8] ), .D(n43), .Z(n17) );
  HS65_LH_AO22X9 U28 ( .A(\MEM_WB_o[ALU_RES][9] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][9] ), .D(n43), .Z(n18) );
  HS65_LH_AO22X9 U29 ( .A(\MEM_WB_o[ALU_RES][10] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][10] ), .D(n43), .Z(n19) );
  HS65_LH_AO22X9 U30 ( .A(\MEM_WB_o[ALU_RES][11] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][11] ), .D(n43), .Z(n20) );
  HS65_LH_AO22X9 U31 ( .A(halt_i), .B(\MEM_WB_o[REGWRITE] ), .C(
        \MEM_WB_i[REGWRITE] ), .D(n42), .Z(n2) );
  HS65_LH_AO22X9 U32 ( .A(\MEM_WB_o[ALU_RES][12] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][12] ), .D(n43), .Z(n21) );
  HS65_LH_AO22X9 U33 ( .A(\MEM_WB_o[ALU_RES][13] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][13] ), .D(n43), .Z(n22) );
  HS65_LH_AO22X9 U34 ( .A(\MEM_WB_o[ALU_RES][14] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][14] ), .D(n43), .Z(n23) );
  HS65_LH_AO22X9 U35 ( .A(\MEM_WB_o[ALU_RES][15] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][15] ), .D(n43), .Z(n24) );
  HS65_LH_AO22X9 U36 ( .A(\MEM_WB_o[ALU_RES][16] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][16] ), .D(n43), .Z(n25) );
  HS65_LH_AO22X9 U37 ( .A(\MEM_WB_o[ALU_RES][17] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][17] ), .D(n44), .Z(n26) );
  HS65_LH_AO22X9 U38 ( .A(\MEM_WB_o[ALU_RES][18] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][18] ), .D(n44), .Z(n27) );
  HS65_LH_AO22X9 U39 ( .A(\MEM_WB_o[ALU_RES][19] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][19] ), .D(n44), .Z(n28) );
  HS65_LH_AO22X9 U40 ( .A(\MEM_WB_o[ALU_RES][20] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][20] ), .D(n44), .Z(n29) );
  HS65_LH_AO22X9 U41 ( .A(\MEM_WB_o[ALU_RES][21] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][21] ), .D(n44), .Z(n30) );
  HS65_LH_AO22X9 U42 ( .A(\MEM_WB_o[ALU_RES][22] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][22] ), .D(n44), .Z(n31) );
  HS65_LH_AO22X9 U43 ( .A(\MEM_WB_o[ALU_RES][23] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][23] ), .D(n44), .Z(n32) );
  HS65_LH_AO22X9 U44 ( .A(\MEM_WB_o[ALU_RES][24] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][24] ), .D(n44), .Z(n33) );
  HS65_LH_AO22X9 U45 ( .A(\MEM_WB_o[ALU_RES][25] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][25] ), .D(n44), .Z(n34) );
  HS65_LH_AO22X9 U46 ( .A(\MEM_WB_o[ALU_RES][26] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][26] ), .D(n44), .Z(n35) );
  HS65_LH_AO22X9 U47 ( .A(\MEM_WB_o[ALU_RES][27] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][27] ), .D(n44), .Z(n36) );
  HS65_LH_AO22X9 U48 ( .A(\MEM_WB_o[ALU_RES][28] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][28] ), .D(n44), .Z(n37) );
  HS65_LH_AO22X9 U49 ( .A(\MEM_WB_o[ALU_RES][29] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][29] ), .D(n45), .Z(n38) );
  HS65_LH_AO22X9 U50 ( .A(\MEM_WB_o[ALU_RES][30] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][30] ), .D(n45), .Z(n39) );
  HS65_LH_AO22X9 U51 ( .A(\MEM_WB_o[ALU_RES][31] ), .B(halt_i), .C(
        \MEM_WB_i[ALU_RES][31] ), .D(n45), .Z(n40) );
  HS65_LH_AO22X9 U52 ( .A(\MEM_WB_o[MEMTOREG] ), .B(halt_i), .C(
        \MEM_WB_i[MEMTOREG] ), .D(n42), .Z(n3) );
  HS65_LH_IVX9 U53 ( .A(halt_i), .Z(n52) );
endmodule


module mini_mips_pipeline ( clk, rst_n, .mini_mips_i({
        \mini_mips_i[DMEM_DATA][31] , \mini_mips_i[DMEM_DATA][30] , 
        \mini_mips_i[DMEM_DATA][29] , \mini_mips_i[DMEM_DATA][28] , 
        \mini_mips_i[DMEM_DATA][27] , \mini_mips_i[DMEM_DATA][26] , 
        \mini_mips_i[DMEM_DATA][25] , \mini_mips_i[DMEM_DATA][24] , 
        \mini_mips_i[DMEM_DATA][23] , \mini_mips_i[DMEM_DATA][22] , 
        \mini_mips_i[DMEM_DATA][21] , \mini_mips_i[DMEM_DATA][20] , 
        \mini_mips_i[DMEM_DATA][19] , \mini_mips_i[DMEM_DATA][18] , 
        \mini_mips_i[DMEM_DATA][17] , \mini_mips_i[DMEM_DATA][16] , 
        \mini_mips_i[DMEM_DATA][15] , \mini_mips_i[DMEM_DATA][14] , 
        \mini_mips_i[DMEM_DATA][13] , \mini_mips_i[DMEM_DATA][12] , 
        \mini_mips_i[DMEM_DATA][11] , \mini_mips_i[DMEM_DATA][10] , 
        \mini_mips_i[DMEM_DATA][9] , \mini_mips_i[DMEM_DATA][8] , 
        \mini_mips_i[DMEM_DATA][7] , \mini_mips_i[DMEM_DATA][6] , 
        \mini_mips_i[DMEM_DATA][5] , \mini_mips_i[DMEM_DATA][4] , 
        \mini_mips_i[DMEM_DATA][3] , \mini_mips_i[DMEM_DATA][2] , 
        \mini_mips_i[DMEM_DATA][1] , \mini_mips_i[DMEM_DATA][0] , 
        \mini_mips_i[IMEM_DATA][31] , \mini_mips_i[IMEM_DATA][30] , 
        \mini_mips_i[IMEM_DATA][29] , \mini_mips_i[IMEM_DATA][28] , 
        \mini_mips_i[IMEM_DATA][27] , \mini_mips_i[IMEM_DATA][26] , 
        \mini_mips_i[IMEM_DATA][25] , \mini_mips_i[IMEM_DATA][24] , 
        \mini_mips_i[IMEM_DATA][23] , \mini_mips_i[IMEM_DATA][22] , 
        \mini_mips_i[IMEM_DATA][21] , \mini_mips_i[IMEM_DATA][20] , 
        \mini_mips_i[IMEM_DATA][19] , \mini_mips_i[IMEM_DATA][18] , 
        \mini_mips_i[IMEM_DATA][17] , \mini_mips_i[IMEM_DATA][16] , 
        \mini_mips_i[IMEM_DATA][15] , \mini_mips_i[IMEM_DATA][14] , 
        \mini_mips_i[IMEM_DATA][13] , \mini_mips_i[IMEM_DATA][12] , 
        \mini_mips_i[IMEM_DATA][11] , \mini_mips_i[IMEM_DATA][10] , 
        \mini_mips_i[IMEM_DATA][9] , \mini_mips_i[IMEM_DATA][8] , 
        \mini_mips_i[IMEM_DATA][7] , \mini_mips_i[IMEM_DATA][6] , 
        \mini_mips_i[IMEM_DATA][5] , \mini_mips_i[IMEM_DATA][4] , 
        \mini_mips_i[IMEM_DATA][3] , \mini_mips_i[IMEM_DATA][2] , 
        \mini_mips_i[IMEM_DATA][1] , \mini_mips_i[IMEM_DATA][0] }), 
    .mini_mips_o({\mini_mips_o[DMEM_ADDR][11] , \mini_mips_o[DMEM_ADDR][10] , 
        \mini_mips_o[DMEM_ADDR][9] , \mini_mips_o[DMEM_ADDR][8] , 
        \mini_mips_o[DMEM_ADDR][7] , \mini_mips_o[DMEM_ADDR][6] , 
        \mini_mips_o[DMEM_ADDR][5] , \mini_mips_o[DMEM_ADDR][4] , 
        \mini_mips_o[DMEM_ADDR][3] , \mini_mips_o[DMEM_ADDR][2] , 
        \mini_mips_o[DMEM_ADDR][1] , \mini_mips_o[DMEM_ADDR][0] , 
        \mini_mips_o[DMEM_DATA][31] , \mini_mips_o[DMEM_DATA][30] , 
        \mini_mips_o[DMEM_DATA][29] , \mini_mips_o[DMEM_DATA][28] , 
        \mini_mips_o[DMEM_DATA][27] , \mini_mips_o[DMEM_DATA][26] , 
        \mini_mips_o[DMEM_DATA][25] , \mini_mips_o[DMEM_DATA][24] , 
        \mini_mips_o[DMEM_DATA][23] , \mini_mips_o[DMEM_DATA][22] , 
        \mini_mips_o[DMEM_DATA][21] , \mini_mips_o[DMEM_DATA][20] , 
        \mini_mips_o[DMEM_DATA][19] , \mini_mips_o[DMEM_DATA][18] , 
        \mini_mips_o[DMEM_DATA][17] , \mini_mips_o[DMEM_DATA][16] , 
        \mini_mips_o[DMEM_DATA][15] , \mini_mips_o[DMEM_DATA][14] , 
        \mini_mips_o[DMEM_DATA][13] , \mini_mips_o[DMEM_DATA][12] , 
        \mini_mips_o[DMEM_DATA][11] , \mini_mips_o[DMEM_DATA][10] , 
        \mini_mips_o[DMEM_DATA][9] , \mini_mips_o[DMEM_DATA][8] , 
        \mini_mips_o[DMEM_DATA][7] , \mini_mips_o[DMEM_DATA][6] , 
        \mini_mips_o[DMEM_DATA][5] , \mini_mips_o[DMEM_DATA][4] , 
        \mini_mips_o[DMEM_DATA][3] , \mini_mips_o[DMEM_DATA][2] , 
        \mini_mips_o[DMEM_DATA][1] , \mini_mips_o[DMEM_DATA][0] , 
        \mini_mips_o[IMEM_ADDR][11] , \mini_mips_o[IMEM_ADDR][10] , 
        \mini_mips_o[IMEM_ADDR][9] , \mini_mips_o[IMEM_ADDR][8] , 
        \mini_mips_o[IMEM_ADDR][7] , \mini_mips_o[IMEM_ADDR][6] , 
        \mini_mips_o[IMEM_ADDR][5] , \mini_mips_o[IMEM_ADDR][4] , 
        \mini_mips_o[IMEM_ADDR][3] , \mini_mips_o[IMEM_ADDR][2] , 
        \mini_mips_o[IMEM_ADDR][1] , \mini_mips_o[IMEM_ADDR][0] , 
        \mini_mips_o[DMEM_WEN_N] }) );
  input clk, rst_n, \mini_mips_i[DMEM_DATA][31] , \mini_mips_i[DMEM_DATA][30] ,
         \mini_mips_i[DMEM_DATA][29] , \mini_mips_i[DMEM_DATA][28] ,
         \mini_mips_i[DMEM_DATA][27] , \mini_mips_i[DMEM_DATA][26] ,
         \mini_mips_i[DMEM_DATA][25] , \mini_mips_i[DMEM_DATA][24] ,
         \mini_mips_i[DMEM_DATA][23] , \mini_mips_i[DMEM_DATA][22] ,
         \mini_mips_i[DMEM_DATA][21] , \mini_mips_i[DMEM_DATA][20] ,
         \mini_mips_i[DMEM_DATA][19] , \mini_mips_i[DMEM_DATA][18] ,
         \mini_mips_i[DMEM_DATA][17] , \mini_mips_i[DMEM_DATA][16] ,
         \mini_mips_i[DMEM_DATA][15] , \mini_mips_i[DMEM_DATA][14] ,
         \mini_mips_i[DMEM_DATA][13] , \mini_mips_i[DMEM_DATA][12] ,
         \mini_mips_i[DMEM_DATA][11] , \mini_mips_i[DMEM_DATA][10] ,
         \mini_mips_i[DMEM_DATA][9] , \mini_mips_i[DMEM_DATA][8] ,
         \mini_mips_i[DMEM_DATA][7] , \mini_mips_i[DMEM_DATA][6] ,
         \mini_mips_i[DMEM_DATA][5] , \mini_mips_i[DMEM_DATA][4] ,
         \mini_mips_i[DMEM_DATA][3] , \mini_mips_i[DMEM_DATA][2] ,
         \mini_mips_i[DMEM_DATA][1] , \mini_mips_i[DMEM_DATA][0] ,
         \mini_mips_i[IMEM_DATA][31] , \mini_mips_i[IMEM_DATA][30] ,
         \mini_mips_i[IMEM_DATA][29] , \mini_mips_i[IMEM_DATA][28] ,
         \mini_mips_i[IMEM_DATA][27] , \mini_mips_i[IMEM_DATA][26] ,
         \mini_mips_i[IMEM_DATA][25] , \mini_mips_i[IMEM_DATA][24] ,
         \mini_mips_i[IMEM_DATA][23] , \mini_mips_i[IMEM_DATA][22] ,
         \mini_mips_i[IMEM_DATA][21] , \mini_mips_i[IMEM_DATA][20] ,
         \mini_mips_i[IMEM_DATA][19] , \mini_mips_i[IMEM_DATA][18] ,
         \mini_mips_i[IMEM_DATA][17] , \mini_mips_i[IMEM_DATA][16] ,
         \mini_mips_i[IMEM_DATA][15] , \mini_mips_i[IMEM_DATA][14] ,
         \mini_mips_i[IMEM_DATA][13] , \mini_mips_i[IMEM_DATA][12] ,
         \mini_mips_i[IMEM_DATA][11] , \mini_mips_i[IMEM_DATA][10] ,
         \mini_mips_i[IMEM_DATA][9] , \mini_mips_i[IMEM_DATA][8] ,
         \mini_mips_i[IMEM_DATA][7] , \mini_mips_i[IMEM_DATA][6] ,
         \mini_mips_i[IMEM_DATA][5] , \mini_mips_i[IMEM_DATA][4] ,
         \mini_mips_i[IMEM_DATA][3] , \mini_mips_i[IMEM_DATA][2] ,
         \mini_mips_i[IMEM_DATA][1] , \mini_mips_i[IMEM_DATA][0] ;
  output \mini_mips_o[DMEM_ADDR][11] , \mini_mips_o[DMEM_ADDR][10] ,
         \mini_mips_o[DMEM_ADDR][9] , \mini_mips_o[DMEM_ADDR][8] ,
         \mini_mips_o[DMEM_ADDR][7] , \mini_mips_o[DMEM_ADDR][6] ,
         \mini_mips_o[DMEM_ADDR][5] , \mini_mips_o[DMEM_ADDR][4] ,
         \mini_mips_o[DMEM_ADDR][3] , \mini_mips_o[DMEM_ADDR][2] ,
         \mini_mips_o[DMEM_ADDR][1] , \mini_mips_o[DMEM_ADDR][0] ,
         \mini_mips_o[DMEM_DATA][31] , \mini_mips_o[DMEM_DATA][30] ,
         \mini_mips_o[DMEM_DATA][29] , \mini_mips_o[DMEM_DATA][28] ,
         \mini_mips_o[DMEM_DATA][27] , \mini_mips_o[DMEM_DATA][26] ,
         \mini_mips_o[DMEM_DATA][25] , \mini_mips_o[DMEM_DATA][24] ,
         \mini_mips_o[DMEM_DATA][23] , \mini_mips_o[DMEM_DATA][22] ,
         \mini_mips_o[DMEM_DATA][21] , \mini_mips_o[DMEM_DATA][20] ,
         \mini_mips_o[DMEM_DATA][19] , \mini_mips_o[DMEM_DATA][18] ,
         \mini_mips_o[DMEM_DATA][17] , \mini_mips_o[DMEM_DATA][16] ,
         \mini_mips_o[DMEM_DATA][15] , \mini_mips_o[DMEM_DATA][14] ,
         \mini_mips_o[DMEM_DATA][13] , \mini_mips_o[DMEM_DATA][12] ,
         \mini_mips_o[DMEM_DATA][11] , \mini_mips_o[DMEM_DATA][10] ,
         \mini_mips_o[DMEM_DATA][9] , \mini_mips_o[DMEM_DATA][8] ,
         \mini_mips_o[DMEM_DATA][7] , \mini_mips_o[DMEM_DATA][6] ,
         \mini_mips_o[DMEM_DATA][5] , \mini_mips_o[DMEM_DATA][4] ,
         \mini_mips_o[DMEM_DATA][3] , \mini_mips_o[DMEM_DATA][2] ,
         \mini_mips_o[DMEM_DATA][1] , \mini_mips_o[DMEM_DATA][0] ,
         \mini_mips_o[IMEM_ADDR][11] , \mini_mips_o[IMEM_ADDR][10] ,
         \mini_mips_o[IMEM_ADDR][9] , \mini_mips_o[IMEM_ADDR][8] ,
         \mini_mips_o[IMEM_ADDR][7] , \mini_mips_o[IMEM_ADDR][6] ,
         \mini_mips_o[IMEM_ADDR][5] , \mini_mips_o[IMEM_ADDR][4] ,
         \mini_mips_o[IMEM_ADDR][3] , \mini_mips_o[IMEM_ADDR][2] ,
         \mini_mips_o[IMEM_ADDR][1] , \mini_mips_o[IMEM_ADDR][0] ,
         \mini_mips_o[DMEM_WEN_N] ;
  wire   s_if_PCSrc, s_exe_out_memtoReg_p, s_exe_out_regWrite_p,
         s_exe_out_memWen_n_p, s_mem_out_memtoReg_p, s_mem_out_regWrite_p,
         s_wb_in_memtoReg_p, s_ctrl_out_RegDst_p, s_ctrl_out_ALUsrc_B_p,
         s_ctrl_out_memtoReg_p, s_ctrl_out_regWrite_p, s_ctrl_out_memWen_n_p,
         s_regfile_forward_A, s_regfile_forward_B, s_wb_in_regWrite_p,
         s_exe_in_ALUsrc_B_p, s_exe_in_RegDst_p, n4, n6, n7, n9, n1, n2, n3,
         n5, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37;
  wire   [11:0] s_id_out_pc_plus1_p;
  wire   [4:0] s_mem_out_write_reg_p;
  wire   [31:12] s_mem_out_alu_res_p;
  wire   [31:0] s_writeback_data;
  wire   [31:0] s_wb_in_alu_res_p;
  wire   [1:0] s_forward_A;
  wire   [31:0] s_src_a;
  wire   [31:0] s_exe_in_regA_p;
  wire   [1:0] s_forward_B;
  wire   [31:0] s_src_b;
  wire   [31:0] s_exe_in_regB_p;
  wire   [5:0] s_id_ctrl_opcode;
  wire   [3:0] s_ctrl_out_cALU_OP_p;
  wire   [11:0] s_exe_if_branch_pc;
  wire   [11:0] s_if_out_pc_plus1_p;
  wire   [4:0] s_wb_in_write_reg_p;
  wire   [31:0] s_id_out_regA_p;
  wire   [31:0] s_id_out_regB_p;
  wire   [4:0] s_id_out_RS_p;
  wire   [4:0] s_id_out_RT_p;
  wire   [4:0] s_id_out_RD_p;
  wire   [4:0] s_id_out_shamt_p;
  wire   [5:0] s_id_out_funct_p;
  wire   [31:0] s_id_out_sign_extend_p;
  wire   [4:0] s_exe_in_shamt_p;
  wire   [5:0] s_exe_in_funct_p;
  wire   [31:0] s_exe_in_sign_extend_p;
  wire   [11:0] s_exe_in_pc_plus1_p;
  wire   [4:0] s_exe_in_RS_p;
  wire   [4:0] s_exe_in_RT_p;
  wire   [4:0] s_exe_in_RD_p;
  wire   [3:0] s_exe_in_cALU_OP_p;
  wire   [31:0] s_exe_out_alu_res_p;
  wire   [4:0] s_exe_out_write_reg_p;
  wire   [31:0] s_exe_out_dmem_data_p;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  controller ctrl_inst ( .ctrl_i(s_id_ctrl_opcode), .ctrl_o({
        s_ctrl_out_RegDst_p, s_ctrl_out_ALUsrc_B_p, s_ctrl_out_memtoReg_p, 
        s_ctrl_out_regWrite_p, s_ctrl_out_memWen_n_p, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, s_ctrl_out_cALU_OP_p[2:0]}) );
  if_top if_top_inst ( .clk(clk), .rst_n(n35), .if_top_i({1'b0, 
        s_exe_if_branch_pc, s_if_PCSrc}), .if_top_o({
        \mini_mips_o[IMEM_ADDR][11] , \mini_mips_o[IMEM_ADDR][10] , 
        \mini_mips_o[IMEM_ADDR][9] , \mini_mips_o[IMEM_ADDR][8] , 
        \mini_mips_o[IMEM_ADDR][7] , \mini_mips_o[IMEM_ADDR][6] , 
        \mini_mips_o[IMEM_ADDR][5] , \mini_mips_o[IMEM_ADDR][4] , 
        \mini_mips_o[IMEM_ADDR][3] , \mini_mips_o[IMEM_ADDR][2] , 
        \mini_mips_o[IMEM_ADDR][1] , \mini_mips_o[IMEM_ADDR][0] , 
        s_if_out_pc_plus1_p}) );
  if_id if_id_inst ( .clk(clk), .rst_n(n34), .halt_i(1'b0), .IF_ID_i(
        s_if_out_pc_plus1_p), .IF_ID_o(s_id_out_pc_plus1_p) );
  id_top id_top_inst ( .clk(clk), .rst_n(n33), .id_top_i({
        \mini_mips_i[IMEM_DATA][31] , \mini_mips_i[IMEM_DATA][30] , 
        \mini_mips_i[IMEM_DATA][29] , \mini_mips_i[IMEM_DATA][28] , 
        \mini_mips_i[IMEM_DATA][27] , \mini_mips_i[IMEM_DATA][26] , 
        \mini_mips_i[IMEM_DATA][25] , \mini_mips_i[IMEM_DATA][24] , 
        \mini_mips_i[IMEM_DATA][23] , \mini_mips_i[IMEM_DATA][22] , 
        \mini_mips_i[IMEM_DATA][21] , \mini_mips_i[IMEM_DATA][20] , 
        \mini_mips_i[IMEM_DATA][19] , \mini_mips_i[IMEM_DATA][18] , 
        \mini_mips_i[IMEM_DATA][17] , \mini_mips_i[IMEM_DATA][16] , 
        \mini_mips_i[IMEM_DATA][15] , \mini_mips_i[IMEM_DATA][14] , 
        \mini_mips_i[IMEM_DATA][13] , \mini_mips_i[IMEM_DATA][12] , 
        \mini_mips_i[IMEM_DATA][11] , \mini_mips_i[IMEM_DATA][10] , 
        \mini_mips_i[IMEM_DATA][9] , \mini_mips_i[IMEM_DATA][8] , 
        \mini_mips_i[IMEM_DATA][7] , \mini_mips_i[IMEM_DATA][6] , 
        \mini_mips_i[IMEM_DATA][5] , \mini_mips_i[IMEM_DATA][4] , 
        \mini_mips_i[IMEM_DATA][3] , \mini_mips_i[IMEM_DATA][2] , 
        \mini_mips_i[IMEM_DATA][1] , \mini_mips_i[IMEM_DATA][0] , 
        s_writeback_data, s_regfile_forward_A, s_regfile_forward_B, 
        s_wb_in_regWrite_p, s_wb_in_write_reg_p}), .id_top_o({s_id_out_regA_p, 
        s_id_out_regB_p, s_id_ctrl_opcode, s_id_out_RS_p, s_id_out_RT_p, 
        s_id_out_RD_p, s_id_out_shamt_p, s_id_out_funct_p, 
        s_id_out_sign_extend_p}) );
  id_exe id_exe_inst ( .clk(clk), .rst_n(n34), .halt_i(1'b0), .ID_EXE_i({
        s_id_out_regA_p, s_id_out_regB_p, s_id_out_shamt_p, s_id_out_funct_p, 
        s_id_out_sign_extend_p, s_id_out_pc_plus1_p, s_id_out_RS_p, 
        s_id_out_RT_p, s_id_out_RD_p, s_ctrl_out_ALUsrc_B_p, 
        s_ctrl_out_memtoReg_p, s_ctrl_out_regWrite_p, s_ctrl_out_memWen_n_p, 
        1'b0, s_ctrl_out_cALU_OP_p[2:0], s_ctrl_out_RegDst_p}), .ID_EXE_o({
        s_exe_in_regA_p, s_exe_in_regB_p, s_exe_in_shamt_p, s_exe_in_funct_p, 
        s_exe_in_sign_extend_p, s_exe_in_pc_plus1_p, s_exe_in_RS_p, 
        s_exe_in_RT_p, s_exe_in_RD_p, s_exe_in_ALUsrc_B_p, 
        s_exe_out_memtoReg_p, s_exe_out_regWrite_p, s_exe_out_memWen_n_p, 
        s_exe_in_cALU_OP_p, s_exe_in_RegDst_p}) );
  exe_top exe_top_inst ( .clk(clk), .rst_n(n33), .exe_top_i({s_exe_in_shamt_p, 
        s_src_a, s_src_b, s_exe_in_ALUsrc_B_p, s_exe_in_sign_extend_p, 
        s_exe_in_cALU_OP_p, s_exe_in_funct_p, s_exe_in_pc_plus1_p, 
        s_exe_in_RegDst_p, s_exe_in_RT_p, s_exe_in_RD_p}), .exe_top_o({
        s_if_PCSrc, s_exe_if_branch_pc, s_exe_out_alu_res_p, 
        s_exe_out_write_reg_p, s_exe_out_dmem_data_p}) );
  forwarding_unit forwarding_unit_inst ( .forwarding_unit_i({s_exe_in_RS_p, 
        s_exe_in_RT_p, s_id_out_RS_p, s_id_out_RT_p, s_mem_out_write_reg_p, 
        s_wb_in_write_reg_p, s_mem_out_regWrite_p, s_wb_in_regWrite_p}), 
        .forwarding_unit_o({s_forward_A, s_forward_B, s_regfile_forward_A, 
        s_regfile_forward_B}) );
  exe_mem exe_mem_inst ( .clk(clk), .rst_n(n33), .halt_i(1'b0), .EXE_MEM_i({
        s_exe_out_alu_res_p, s_exe_out_dmem_data_p, s_exe_out_write_reg_p, 
        s_exe_out_memtoReg_p, s_exe_out_regWrite_p, s_exe_out_memWen_n_p}), 
        .EXE_MEM_o({s_mem_out_alu_res_p, \mini_mips_o[DMEM_ADDR][11] , 
        \mini_mips_o[DMEM_ADDR][10] , \mini_mips_o[DMEM_ADDR][9] , 
        \mini_mips_o[DMEM_ADDR][8] , \mini_mips_o[DMEM_ADDR][7] , 
        \mini_mips_o[DMEM_ADDR][6] , \mini_mips_o[DMEM_ADDR][5] , 
        \mini_mips_o[DMEM_ADDR][4] , \mini_mips_o[DMEM_ADDR][3] , 
        \mini_mips_o[DMEM_ADDR][2] , \mini_mips_o[DMEM_ADDR][1] , 
        \mini_mips_o[DMEM_ADDR][0] , \mini_mips_o[DMEM_DATA][31] , 
        \mini_mips_o[DMEM_DATA][30] , \mini_mips_o[DMEM_DATA][29] , 
        \mini_mips_o[DMEM_DATA][28] , \mini_mips_o[DMEM_DATA][27] , 
        \mini_mips_o[DMEM_DATA][26] , \mini_mips_o[DMEM_DATA][25] , 
        \mini_mips_o[DMEM_DATA][24] , \mini_mips_o[DMEM_DATA][23] , 
        \mini_mips_o[DMEM_DATA][22] , \mini_mips_o[DMEM_DATA][21] , 
        \mini_mips_o[DMEM_DATA][20] , \mini_mips_o[DMEM_DATA][19] , 
        \mini_mips_o[DMEM_DATA][18] , \mini_mips_o[DMEM_DATA][17] , 
        \mini_mips_o[DMEM_DATA][16] , \mini_mips_o[DMEM_DATA][15] , 
        \mini_mips_o[DMEM_DATA][14] , \mini_mips_o[DMEM_DATA][13] , 
        \mini_mips_o[DMEM_DATA][12] , \mini_mips_o[DMEM_DATA][11] , 
        \mini_mips_o[DMEM_DATA][10] , \mini_mips_o[DMEM_DATA][9] , 
        \mini_mips_o[DMEM_DATA][8] , \mini_mips_o[DMEM_DATA][7] , 
        \mini_mips_o[DMEM_DATA][6] , \mini_mips_o[DMEM_DATA][5] , 
        \mini_mips_o[DMEM_DATA][4] , \mini_mips_o[DMEM_DATA][3] , 
        \mini_mips_o[DMEM_DATA][2] , \mini_mips_o[DMEM_DATA][1] , 
        \mini_mips_o[DMEM_DATA][0] , s_mem_out_write_reg_p, 
        s_mem_out_memtoReg_p, s_mem_out_regWrite_p, \mini_mips_o[DMEM_WEN_N] }) );
  mem_wb mem_wb_inst ( .clk(clk), .rst_n(n34), .halt_i(1'b0), .MEM_WB_i({
        s_mem_out_alu_res_p, \mini_mips_o[DMEM_ADDR][11] , 
        \mini_mips_o[DMEM_ADDR][10] , \mini_mips_o[DMEM_ADDR][9] , 
        \mini_mips_o[DMEM_ADDR][8] , \mini_mips_o[DMEM_ADDR][7] , 
        \mini_mips_o[DMEM_ADDR][6] , \mini_mips_o[DMEM_ADDR][5] , 
        \mini_mips_o[DMEM_ADDR][4] , \mini_mips_o[DMEM_ADDR][3] , 
        \mini_mips_o[DMEM_ADDR][2] , \mini_mips_o[DMEM_ADDR][1] , 
        \mini_mips_o[DMEM_ADDR][0] , s_mem_out_write_reg_p, 
        s_mem_out_memtoReg_p, s_mem_out_regWrite_p}), .MEM_WB_o({
        s_wb_in_alu_res_p, s_wb_in_write_reg_p, s_wb_in_memtoReg_p, 
        s_wb_in_regWrite_p}) );
  HS65_LHS_XNOR2X6 U2 ( .A(s_forward_A[0]), .B(s_forward_A[1]), .Z(n1) );
  HS65_LHS_XNOR2X6 U3 ( .A(s_forward_B[0]), .B(s_forward_B[1]), .Z(n2) );
  HS65_LH_AND2X4 U4 ( .A(s_forward_A[1]), .B(n36), .Z(n9) );
  HS65_LH_AND2X4 U5 ( .A(s_forward_B[1]), .B(n37), .Z(n6) );
  HS65_LH_BFX9 U6 ( .A(n9), .Z(n5) );
  HS65_LH_BFX9 U7 ( .A(n9), .Z(n8) );
  HS65_LH_BFX9 U8 ( .A(n13), .Z(n15) );
  HS65_LH_BFX9 U9 ( .A(n1), .Z(n11) );
  HS65_LH_BFX9 U10 ( .A(n1), .Z(n12) );
  HS65_LH_BFX9 U11 ( .A(n31), .Z(n29) );
  HS65_LH_BFX9 U12 ( .A(n9), .Z(n3) );
  HS65_LH_BFX9 U13 ( .A(n6), .Z(n17) );
  HS65_LH_BFX9 U14 ( .A(n6), .Z(n18) );
  HS65_LH_BFX9 U15 ( .A(n6), .Z(n19) );
  HS65_LH_BFX9 U16 ( .A(n13), .Z(n14) );
  HS65_LH_BFX9 U17 ( .A(n23), .Z(n24) );
  HS65_LH_BFX9 U18 ( .A(n23), .Z(n25) );
  HS65_LH_BFX9 U19 ( .A(n1), .Z(n10) );
  HS65_LH_BFX9 U20 ( .A(n2), .Z(n20) );
  HS65_LH_BFX9 U21 ( .A(n2), .Z(n21) );
  HS65_LH_IVX9 U22 ( .A(n28), .Z(n27) );
  HS65_LH_BFX9 U23 ( .A(n23), .Z(n26) );
  HS65_LH_BFX9 U24 ( .A(n13), .Z(n16) );
  HS65_LH_BFX9 U25 ( .A(n2), .Z(n22) );
  HS65_LH_BFX9 U26 ( .A(n31), .Z(n30) );
  HS65_LH_IVX9 U27 ( .A(s_forward_A[0]), .Z(n36) );
  HS65_LH_BFX9 U28 ( .A(n7), .Z(n13) );
  HS65_LH_NOR2X6 U29 ( .A(n36), .B(s_forward_A[1]), .Z(n7) );
  HS65_LH_IVX9 U30 ( .A(s_forward_B[0]), .Z(n37) );
  HS65_LH_BFX9 U31 ( .A(n31), .Z(n28) );
  HS65_LH_IVX9 U32 ( .A(s_wb_in_memtoReg_p), .Z(n31) );
  HS65_LH_BFX9 U33 ( .A(n4), .Z(n23) );
  HS65_LH_NOR2X6 U34 ( .A(n37), .B(s_forward_B[1]), .Z(n4) );
  HS65_LH_BFX9 U35 ( .A(n32), .Z(n33) );
  HS65_LH_BFX9 U36 ( .A(n32), .Z(n34) );
  HS65_LH_BFX9 U37 ( .A(n32), .Z(n35) );
  HS65_LH_AO222X4 U38 ( .A(n25), .B(s_writeback_data[2]), .C(
        s_exe_in_regB_p[2]), .D(n21), .E(\mini_mips_o[DMEM_ADDR][2] ), .F(n18), 
        .Z(s_src_b[2]) );
  HS65_LH_AO222X4 U39 ( .A(n24), .B(s_writeback_data[0]), .C(
        s_exe_in_regB_p[0]), .D(n20), .E(\mini_mips_o[DMEM_ADDR][0] ), .F(n17), 
        .Z(s_src_b[0]) );
  HS65_LH_AO22X9 U40 ( .A(s_wb_in_alu_res_p[1]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][1] ), .D(n27), .Z(s_writeback_data[1]) );
  HS65_LH_AO22X9 U41 ( .A(s_wb_in_alu_res_p[2]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][2] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[2]) );
  HS65_LH_AO22X9 U42 ( .A(s_wb_in_alu_res_p[4]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][4] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[4]) );
  HS65_LH_AO22X9 U43 ( .A(s_wb_in_alu_res_p[3]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][3] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[3]) );
  HS65_LH_AO22X9 U44 ( .A(s_wb_in_alu_res_p[5]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][5] ), .D(n27), .Z(s_writeback_data[5]) );
  HS65_LH_AO22X9 U45 ( .A(s_wb_in_alu_res_p[8]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][8] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[8]) );
  HS65_LH_AO22X9 U46 ( .A(s_wb_in_alu_res_p[0]), .B(n28), .C(
        \mini_mips_i[DMEM_DATA][0] ), .D(n27), .Z(s_writeback_data[0]) );
  HS65_LH_AO222X4 U47 ( .A(n14), .B(s_writeback_data[1]), .C(
        s_exe_in_regA_p[1]), .D(n10), .E(n3), .F(\mini_mips_o[DMEM_ADDR][1] ), 
        .Z(s_src_a[1]) );
  HS65_LH_AO222X4 U48 ( .A(n15), .B(s_writeback_data[2]), .C(
        s_exe_in_regA_p[2]), .D(n11), .E(n5), .F(\mini_mips_o[DMEM_ADDR][2] ), 
        .Z(s_src_a[2]) );
  HS65_LH_AO222X4 U49 ( .A(n16), .B(s_writeback_data[4]), .C(
        s_exe_in_regA_p[4]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][4] ), 
        .Z(s_src_a[4]) );
  HS65_LH_AO222X4 U50 ( .A(n16), .B(s_writeback_data[3]), .C(
        s_exe_in_regA_p[3]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][3] ), 
        .Z(s_src_a[3]) );
  HS65_LH_AO222X4 U51 ( .A(n16), .B(s_writeback_data[5]), .C(
        s_exe_in_regA_p[5]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][5] ), 
        .Z(s_src_a[5]) );
  HS65_LH_AO222X4 U52 ( .A(n16), .B(s_writeback_data[8]), .C(
        s_exe_in_regA_p[8]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][8] ), 
        .Z(s_src_a[8]) );
  HS65_LH_AO222X4 U53 ( .A(n14), .B(s_writeback_data[0]), .C(
        s_exe_in_regA_p[0]), .D(n10), .E(n3), .F(\mini_mips_o[DMEM_ADDR][0] ), 
        .Z(s_src_a[0]) );
  HS65_LH_AO222X4 U54 ( .A(n14), .B(s_writeback_data[16]), .C(
        s_exe_in_regA_p[16]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[16]), 
        .Z(s_src_a[16]) );
  HS65_LH_AO222X4 U55 ( .A(n14), .B(s_writeback_data[15]), .C(
        s_exe_in_regA_p[15]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[15]), 
        .Z(s_src_a[15]) );
  HS65_LH_AO222X4 U56 ( .A(n14), .B(s_writeback_data[13]), .C(
        s_exe_in_regA_p[13]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[13]), 
        .Z(s_src_a[13]) );
  HS65_LH_AO222X4 U57 ( .A(n14), .B(s_writeback_data[14]), .C(
        s_exe_in_regA_p[14]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[14]), 
        .Z(s_src_a[14]) );
  HS65_LH_AO222X4 U58 ( .A(n14), .B(s_writeback_data[17]), .C(
        s_exe_in_regA_p[17]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[17]), 
        .Z(s_src_a[17]) );
  HS65_LH_AO222X4 U59 ( .A(n15), .B(s_writeback_data[20]), .C(
        s_exe_in_regA_p[20]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[20]), 
        .Z(s_src_a[20]) );
  HS65_LH_AO222X4 U60 ( .A(n26), .B(s_writeback_data[3]), .C(
        s_exe_in_regB_p[3]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][3] ), .F(n19), 
        .Z(s_src_b[3]) );
  HS65_LH_AO222X4 U61 ( .A(n24), .B(s_writeback_data[1]), .C(
        s_exe_in_regB_p[1]), .D(n20), .E(\mini_mips_o[DMEM_ADDR][1] ), .F(n17), 
        .Z(s_src_b[1]) );
  HS65_LH_AO222X4 U62 ( .A(n26), .B(s_writeback_data[4]), .C(
        s_exe_in_regB_p[4]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][4] ), .F(n19), 
        .Z(s_src_b[4]) );
  HS65_LH_AO222X4 U63 ( .A(n26), .B(s_writeback_data[5]), .C(
        s_exe_in_regB_p[5]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][5] ), .F(n19), 
        .Z(s_src_b[5]) );
  HS65_LH_AO222X4 U64 ( .A(n26), .B(s_writeback_data[6]), .C(
        s_exe_in_regB_p[6]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][6] ), .F(n19), 
        .Z(s_src_b[6]) );
  HS65_LH_AO222X4 U65 ( .A(n26), .B(s_writeback_data[7]), .C(
        s_exe_in_regB_p[7]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][7] ), .F(n19), 
        .Z(s_src_b[7]) );
  HS65_LH_AO222X4 U66 ( .A(n26), .B(s_writeback_data[8]), .C(
        s_exe_in_regB_p[8]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][8] ), .F(n19), 
        .Z(s_src_b[8]) );
  HS65_LH_AO22X9 U67 ( .A(s_wb_in_alu_res_p[20]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][20] ), .D(n27), .Z(s_writeback_data[20]) );
  HS65_LH_AO22X9 U68 ( .A(s_wb_in_alu_res_p[14]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][14] ), .D(n27), .Z(s_writeback_data[14]) );
  HS65_LH_AO22X9 U69 ( .A(s_wb_in_alu_res_p[17]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][17] ), .D(n27), .Z(s_writeback_data[17]) );
  HS65_LH_AO22X9 U70 ( .A(s_wb_in_alu_res_p[6]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][6] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[6]) );
  HS65_LH_AO22X9 U71 ( .A(s_wb_in_alu_res_p[7]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][7] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[7]) );
  HS65_LH_AO22X9 U72 ( .A(s_wb_in_alu_res_p[9]), .B(n30), .C(
        s_wb_in_memtoReg_p), .D(\mini_mips_i[DMEM_DATA][9] ), .Z(
        s_writeback_data[9]) );
  HS65_LH_AO22X9 U73 ( .A(s_wb_in_alu_res_p[10]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][10] ), .D(n27), .Z(s_writeback_data[10]) );
  HS65_LH_AO22X9 U74 ( .A(s_wb_in_alu_res_p[11]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][11] ), .D(n27), .Z(s_writeback_data[11]) );
  HS65_LH_AO22X9 U75 ( .A(s_wb_in_alu_res_p[12]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][12] ), .D(n27), .Z(s_writeback_data[12]) );
  HS65_LH_AO22X9 U76 ( .A(s_wb_in_alu_res_p[13]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][13] ), .D(n27), .Z(s_writeback_data[13]) );
  HS65_LH_AO22X9 U77 ( .A(s_wb_in_alu_res_p[15]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][15] ), .D(n27), .Z(s_writeback_data[15]) );
  HS65_LH_AO22X9 U78 ( .A(s_wb_in_alu_res_p[16]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][16] ), .D(n27), .Z(s_writeback_data[16]) );
  HS65_LH_AO22X9 U79 ( .A(s_wb_in_alu_res_p[18]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][18] ), .D(n27), .Z(s_writeback_data[18]) );
  HS65_LH_AO222X4 U80 ( .A(n16), .B(s_writeback_data[6]), .C(
        s_exe_in_regA_p[6]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][6] ), 
        .Z(s_src_a[6]) );
  HS65_LH_AO222X4 U81 ( .A(n16), .B(s_writeback_data[7]), .C(
        s_exe_in_regA_p[7]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][7] ), 
        .Z(s_src_a[7]) );
  HS65_LH_AO222X4 U82 ( .A(n16), .B(s_writeback_data[9]), .C(
        s_exe_in_regA_p[9]), .D(n12), .E(n8), .F(\mini_mips_o[DMEM_ADDR][9] ), 
        .Z(s_src_a[9]) );
  HS65_LH_AO222X4 U83 ( .A(n14), .B(s_writeback_data[10]), .C(
        s_exe_in_regA_p[10]), .D(n10), .E(n3), .F(\mini_mips_o[DMEM_ADDR][10] ), .Z(s_src_a[10]) );
  HS65_LH_AO222X4 U84 ( .A(n14), .B(s_writeback_data[11]), .C(
        s_exe_in_regA_p[11]), .D(n10), .E(n3), .F(\mini_mips_o[DMEM_ADDR][11] ), .Z(s_src_a[11]) );
  HS65_LH_AO222X4 U85 ( .A(n14), .B(s_writeback_data[12]), .C(
        s_exe_in_regA_p[12]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[12]), 
        .Z(s_src_a[12]) );
  HS65_LH_AO222X4 U86 ( .A(n14), .B(s_writeback_data[18]), .C(
        s_exe_in_regA_p[18]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[18]), 
        .Z(s_src_a[18]) );
  HS65_LH_AO222X4 U87 ( .A(n15), .B(s_writeback_data[28]), .C(
        s_exe_in_regA_p[28]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[28]), 
        .Z(s_src_a[28]) );
  HS65_LH_AO222X4 U88 ( .A(n15), .B(s_writeback_data[22]), .C(
        s_exe_in_regA_p[22]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[22]), 
        .Z(s_src_a[22]) );
  HS65_LH_AO222X4 U89 ( .A(n15), .B(s_writeback_data[24]), .C(
        s_exe_in_regA_p[24]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[24]), 
        .Z(s_src_a[24]) );
  HS65_LH_AO222X4 U90 ( .A(n15), .B(s_writeback_data[21]), .C(
        s_exe_in_regA_p[21]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[21]), 
        .Z(s_src_a[21]) );
  HS65_LH_AO222X4 U91 ( .A(n15), .B(s_writeback_data[27]), .C(
        s_exe_in_regA_p[27]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[27]), 
        .Z(s_src_a[27]) );
  HS65_LH_AO222X4 U92 ( .A(n15), .B(s_writeback_data[25]), .C(
        s_exe_in_regA_p[25]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[25]), 
        .Z(s_src_a[25]) );
  HS65_LH_AO222X4 U93 ( .A(n14), .B(s_writeback_data[19]), .C(
        s_exe_in_regA_p[19]), .D(n10), .E(n3), .F(s_mem_out_alu_res_p[19]), 
        .Z(s_src_a[19]) );
  HS65_LH_AO222X4 U94 ( .A(n15), .B(s_writeback_data[23]), .C(
        s_exe_in_regA_p[23]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[23]), 
        .Z(s_src_a[23]) );
  HS65_LH_AO222X4 U95 ( .A(n15), .B(s_writeback_data[26]), .C(
        s_exe_in_regA_p[26]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[26]), 
        .Z(s_src_a[26]) );
  HS65_LH_AO222X4 U96 ( .A(n26), .B(s_writeback_data[9]), .C(
        s_exe_in_regB_p[9]), .D(n22), .E(\mini_mips_o[DMEM_ADDR][9] ), .F(n19), 
        .Z(s_src_b[9]) );
  HS65_LH_AO222X4 U97 ( .A(n24), .B(s_writeback_data[10]), .C(
        s_exe_in_regB_p[10]), .D(n20), .E(\mini_mips_o[DMEM_ADDR][10] ), .F(
        n17), .Z(s_src_b[10]) );
  HS65_LH_AO222X4 U98 ( .A(n24), .B(s_writeback_data[11]), .C(
        s_exe_in_regB_p[11]), .D(n20), .E(\mini_mips_o[DMEM_ADDR][11] ), .F(
        n17), .Z(s_src_b[11]) );
  HS65_LH_AO222X4 U99 ( .A(n24), .B(s_writeback_data[12]), .C(
        s_exe_in_regB_p[12]), .D(n20), .E(s_mem_out_alu_res_p[12]), .F(n17), 
        .Z(s_src_b[12]) );
  HS65_LH_AO222X4 U100 ( .A(n24), .B(s_writeback_data[13]), .C(
        s_exe_in_regB_p[13]), .D(n20), .E(s_mem_out_alu_res_p[13]), .F(n17), 
        .Z(s_src_b[13]) );
  HS65_LH_AO222X4 U101 ( .A(n24), .B(s_writeback_data[14]), .C(
        s_exe_in_regB_p[14]), .D(n20), .E(s_mem_out_alu_res_p[14]), .F(n17), 
        .Z(s_src_b[14]) );
  HS65_LH_AO22X9 U102 ( .A(s_wb_in_alu_res_p[27]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][27] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[27]) );
  HS65_LH_AO22X9 U103 ( .A(s_wb_in_alu_res_p[23]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][23] ), .D(n27), .Z(s_writeback_data[23]) );
  HS65_LH_AO22X9 U104 ( .A(s_wb_in_alu_res_p[26]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][26] ), .D(n27), .Z(s_writeback_data[26]) );
  HS65_LH_AO22X9 U105 ( .A(s_wb_in_alu_res_p[29]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][29] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[29]) );
  HS65_LH_AO22X9 U106 ( .A(s_wb_in_alu_res_p[28]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][28] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[28]) );
  HS65_LH_AO22X9 U107 ( .A(s_wb_in_alu_res_p[19]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][19] ), .D(n27), .Z(s_writeback_data[19]) );
  HS65_LH_AO22X9 U108 ( .A(s_wb_in_alu_res_p[21]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][21] ), .D(n27), .Z(s_writeback_data[21]) );
  HS65_LH_AO22X9 U109 ( .A(s_wb_in_alu_res_p[22]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][22] ), .D(n27), .Z(s_writeback_data[22]) );
  HS65_LH_AO22X9 U110 ( .A(s_wb_in_alu_res_p[24]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][24] ), .D(n27), .Z(s_writeback_data[24]) );
  HS65_LH_AO22X9 U111 ( .A(s_wb_in_alu_res_p[25]), .B(n29), .C(
        \mini_mips_i[DMEM_DATA][25] ), .D(n27), .Z(s_writeback_data[25]) );
  HS65_LH_AO222X4 U112 ( .A(n15), .B(s_writeback_data[29]), .C(
        s_exe_in_regA_p[29]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[29]), 
        .Z(s_src_a[29]) );
  HS65_LH_AO222X4 U113 ( .A(n15), .B(s_writeback_data[30]), .C(
        s_exe_in_regA_p[30]), .D(n11), .E(n5), .F(s_mem_out_alu_res_p[30]), 
        .Z(s_src_a[30]) );
  HS65_LH_AO222X4 U114 ( .A(n24), .B(s_writeback_data[15]), .C(
        s_exe_in_regB_p[15]), .D(n20), .E(s_mem_out_alu_res_p[15]), .F(n17), 
        .Z(s_src_b[15]) );
  HS65_LH_AO222X4 U115 ( .A(n24), .B(s_writeback_data[16]), .C(
        s_exe_in_regB_p[16]), .D(n20), .E(s_mem_out_alu_res_p[16]), .F(n17), 
        .Z(s_src_b[16]) );
  HS65_LH_AO222X4 U116 ( .A(n24), .B(s_writeback_data[17]), .C(
        s_exe_in_regB_p[17]), .D(n20), .E(s_mem_out_alu_res_p[17]), .F(n17), 
        .Z(s_src_b[17]) );
  HS65_LH_AO222X4 U117 ( .A(n24), .B(s_writeback_data[18]), .C(
        s_exe_in_regB_p[18]), .D(n20), .E(s_mem_out_alu_res_p[18]), .F(n17), 
        .Z(s_src_b[18]) );
  HS65_LH_AO222X4 U118 ( .A(n24), .B(s_writeback_data[19]), .C(
        s_exe_in_regB_p[19]), .D(n20), .E(s_mem_out_alu_res_p[19]), .F(n17), 
        .Z(s_src_b[19]) );
  HS65_LH_AO222X4 U119 ( .A(n25), .B(s_writeback_data[20]), .C(
        s_exe_in_regB_p[20]), .D(n21), .E(s_mem_out_alu_res_p[20]), .F(n18), 
        .Z(s_src_b[20]) );
  HS65_LH_AO222X4 U120 ( .A(n25), .B(s_writeback_data[21]), .C(
        s_exe_in_regB_p[21]), .D(n21), .E(s_mem_out_alu_res_p[21]), .F(n18), 
        .Z(s_src_b[21]) );
  HS65_LH_AO22X9 U121 ( .A(s_wb_in_alu_res_p[30]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][30] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[30]) );
  HS65_LH_AO22X9 U122 ( .A(s_wb_in_alu_res_p[31]), .B(n30), .C(
        \mini_mips_i[DMEM_DATA][31] ), .D(s_wb_in_memtoReg_p), .Z(
        s_writeback_data[31]) );
  HS65_LH_AO222X4 U123 ( .A(n16), .B(s_writeback_data[31]), .C(
        s_exe_in_regA_p[31]), .D(n12), .E(n8), .F(s_mem_out_alu_res_p[31]), 
        .Z(s_src_a[31]) );
  HS65_LH_AO222X4 U124 ( .A(n25), .B(s_writeback_data[28]), .C(
        s_exe_in_regB_p[28]), .D(n21), .E(s_mem_out_alu_res_p[28]), .F(n18), 
        .Z(s_src_b[28]) );
  HS65_LH_AO222X4 U125 ( .A(n25), .B(s_writeback_data[22]), .C(
        s_exe_in_regB_p[22]), .D(n21), .E(s_mem_out_alu_res_p[22]), .F(n18), 
        .Z(s_src_b[22]) );
  HS65_LH_AO222X4 U126 ( .A(n25), .B(s_writeback_data[23]), .C(
        s_exe_in_regB_p[23]), .D(n21), .E(s_mem_out_alu_res_p[23]), .F(n18), 
        .Z(s_src_b[23]) );
  HS65_LH_AO222X4 U127 ( .A(n25), .B(s_writeback_data[24]), .C(
        s_exe_in_regB_p[24]), .D(n21), .E(s_mem_out_alu_res_p[24]), .F(n18), 
        .Z(s_src_b[24]) );
  HS65_LH_AO222X4 U128 ( .A(n25), .B(s_writeback_data[25]), .C(
        s_exe_in_regB_p[25]), .D(n21), .E(s_mem_out_alu_res_p[25]), .F(n18), 
        .Z(s_src_b[25]) );
  HS65_LH_AO222X4 U129 ( .A(n25), .B(s_writeback_data[26]), .C(
        s_exe_in_regB_p[26]), .D(n21), .E(s_mem_out_alu_res_p[26]), .F(n18), 
        .Z(s_src_b[26]) );
  HS65_LH_AO222X4 U130 ( .A(n25), .B(s_writeback_data[27]), .C(
        s_exe_in_regB_p[27]), .D(n21), .E(s_mem_out_alu_res_p[27]), .F(n18), 
        .Z(s_src_b[27]) );
  HS65_LH_AO222X4 U131 ( .A(n26), .B(s_writeback_data[31]), .C(
        s_exe_in_regB_p[31]), .D(n22), .E(s_mem_out_alu_res_p[31]), .F(n19), 
        .Z(s_src_b[31]) );
  HS65_LH_AO222X4 U132 ( .A(n25), .B(s_writeback_data[29]), .C(
        s_exe_in_regB_p[29]), .D(n21), .E(s_mem_out_alu_res_p[29]), .F(n18), 
        .Z(s_src_b[29]) );
  HS65_LH_AO222X4 U133 ( .A(n25), .B(s_writeback_data[30]), .C(
        s_exe_in_regB_p[30]), .D(n21), .E(s_mem_out_alu_res_p[30]), .F(n18), 
        .Z(s_src_b[30]) );
  HS65_LH_BFX9 U134 ( .A(rst_n), .Z(n32) );
endmodule


module mini_mips_p ( clk, rst_n );
  inout clk,  rst_n;
  wire   clk_i, rst_n_i, \s_mini_mips_i[DMEM_DATA][31] ,
         \s_mini_mips_i[DMEM_DATA][30] , \s_mini_mips_i[DMEM_DATA][29] ,
         \s_mini_mips_i[DMEM_DATA][28] , \s_mini_mips_i[DMEM_DATA][27] ,
         \s_mini_mips_i[DMEM_DATA][26] , \s_mini_mips_i[DMEM_DATA][25] ,
         \s_mini_mips_i[DMEM_DATA][24] , \s_mini_mips_i[DMEM_DATA][23] ,
         \s_mini_mips_i[DMEM_DATA][22] , \s_mini_mips_i[DMEM_DATA][21] ,
         \s_mini_mips_i[DMEM_DATA][20] , \s_mini_mips_i[DMEM_DATA][19] ,
         \s_mini_mips_i[DMEM_DATA][18] , \s_mini_mips_i[DMEM_DATA][17] ,
         \s_mini_mips_i[DMEM_DATA][16] , \s_mini_mips_i[DMEM_DATA][15] ,
         \s_mini_mips_i[DMEM_DATA][14] , \s_mini_mips_i[DMEM_DATA][13] ,
         \s_mini_mips_i[DMEM_DATA][12] , \s_mini_mips_i[DMEM_DATA][11] ,
         \s_mini_mips_i[DMEM_DATA][10] , \s_mini_mips_i[DMEM_DATA][9] ,
         \s_mini_mips_i[DMEM_DATA][8] , \s_mini_mips_i[DMEM_DATA][7] ,
         \s_mini_mips_i[DMEM_DATA][6] , \s_mini_mips_i[DMEM_DATA][5] ,
         \s_mini_mips_i[DMEM_DATA][4] , \s_mini_mips_i[DMEM_DATA][3] ,
         \s_mini_mips_i[DMEM_DATA][2] , \s_mini_mips_i[DMEM_DATA][1] ,
         \s_mini_mips_i[DMEM_DATA][0] , \s_mini_mips_i[IMEM_DATA][31] ,
         \s_mini_mips_i[IMEM_DATA][30] , \s_mini_mips_i[IMEM_DATA][29] ,
         \s_mini_mips_i[IMEM_DATA][28] , \s_mini_mips_i[IMEM_DATA][27] ,
         \s_mini_mips_i[IMEM_DATA][26] , \s_mini_mips_i[IMEM_DATA][25] ,
         \s_mini_mips_i[IMEM_DATA][24] , \s_mini_mips_i[IMEM_DATA][23] ,
         \s_mini_mips_i[IMEM_DATA][22] , \s_mini_mips_i[IMEM_DATA][21] ,
         \s_mini_mips_i[IMEM_DATA][20] , \s_mini_mips_i[IMEM_DATA][19] ,
         \s_mini_mips_i[IMEM_DATA][18] , \s_mini_mips_i[IMEM_DATA][17] ,
         \s_mini_mips_i[IMEM_DATA][16] , \s_mini_mips_i[IMEM_DATA][15] ,
         \s_mini_mips_i[IMEM_DATA][14] , \s_mini_mips_i[IMEM_DATA][13] ,
         \s_mini_mips_i[IMEM_DATA][12] , \s_mini_mips_i[IMEM_DATA][11] ,
         \s_mini_mips_i[IMEM_DATA][10] , \s_mini_mips_i[IMEM_DATA][9] ,
         \s_mini_mips_i[IMEM_DATA][8] , \s_mini_mips_i[IMEM_DATA][7] ,
         \s_mini_mips_i[IMEM_DATA][6] , \s_mini_mips_i[IMEM_DATA][5] ,
         \s_mini_mips_i[IMEM_DATA][4] , \s_mini_mips_i[IMEM_DATA][3] ,
         \s_mini_mips_i[IMEM_DATA][2] , \s_mini_mips_i[IMEM_DATA][1] ,
         \s_mini_mips_i[IMEM_DATA][0] , \s_mini_mips_o[DMEM_ADDR][11] ,
         \s_mini_mips_o[DMEM_ADDR][10] , \s_mini_mips_o[DMEM_ADDR][9] ,
         \s_mini_mips_o[DMEM_ADDR][8] , \s_mini_mips_o[DMEM_ADDR][7] ,
         \s_mini_mips_o[DMEM_ADDR][6] , \s_mini_mips_o[DMEM_ADDR][5] ,
         \s_mini_mips_o[DMEM_ADDR][4] , \s_mini_mips_o[DMEM_ADDR][3] ,
         \s_mini_mips_o[DMEM_ADDR][2] , \s_mini_mips_o[DMEM_ADDR][1] ,
         \s_mini_mips_o[DMEM_ADDR][0] , \s_mini_mips_o[IMEM_ADDR][11] ,
         \s_mini_mips_o[IMEM_ADDR][10] , \s_mini_mips_o[IMEM_ADDR][9] ,
         \s_mini_mips_o[IMEM_ADDR][8] , \s_mini_mips_o[IMEM_ADDR][7] ,
         \s_mini_mips_o[IMEM_ADDR][6] , \s_mini_mips_o[IMEM_ADDR][5] ,
         \s_mini_mips_o[IMEM_ADDR][4] , \s_mini_mips_o[IMEM_ADDR][3] ,
         \s_mini_mips_o[IMEM_ADDR][2] , \s_mini_mips_o[IMEM_ADDR][1] ,
         \s_mini_mips_o[IMEM_ADDR][0] , \s_mini_mips_o[DMEM_WEN_N] ;
  tri   clk;
  tri   rst_n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;

  ST_SPHDL_4096x32m8_L imem_inst ( .A({\s_mini_mips_o[IMEM_ADDR][11] , 
        \s_mini_mips_o[IMEM_ADDR][10] , \s_mini_mips_o[IMEM_ADDR][9] , 
        \s_mini_mips_o[IMEM_ADDR][8] , \s_mini_mips_o[IMEM_ADDR][7] , 
        \s_mini_mips_o[IMEM_ADDR][6] , \s_mini_mips_o[IMEM_ADDR][5] , 
        \s_mini_mips_o[IMEM_ADDR][4] , \s_mini_mips_o[IMEM_ADDR][3] , 
        \s_mini_mips_o[IMEM_ADDR][2] , \s_mini_mips_o[IMEM_ADDR][1] , 
        \s_mini_mips_o[IMEM_ADDR][0] }), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .Q({\s_mini_mips_i[IMEM_DATA][31] , 
        \s_mini_mips_i[IMEM_DATA][30] , \s_mini_mips_i[IMEM_DATA][29] , 
        \s_mini_mips_i[IMEM_DATA][28] , \s_mini_mips_i[IMEM_DATA][27] , 
        \s_mini_mips_i[IMEM_DATA][26] , \s_mini_mips_i[IMEM_DATA][25] , 
        \s_mini_mips_i[IMEM_DATA][24] , \s_mini_mips_i[IMEM_DATA][23] , 
        \s_mini_mips_i[IMEM_DATA][22] , \s_mini_mips_i[IMEM_DATA][21] , 
        \s_mini_mips_i[IMEM_DATA][20] , \s_mini_mips_i[IMEM_DATA][19] , 
        \s_mini_mips_i[IMEM_DATA][18] , \s_mini_mips_i[IMEM_DATA][17] , 
        \s_mini_mips_i[IMEM_DATA][16] , \s_mini_mips_i[IMEM_DATA][15] , 
        \s_mini_mips_i[IMEM_DATA][14] , \s_mini_mips_i[IMEM_DATA][13] , 
        \s_mini_mips_i[IMEM_DATA][12] , \s_mini_mips_i[IMEM_DATA][11] , 
        \s_mini_mips_i[IMEM_DATA][10] , \s_mini_mips_i[IMEM_DATA][9] , 
        \s_mini_mips_i[IMEM_DATA][8] , \s_mini_mips_i[IMEM_DATA][7] , 
        \s_mini_mips_i[IMEM_DATA][6] , \s_mini_mips_i[IMEM_DATA][5] , 
        \s_mini_mips_i[IMEM_DATA][4] , \s_mini_mips_i[IMEM_DATA][3] , 
        \s_mini_mips_i[IMEM_DATA][2] , \s_mini_mips_i[IMEM_DATA][1] , 
        \s_mini_mips_i[IMEM_DATA][0] }), .CK(clk_i), .CSN(1'b0), .TBYPASS(1'b0), .WEN(1'b1) );
  ST_SPHDL_4096x32m8_L dmem_inst ( .A({\s_mini_mips_o[DMEM_ADDR][11] , 
        \s_mini_mips_o[DMEM_ADDR][10] , \s_mini_mips_o[DMEM_ADDR][9] , 
        \s_mini_mips_o[DMEM_ADDR][8] , \s_mini_mips_o[DMEM_ADDR][7] , 
        \s_mini_mips_o[DMEM_ADDR][6] , \s_mini_mips_o[DMEM_ADDR][5] , 
        \s_mini_mips_o[DMEM_ADDR][4] , \s_mini_mips_o[DMEM_ADDR][3] , 
        \s_mini_mips_o[DMEM_ADDR][2] , \s_mini_mips_o[DMEM_ADDR][1] , 
        \s_mini_mips_o[DMEM_ADDR][0] }), .D({\s_mini_mips_i[DMEM_DATA][31] , 
        \s_mini_mips_i[DMEM_DATA][30] , \s_mini_mips_i[DMEM_DATA][29] , 
        \s_mini_mips_i[DMEM_DATA][28] , \s_mini_mips_i[DMEM_DATA][27] , 
        \s_mini_mips_i[DMEM_DATA][26] , \s_mini_mips_i[DMEM_DATA][25] , 
        \s_mini_mips_i[DMEM_DATA][24] , \s_mini_mips_i[DMEM_DATA][23] , 
        \s_mini_mips_i[DMEM_DATA][22] , \s_mini_mips_i[DMEM_DATA][21] , 
        \s_mini_mips_i[DMEM_DATA][20] , \s_mini_mips_i[DMEM_DATA][19] , 
        \s_mini_mips_i[DMEM_DATA][18] , \s_mini_mips_i[DMEM_DATA][17] , 
        \s_mini_mips_i[DMEM_DATA][16] , \s_mini_mips_i[DMEM_DATA][15] , 
        \s_mini_mips_i[DMEM_DATA][14] , \s_mini_mips_i[DMEM_DATA][13] , 
        \s_mini_mips_i[DMEM_DATA][12] , \s_mini_mips_i[DMEM_DATA][11] , 
        \s_mini_mips_i[DMEM_DATA][10] , \s_mini_mips_i[DMEM_DATA][9] , 
        \s_mini_mips_i[DMEM_DATA][8] , \s_mini_mips_i[DMEM_DATA][7] , 
        \s_mini_mips_i[DMEM_DATA][6] , \s_mini_mips_i[DMEM_DATA][5] , 
        \s_mini_mips_i[DMEM_DATA][4] , \s_mini_mips_i[DMEM_DATA][3] , 
        \s_mini_mips_i[DMEM_DATA][2] , \s_mini_mips_i[DMEM_DATA][1] , 
        \s_mini_mips_i[DMEM_DATA][0] }), .Q({\s_mini_mips_i[DMEM_DATA][31] , 
        \s_mini_mips_i[DMEM_DATA][30] , \s_mini_mips_i[DMEM_DATA][29] , 
        \s_mini_mips_i[DMEM_DATA][28] , \s_mini_mips_i[DMEM_DATA][27] , 
        \s_mini_mips_i[DMEM_DATA][26] , \s_mini_mips_i[DMEM_DATA][25] , 
        \s_mini_mips_i[DMEM_DATA][24] , \s_mini_mips_i[DMEM_DATA][23] , 
        \s_mini_mips_i[DMEM_DATA][22] , \s_mini_mips_i[DMEM_DATA][21] , 
        \s_mini_mips_i[DMEM_DATA][20] , \s_mini_mips_i[DMEM_DATA][19] , 
        \s_mini_mips_i[DMEM_DATA][18] , \s_mini_mips_i[DMEM_DATA][17] , 
        \s_mini_mips_i[DMEM_DATA][16] , \s_mini_mips_i[DMEM_DATA][15] , 
        \s_mini_mips_i[DMEM_DATA][14] , \s_mini_mips_i[DMEM_DATA][13] , 
        \s_mini_mips_i[DMEM_DATA][12] , \s_mini_mips_i[DMEM_DATA][11] , 
        \s_mini_mips_i[DMEM_DATA][10] , \s_mini_mips_i[DMEM_DATA][9] , 
        \s_mini_mips_i[DMEM_DATA][8] , \s_mini_mips_i[DMEM_DATA][7] , 
        \s_mini_mips_i[DMEM_DATA][6] , \s_mini_mips_i[DMEM_DATA][5] , 
        \s_mini_mips_i[DMEM_DATA][4] , \s_mini_mips_i[DMEM_DATA][3] , 
        \s_mini_mips_i[DMEM_DATA][2] , \s_mini_mips_i[DMEM_DATA][1] , 
        \s_mini_mips_i[DMEM_DATA][0] }), .CK(clk_i), .CSN(1'b0), .TBYPASS(1'b0), .WEN(\s_mini_mips_o[DMEM_WEN_N] ) );
  BD2SCARUDQP_1V8_SF_LIN clk_pad_in ( .A(1'b0), .TA(1'b0), .TM(1'b0), .EN(1'b1), .TEN(1'b1), .IO(clk), .HYST(1'b0), .PDN(1'b0), .PUN(1'b0), .ZI(clk_i) );
  BD2SCARUDQP_1V8_SF_LIN rst_n_pad_in ( .A(1'b0), .TA(1'b0), .TM(1'b0), .EN(
        1'b1), .TEN(1'b1), .IO(rst_n), .HYST(1'b0), .PDN(1'b0), .PUN(1'b0), 
        .ZI(rst_n_i) );
  mini_mips_pipeline mini_mips_inst ( .clk(clk_i), .rst_n(rst_n_i), 
        .mini_mips_i({\s_mini_mips_i[DMEM_DATA][31] , 
        \s_mini_mips_i[DMEM_DATA][30] , \s_mini_mips_i[DMEM_DATA][29] , 
        \s_mini_mips_i[DMEM_DATA][28] , \s_mini_mips_i[DMEM_DATA][27] , 
        \s_mini_mips_i[DMEM_DATA][26] , \s_mini_mips_i[DMEM_DATA][25] , 
        \s_mini_mips_i[DMEM_DATA][24] , \s_mini_mips_i[DMEM_DATA][23] , 
        \s_mini_mips_i[DMEM_DATA][22] , \s_mini_mips_i[DMEM_DATA][21] , 
        \s_mini_mips_i[DMEM_DATA][20] , \s_mini_mips_i[DMEM_DATA][19] , 
        \s_mini_mips_i[DMEM_DATA][18] , \s_mini_mips_i[DMEM_DATA][17] , 
        \s_mini_mips_i[DMEM_DATA][16] , \s_mini_mips_i[DMEM_DATA][15] , 
        \s_mini_mips_i[DMEM_DATA][14] , \s_mini_mips_i[DMEM_DATA][13] , 
        \s_mini_mips_i[DMEM_DATA][12] , \s_mini_mips_i[DMEM_DATA][11] , 
        \s_mini_mips_i[DMEM_DATA][10] , \s_mini_mips_i[DMEM_DATA][9] , 
        \s_mini_mips_i[DMEM_DATA][8] , \s_mini_mips_i[DMEM_DATA][7] , 
        \s_mini_mips_i[DMEM_DATA][6] , \s_mini_mips_i[DMEM_DATA][5] , 
        \s_mini_mips_i[DMEM_DATA][4] , \s_mini_mips_i[DMEM_DATA][3] , 
        \s_mini_mips_i[DMEM_DATA][2] , \s_mini_mips_i[DMEM_DATA][1] , 
        \s_mini_mips_i[DMEM_DATA][0] , \s_mini_mips_i[IMEM_DATA][31] , 
        \s_mini_mips_i[IMEM_DATA][30] , \s_mini_mips_i[IMEM_DATA][29] , 
        \s_mini_mips_i[IMEM_DATA][28] , \s_mini_mips_i[IMEM_DATA][27] , 
        \s_mini_mips_i[IMEM_DATA][26] , \s_mini_mips_i[IMEM_DATA][25] , 
        \s_mini_mips_i[IMEM_DATA][24] , \s_mini_mips_i[IMEM_DATA][23] , 
        \s_mini_mips_i[IMEM_DATA][22] , \s_mini_mips_i[IMEM_DATA][21] , 
        \s_mini_mips_i[IMEM_DATA][20] , \s_mini_mips_i[IMEM_DATA][19] , 
        \s_mini_mips_i[IMEM_DATA][18] , \s_mini_mips_i[IMEM_DATA][17] , 
        \s_mini_mips_i[IMEM_DATA][16] , \s_mini_mips_i[IMEM_DATA][15] , 
        \s_mini_mips_i[IMEM_DATA][14] , \s_mini_mips_i[IMEM_DATA][13] , 
        \s_mini_mips_i[IMEM_DATA][12] , \s_mini_mips_i[IMEM_DATA][11] , 
        \s_mini_mips_i[IMEM_DATA][10] , \s_mini_mips_i[IMEM_DATA][9] , 
        \s_mini_mips_i[IMEM_DATA][8] , \s_mini_mips_i[IMEM_DATA][7] , 
        \s_mini_mips_i[IMEM_DATA][6] , \s_mini_mips_i[IMEM_DATA][5] , 
        \s_mini_mips_i[IMEM_DATA][4] , \s_mini_mips_i[IMEM_DATA][3] , 
        \s_mini_mips_i[IMEM_DATA][2] , \s_mini_mips_i[IMEM_DATA][1] , 
        \s_mini_mips_i[IMEM_DATA][0] }), .mini_mips_o({
        \s_mini_mips_o[DMEM_ADDR][11] , \s_mini_mips_o[DMEM_ADDR][10] , 
        \s_mini_mips_o[DMEM_ADDR][9] , \s_mini_mips_o[DMEM_ADDR][8] , 
        \s_mini_mips_o[DMEM_ADDR][7] , \s_mini_mips_o[DMEM_ADDR][6] , 
        \s_mini_mips_o[DMEM_ADDR][5] , \s_mini_mips_o[DMEM_ADDR][4] , 
        \s_mini_mips_o[DMEM_ADDR][3] , \s_mini_mips_o[DMEM_ADDR][2] , 
        \s_mini_mips_o[DMEM_ADDR][1] , \s_mini_mips_o[DMEM_ADDR][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        \s_mini_mips_o[IMEM_ADDR][11] , \s_mini_mips_o[IMEM_ADDR][10] , 
        \s_mini_mips_o[IMEM_ADDR][9] , \s_mini_mips_o[IMEM_ADDR][8] , 
        \s_mini_mips_o[IMEM_ADDR][7] , \s_mini_mips_o[IMEM_ADDR][6] , 
        \s_mini_mips_o[IMEM_ADDR][5] , \s_mini_mips_o[IMEM_ADDR][4] , 
        \s_mini_mips_o[IMEM_ADDR][3] , \s_mini_mips_o[IMEM_ADDR][2] , 
        \s_mini_mips_o[IMEM_ADDR][1] , \s_mini_mips_o[IMEM_ADDR][0] , 
        \s_mini_mips_o[DMEM_WEN_N] }) );
endmodule

