
library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_mult_uns_0 is

   port( a, b : in std_logic_vector (31 downto 0);  product : out 
         std_logic_vector (63 downto 0));

end alu_DW_mult_uns_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_mult_uns_0 is

   component HS65_LHS_XOR2X3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X4
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_HA1X4
      port( A0, B0 : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   signal n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n292, n293, n294, n295, n296, n297, n299, n300, 
      n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n330, n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n354, 
      n355, n356, n357, n358, n359, n360, n361, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094 : std_logic;

begin
   
   U228 : HS65_LH_FA1X4 port map( A0 => n293, B0 => n292, CI => n228, CO => 
                           n227, S0 => product(62));
   U229 : HS65_LH_FA1X4 port map( A0 => n295, B0 => n294, CI => n229, CO => 
                           n228, S0 => product(61));
   U230 : HS65_LH_FA1X4 port map( A0 => n296, B0 => n299, CI => n230, CO => 
                           n229, S0 => product(60));
   U231 : HS65_LH_FA1X4 port map( A0 => n300, B0 => n302, CI => n231, CO => 
                           n230, S0 => product(59));
   U232 : HS65_LH_FA1X4 port map( A0 => n303, B0 => n305, CI => n232, CO => 
                           n231, S0 => product(58));
   U233 : HS65_LH_FA1X4 port map( A0 => n306, B0 => n311, CI => n233, CO => 
                           n232, S0 => product(57));
   U234 : HS65_LH_FA1X4 port map( A0 => n312, B0 => n316, CI => n234, CO => 
                           n233, S0 => product(56));
   U235 : HS65_LH_FA1X4 port map( A0 => n317, B0 => n322, CI => n235, CO => 
                           n234, S0 => product(55));
   U236 : HS65_LH_FA1X4 port map( A0 => n323, B0 => n330, CI => n236, CO => 
                           n235, S0 => product(54));
   U237 : HS65_LH_FA1X4 port map( A0 => n331, B0 => n337, CI => n237, CO => 
                           n236, S0 => product(53));
   U238 : HS65_LH_FA1X4 port map( A0 => n338, B0 => n344, CI => n238, CO => 
                           n237, S0 => product(52));
   U239 : HS65_LH_FA1X4 port map( A0 => n345, B0 => n354, CI => n239, CO => 
                           n238, S0 => product(51));
   U240 : HS65_LH_FA1X4 port map( A0 => n355, B0 => n363, CI => n240, CO => 
                           n239, S0 => product(50));
   U241 : HS65_LH_FA1X4 port map( A0 => n364, B0 => n373, CI => n241, CO => 
                           n240, S0 => product(49));
   U242 : HS65_LH_FA1X4 port map( A0 => n374, B0 => n385, CI => n242, CO => 
                           n241, S0 => product(48));
   U243 : HS65_LH_FA1X4 port map( A0 => n386, B0 => n396, CI => n243, CO => 
                           n242, S0 => product(47));
   U244 : HS65_LH_FA1X4 port map( A0 => n397, B0 => n407, CI => n244, CO => 
                           n243, S0 => product(46));
   U245 : HS65_LH_FA1X4 port map( A0 => n408, B0 => n421, CI => n245, CO => 
                           n244, S0 => product(45));
   U246 : HS65_LH_FA1X4 port map( A0 => n422, B0 => n434, CI => n246, CO => 
                           n245, S0 => product(44));
   U247 : HS65_LH_FA1X4 port map( A0 => n435, B0 => n448, CI => n247, CO => 
                           n246, S0 => product(43));
   U248 : HS65_LH_FA1X4 port map( A0 => n449, B0 => n464, CI => n248, CO => 
                           n247, S0 => product(42));
   U249 : HS65_LH_FA1X4 port map( A0 => n465, B0 => n479, CI => n249, CO => 
                           n248, S0 => product(41));
   U250 : HS65_LH_FA1X4 port map( A0 => n480, B0 => n494, CI => n250, CO => 
                           n249, S0 => product(40));
   U251 : HS65_LH_FA1X4 port map( A0 => n495, B0 => n512, CI => n251, CO => 
                           n250, S0 => product(39));
   U252 : HS65_LH_FA1X4 port map( A0 => n513, B0 => n529, CI => n252, CO => 
                           n251, S0 => product(38));
   U253 : HS65_LH_FA1X4 port map( A0 => n530, B0 => n546, CI => n253, CO => 
                           n252, S0 => product(37));
   U254 : HS65_LH_FA1X4 port map( A0 => n547, B0 => n564, CI => n254, CO => 
                           n253, S0 => product(36));
   U255 : HS65_LH_FA1X4 port map( A0 => n565, B0 => n582, CI => n255, CO => 
                           n254, S0 => product(35));
   U256 : HS65_LH_FA1X4 port map( A0 => n583, B0 => n600, CI => n256, CO => 
                           n255, S0 => product(34));
   U257 : HS65_LH_FA1X4 port map( A0 => n601, B0 => n1386, CI => n257, CO => 
                           n256, S0 => product(33));
   U258 : HS65_LH_FA1X4 port map( A0 => n1387, B0 => n619, CI => n258, CO => 
                           n257, S0 => product(32));
   U259 : HS65_LH_FA1X4 port map( A0 => n1388, B0 => n637, CI => n259, CO => 
                           n258, S0 => product(31));
   U260 : HS65_LH_FA1X4 port map( A0 => n1389, B0 => n655, CI => n260, CO => 
                           n259, S0 => product(30));
   U261 : HS65_LH_FA1X4 port map( A0 => n1390, B0 => n673, CI => n261, CO => 
                           n260, S0 => product(29));
   U262 : HS65_LH_FA1X4 port map( A0 => n1391, B0 => n691, CI => n262, CO => 
                           n261, S0 => product(28));
   U263 : HS65_LH_FA1X4 port map( A0 => n1392, B0 => n709, CI => n263, CO => 
                           n262, S0 => product(27));
   U264 : HS65_LH_FA1X4 port map( A0 => n1393, B0 => n727, CI => n264, CO => 
                           n263, S0 => product(26));
   U265 : HS65_LH_FA1X4 port map( A0 => n1394, B0 => n743, CI => n265, CO => 
                           n264, S0 => product(25));
   U266 : HS65_LH_FA1X4 port map( A0 => n1395, B0 => n759, CI => n266, CO => 
                           n265, S0 => product(24));
   U267 : HS65_LH_FA1X4 port map( A0 => n1396, B0 => n775, CI => n267, CO => 
                           n266, S0 => product(23));
   U268 : HS65_LH_FA1X4 port map( A0 => n1397, B0 => n789, CI => n268, CO => 
                           n267, S0 => product(22));
   U269 : HS65_LH_FA1X4 port map( A0 => n1398, B0 => n803, CI => n269, CO => 
                           n268, S0 => product(21));
   U270 : HS65_LH_FA1X4 port map( A0 => n1399, B0 => n817, CI => n270, CO => 
                           n269, S0 => product(20));
   U271 : HS65_LH_FA1X4 port map( A0 => n1400, B0 => n829, CI => n271, CO => 
                           n270, S0 => product(19));
   U272 : HS65_LH_FA1X4 port map( A0 => n1401, B0 => n841, CI => n272, CO => 
                           n271, S0 => product(18));
   U273 : HS65_LH_FA1X4 port map( A0 => n1402, B0 => n853, CI => n273, CO => 
                           n272, S0 => product(17));
   U274 : HS65_LH_FA1X4 port map( A0 => n1403, B0 => n863, CI => n274, CO => 
                           n273, S0 => product(16));
   U275 : HS65_LH_FA1X4 port map( A0 => n1404, B0 => n873, CI => n275, CO => 
                           n274, S0 => product(15));
   U276 : HS65_LH_FA1X4 port map( A0 => n1405, B0 => n883, CI => n276, CO => 
                           n275, S0 => product(14));
   U277 : HS65_LH_FA1X4 port map( A0 => n1406, B0 => n891, CI => n277, CO => 
                           n276, S0 => product(13));
   U278 : HS65_LH_FA1X4 port map( A0 => n1407, B0 => n899, CI => n278, CO => 
                           n277, S0 => product(12));
   U279 : HS65_LH_FA1X4 port map( A0 => n1408, B0 => n907, CI => n279, CO => 
                           n278, S0 => product(11));
   U280 : HS65_LH_FA1X4 port map( A0 => n1409, B0 => n913, CI => n280, CO => 
                           n279, S0 => product(10));
   U281 : HS65_LH_FA1X4 port map( A0 => n1410, B0 => n919, CI => n281, CO => 
                           n280, S0 => product(9));
   U282 : HS65_LH_FA1X4 port map( A0 => n1411, B0 => n925, CI => n282, CO => 
                           n281, S0 => product(8));
   U283 : HS65_LH_FA1X4 port map( A0 => n1412, B0 => n929, CI => n283, CO => 
                           n282, S0 => product(7));
   U284 : HS65_LH_FA1X4 port map( A0 => n1413, B0 => n933, CI => n284, CO => 
                           n283, S0 => product(6));
   U285 : HS65_LH_FA1X4 port map( A0 => n1414, B0 => n937, CI => n285, CO => 
                           n284, S0 => product(5));
   U286 : HS65_LH_FA1X4 port map( A0 => n1415, B0 => n939, CI => n286, CO => 
                           n285, S0 => product(4));
   U287 : HS65_LH_FA1X4 port map( A0 => n1416, B0 => n941, CI => n287, CO => 
                           n286, S0 => product(3));
   U288 : HS65_LH_HA1X4 port map( A0 => n1417, B0 => n288, CO => n287, S0 => 
                           product(2));
   U289 : HS65_LH_HA1X4 port map( A0 => n1418, B0 => n289, CO => n288, S0 => 
                           product(1));
   U290 : HS65_LH_HA1X4 port map( A0 => a(2), B0 => n1419, CO => n289, S0 => 
                           product(0));
   U293 : HS65_LH_FA1X4 port map( A0 => n297, B0 => n2646, CI => n1041, CO => 
                           n293, S0 => n294);
   U294 : HS65_LH_FA1X4 port map( A0 => n1042, B0 => n2647, CI => n1071, CO => 
                           n295, S0 => n296);
   U296 : HS65_LH_FA1X4 port map( A0 => n2647, B0 => n1043, CI => n1072, CO => 
                           n299, S0 => n300);
   U298 : HS65_LH_FA1X4 port map( A0 => n1073, B0 => n304, CI => n307, CO => 
                           n302, S0 => n303);
   U299 : HS65_LH_FA1X4 port map( A0 => n309, B0 => n2644, CI => n1044, CO => 
                           n297, S0 => n304);
   U300 : HS65_LH_FA1X4 port map( A0 => n1106, B0 => n1074, CI => n308, CO => 
                           n305, S0 => n306);
   U301 : HS65_LH_FA1X4 port map( A0 => n1045, B0 => n2652, CI => n313, CO => 
                           n307, S0 => n308);
   U303 : HS65_LH_FA1X4 port map( A0 => n314, B0 => n318, CI => n1107, CO => 
                           n311, S0 => n312);
   U304 : HS65_LH_FA1X4 port map( A0 => n2652, B0 => n320, CI => n1075, CO => 
                           n313, S0 => n314);
   U306 : HS65_LH_FA1X4 port map( A0 => n1108, B0 => n319, CI => n324, CO => 
                           n316, S0 => n317);
   U307 : HS65_LH_FA1X4 port map( A0 => n326, B0 => n321, CI => n1076, CO => 
                           n318, S0 => n319);
   U308 : HS65_LH_FA1X4 port map( A0 => n328, B0 => n2642, CI => n1046, CO => 
                           n320, S0 => n321);
   U309 : HS65_LH_FA1X4 port map( A0 => n1141, B0 => n1109, CI => n325, CO => 
                           n322, S0 => n323);
   U310 : HS65_LH_FA1X4 port map( A0 => n327, B0 => n334, CI => n332, CO => 
                           n324, S0 => n325);
   U311 : HS65_LH_FA1X4 port map( A0 => n1047, B0 => n2648, CI => n1077, CO => 
                           n326, S0 => n327);
   U313 : HS65_LH_FA1X4 port map( A0 => n333, B0 => n339, CI => n1142, CO => 
                           n330, S0 => n331);
   U314 : HS65_LH_FA1X4 port map( A0 => n335, B0 => n341, CI => n1110, CO => 
                           n332, S0 => n333);
   U315 : HS65_LH_FA1X4 port map( A0 => n2648, B0 => n1048, CI => n1078, CO => 
                           n334, S0 => n335);
   U317 : HS65_LH_FA1X4 port map( A0 => n1143, B0 => n340, CI => n346, CO => 
                           n337, S0 => n338);
   U318 : HS65_LH_FA1X4 port map( A0 => n348, B0 => n342, CI => n1111, CO => 
                           n339, S0 => n340);
   U319 : HS65_LH_FA1X4 port map( A0 => n1079, B0 => n343, CI => n350, CO => 
                           n341, S0 => n342);
   U320 : HS65_LH_FA1X4 port map( A0 => n352, B0 => n2640, CI => n1049, CO => 
                           n328, S0 => n343);
   U321 : HS65_LH_FA1X4 port map( A0 => n1176, B0 => n1144, CI => n347, CO => 
                           n344, S0 => n345);
   U322 : HS65_LH_FA1X4 port map( A0 => n349, B0 => n358, CI => n356, CO => 
                           n346, S0 => n347);
   U323 : HS65_LH_FA1X4 port map( A0 => n351, B0 => n1080, CI => n1112, CO => 
                           n348, S0 => n349);
   U324 : HS65_LH_FA1X4 port map( A0 => n1050, B0 => n2653, CI => n360, CO => 
                           n350, S0 => n351);
   U326 : HS65_LH_FA1X4 port map( A0 => n357, B0 => n365, CI => n1177, CO => 
                           n354, S0 => n355);
   U327 : HS65_LH_FA1X4 port map( A0 => n359, B0 => n367, CI => n1145, CO => 
                           n356, S0 => n357);
   U328 : HS65_LH_FA1X4 port map( A0 => n361, B0 => n369, CI => n1113, CO => 
                           n358, S0 => n359);
   U329 : HS65_LH_FA1X4 port map( A0 => n2653, B0 => n371, CI => n1081, CO => 
                           n360, S0 => n361);
   U331 : HS65_LH_FA1X4 port map( A0 => n1178, B0 => n366, CI => n375, CO => 
                           n363, S0 => n364);
   U332 : HS65_LH_FA1X4 port map( A0 => n377, B0 => n368, CI => n1146, CO => 
                           n365, S0 => n366);
   U333 : HS65_LH_FA1X4 port map( A0 => n1114, B0 => n370, CI => n379, CO => 
                           n367, S0 => n368);
   U334 : HS65_LH_FA1X4 port map( A0 => n381, B0 => n372, CI => n1082, CO => 
                           n369, S0 => n370);
   U335 : HS65_LH_FA1X4 port map( A0 => n383, B0 => n2638, CI => n1051, CO => 
                           n371, S0 => n372);
   U336 : HS65_LH_FA1X4 port map( A0 => n1211, B0 => n1179, CI => n376, CO => 
                           n373, S0 => n374);
   U337 : HS65_LH_FA1X4 port map( A0 => n378, B0 => n389, CI => n387, CO => 
                           n375, S0 => n376);
   U338 : HS65_LH_FA1X4 port map( A0 => n380, B0 => n1115, CI => n1147, CO => 
                           n377, S0 => n378);
   U339 : HS65_LH_FA1X4 port map( A0 => n382, B0 => n393, CI => n391, CO => 
                           n379, S0 => n380);
   U340 : HS65_LH_FA1X4 port map( A0 => n1052, B0 => n2649, CI => n1083, CO => 
                           n381, S0 => n382);
   U342 : HS65_LH_FA1X4 port map( A0 => n388, B0 => n398, CI => n1212, CO => 
                           n385, S0 => n386);
   U343 : HS65_LH_FA1X4 port map( A0 => n390, B0 => n400, CI => n1180, CO => 
                           n387, S0 => n388);
   U344 : HS65_LH_FA1X4 port map( A0 => n392, B0 => n402, CI => n1148, CO => 
                           n389, S0 => n390);
   U345 : HS65_LH_FA1X4 port map( A0 => n394, B0 => n404, CI => n1116, CO => 
                           n391, S0 => n392);
   U346 : HS65_LH_FA1X4 port map( A0 => n2649, B0 => n1053, CI => n1084, CO => 
                           n393, S0 => n394);
   U348 : HS65_LH_FA1X4 port map( A0 => n1213, B0 => n399, CI => n409, CO => 
                           n396, S0 => n397);
   U349 : HS65_LH_FA1X4 port map( A0 => n411, B0 => n401, CI => n1181, CO => 
                           n398, S0 => n399);
   U350 : HS65_LH_FA1X4 port map( A0 => n1149, B0 => n403, CI => n413, CO => 
                           n400, S0 => n401);
   U351 : HS65_LH_FA1X4 port map( A0 => n415, B0 => n405, CI => n1117, CO => 
                           n402, S0 => n403);
   U352 : HS65_LH_FA1X4 port map( A0 => n1085, B0 => n406, CI => n417, CO => 
                           n404, S0 => n405);
   U353 : HS65_LH_FA1X4 port map( A0 => n419, B0 => n2636, CI => n1054, CO => 
                           n383, S0 => n406);
   U354 : HS65_LH_FA1X4 port map( A0 => n1246, B0 => n1214, CI => n410, CO => 
                           n407, S0 => n408);
   U355 : HS65_LH_FA1X4 port map( A0 => n412, B0 => n425, CI => n423, CO => 
                           n409, S0 => n410);
   U356 : HS65_LH_FA1X4 port map( A0 => n414, B0 => n1150, CI => n1182, CO => 
                           n411, S0 => n412);
   U357 : HS65_LH_FA1X4 port map( A0 => n416, B0 => n429, CI => n427, CO => 
                           n413, S0 => n414);
   U358 : HS65_LH_FA1X4 port map( A0 => n418, B0 => n1086, CI => n1118, CO => 
                           n415, S0 => n416);
   U359 : HS65_LH_FA1X4 port map( A0 => n1055, B0 => n2654, CI => n431, CO => 
                           n417, S0 => n418);
   U361 : HS65_LH_FA1X4 port map( A0 => n424, B0 => n436, CI => n1247, CO => 
                           n421, S0 => n422);
   U362 : HS65_LH_FA1X4 port map( A0 => n426, B0 => n438, CI => n1215, CO => 
                           n423, S0 => n424);
   U363 : HS65_LH_FA1X4 port map( A0 => n428, B0 => n440, CI => n1183, CO => 
                           n425, S0 => n426);
   U364 : HS65_LH_FA1X4 port map( A0 => n430, B0 => n442, CI => n1151, CO => 
                           n427, S0 => n428);
   U365 : HS65_LH_FA1X4 port map( A0 => n432, B0 => n444, CI => n1119, CO => 
                           n429, S0 => n430);
   U366 : HS65_LH_FA1X4 port map( A0 => n2654, B0 => n446, CI => n1087, CO => 
                           n431, S0 => n432);
   U368 : HS65_LH_FA1X4 port map( A0 => n1248, B0 => n437, CI => n450, CO => 
                           n434, S0 => n435);
   U369 : HS65_LH_FA1X4 port map( A0 => n452, B0 => n439, CI => n1216, CO => 
                           n436, S0 => n437);
   U370 : HS65_LH_FA1X4 port map( A0 => n1184, B0 => n441, CI => n454, CO => 
                           n438, S0 => n439);
   U371 : HS65_LH_FA1X4 port map( A0 => n456, B0 => n443, CI => n1152, CO => 
                           n440, S0 => n441);
   U372 : HS65_LH_FA1X4 port map( A0 => n1120, B0 => n445, CI => n458, CO => 
                           n442, S0 => n443);
   U373 : HS65_LH_FA1X4 port map( A0 => n460, B0 => n447, CI => n1088, CO => 
                           n444, S0 => n445);
   U374 : HS65_LH_FA1X4 port map( A0 => n462, B0 => n2634, CI => n1056, CO => 
                           n446, S0 => n447);
   U375 : HS65_LH_FA1X4 port map( A0 => n1281, B0 => n1249, CI => n451, CO => 
                           n448, S0 => n449);
   U376 : HS65_LH_FA1X4 port map( A0 => n453, B0 => n468, CI => n466, CO => 
                           n450, S0 => n451);
   U377 : HS65_LH_FA1X4 port map( A0 => n455, B0 => n1185, CI => n1217, CO => 
                           n452, S0 => n453);
   U378 : HS65_LH_FA1X4 port map( A0 => n457, B0 => n472, CI => n470, CO => 
                           n454, S0 => n455);
   U379 : HS65_LH_FA1X4 port map( A0 => n459, B0 => n1121, CI => n1153, CO => 
                           n456, S0 => n457);
   U380 : HS65_LH_FA1X4 port map( A0 => n461, B0 => n476, CI => n474, CO => 
                           n458, S0 => n459);
   U381 : HS65_LH_FA1X4 port map( A0 => n1057, B0 => n2650, CI => n1089, CO => 
                           n460, S0 => n461);
   U383 : HS65_LH_FA1X4 port map( A0 => n467, B0 => n481, CI => n1282, CO => 
                           n464, S0 => n465);
   U384 : HS65_LH_FA1X4 port map( A0 => n469, B0 => n483, CI => n1250, CO => 
                           n466, S0 => n467);
   U385 : HS65_LH_FA1X4 port map( A0 => n471, B0 => n485, CI => n1218, CO => 
                           n468, S0 => n469);
   U386 : HS65_LH_FA1X4 port map( A0 => n473, B0 => n487, CI => n1186, CO => 
                           n470, S0 => n471);
   U387 : HS65_LH_FA1X4 port map( A0 => n475, B0 => n489, CI => n1154, CO => 
                           n472, S0 => n473);
   U388 : HS65_LH_FA1X4 port map( A0 => n477, B0 => n491, CI => n1122, CO => 
                           n474, S0 => n475);
   U389 : HS65_LH_FA1X4 port map( A0 => n2650, B0 => n1058, CI => n1090, CO => 
                           n476, S0 => n477);
   U391 : HS65_LH_FA1X4 port map( A0 => n1283, B0 => n482, CI => n496, CO => 
                           n479, S0 => n480);
   U392 : HS65_LH_FA1X4 port map( A0 => n498, B0 => n484, CI => n1251, CO => 
                           n481, S0 => n482);
   U393 : HS65_LH_FA1X4 port map( A0 => n1219, B0 => n486, CI => n500, CO => 
                           n483, S0 => n484);
   U394 : HS65_LH_FA1X4 port map( A0 => n502, B0 => n488, CI => n1187, CO => 
                           n485, S0 => n486);
   U395 : HS65_LH_FA1X4 port map( A0 => n1155, B0 => n490, CI => n504, CO => 
                           n487, S0 => n488);
   U396 : HS65_LH_FA1X4 port map( A0 => n506, B0 => n492, CI => n1123, CO => 
                           n489, S0 => n490);
   U397 : HS65_LH_FA1X4 port map( A0 => n1091, B0 => n493, CI => n508, CO => 
                           n491, S0 => n492);
   U398 : HS65_LH_FA1X4 port map( A0 => n510, B0 => n2632, CI => n1059, CO => 
                           n462, S0 => n493);
   U399 : HS65_LH_FA1X4 port map( A0 => n1316, B0 => n1284, CI => n497, CO => 
                           n494, S0 => n495);
   U400 : HS65_LH_FA1X4 port map( A0 => n499, B0 => n516, CI => n514, CO => 
                           n496, S0 => n497);
   U401 : HS65_LH_FA1X4 port map( A0 => n501, B0 => n1220, CI => n1252, CO => 
                           n498, S0 => n499);
   U402 : HS65_LH_FA1X4 port map( A0 => n503, B0 => n520, CI => n518, CO => 
                           n500, S0 => n501);
   U403 : HS65_LH_FA1X4 port map( A0 => n505, B0 => n1156, CI => n1188, CO => 
                           n502, S0 => n503);
   U404 : HS65_LH_FA1X4 port map( A0 => n507, B0 => n524, CI => n522, CO => 
                           n504, S0 => n505);
   U405 : HS65_LH_FA1X4 port map( A0 => n509, B0 => n1092, CI => n1124, CO => 
                           n506, S0 => n507);
   U406 : HS65_LH_FA1X4 port map( A0 => n1060, B0 => n2651, CI => n526, CO => 
                           n508, S0 => n509);
   U408 : HS65_LH_FA1X4 port map( A0 => n515, B0 => n531, CI => n1317, CO => 
                           n512, S0 => n513);
   U409 : HS65_LH_FA1X4 port map( A0 => n517, B0 => n533, CI => n1285, CO => 
                           n514, S0 => n515);
   U410 : HS65_LH_FA1X4 port map( A0 => n519, B0 => n535, CI => n1253, CO => 
                           n516, S0 => n517);
   U411 : HS65_LH_FA1X4 port map( A0 => n521, B0 => n537, CI => n1221, CO => 
                           n518, S0 => n519);
   U412 : HS65_LH_FA1X4 port map( A0 => n523, B0 => n539, CI => n1189, CO => 
                           n520, S0 => n521);
   U413 : HS65_LH_FA1X4 port map( A0 => n525, B0 => n541, CI => n1157, CO => 
                           n522, S0 => n523);
   U414 : HS65_LH_FA1X4 port map( A0 => n527, B0 => n543, CI => n1125, CO => 
                           n524, S0 => n525);
   U415 : HS65_LH_FA1X4 port map( A0 => n2651, B0 => n1061, CI => n1093, CO => 
                           n526, S0 => n527);
   U417 : HS65_LH_FA1X4 port map( A0 => n1318, B0 => n532, CI => n548, CO => 
                           n529, S0 => n530);
   U418 : HS65_LH_FA1X4 port map( A0 => n550, B0 => n534, CI => n1286, CO => 
                           n531, S0 => n532);
   U419 : HS65_LH_FA1X4 port map( A0 => n1254, B0 => n536, CI => n552, CO => 
                           n533, S0 => n534);
   U420 : HS65_LH_FA1X4 port map( A0 => n554, B0 => n538, CI => n1222, CO => 
                           n535, S0 => n536);
   U421 : HS65_LH_FA1X4 port map( A0 => n1190, B0 => n540, CI => n556, CO => 
                           n537, S0 => n538);
   U422 : HS65_LH_FA1X4 port map( A0 => n1158, B0 => n542, CI => n558, CO => 
                           n539, S0 => n540);
   U423 : HS65_LH_FA1X4 port map( A0 => n1126, B0 => n544, CI => n560, CO => 
                           n541, S0 => n542);
   U424 : HS65_LH_FA1X4 port map( A0 => n562, B0 => n545, CI => n1094, CO => 
                           n543, S0 => n544);
   U425 : HS65_LH_FA1X4 port map( A0 => n2630, B0 => n2628, CI => n1062, CO => 
                           n510, S0 => n545);
   U426 : HS65_LH_FA1X4 port map( A0 => n1351, B0 => n1319, CI => n549, CO => 
                           n546, S0 => n547);
   U427 : HS65_LH_FA1X4 port map( A0 => n551, B0 => n1287, CI => n566, CO => 
                           n548, S0 => n549);
   U428 : HS65_LH_FA1X4 port map( A0 => n553, B0 => n1255, CI => n568, CO => 
                           n550, S0 => n551);
   U429 : HS65_LH_FA1X4 port map( A0 => n555, B0 => n572, CI => n570, CO => 
                           n552, S0 => n553);
   U430 : HS65_LH_FA1X4 port map( A0 => n557, B0 => n1191, CI => n1223, CO => 
                           n554, S0 => n555);
   U431 : HS65_LH_FA1X4 port map( A0 => n559, B0 => n576, CI => n574, CO => 
                           n556, S0 => n557);
   U432 : HS65_LH_FA1X4 port map( A0 => n561, B0 => n1127, CI => n1159, CO => 
                           n558, S0 => n559);
   U433 : HS65_LH_FA1X4 port map( A0 => n563, B0 => n1095, CI => n578, CO => 
                           n560, S0 => n561);
   U434 : HS65_LH_FA1X4 port map( A0 => n1063, B0 => a(2), CI => n580, CO => 
                           n562, S0 => n563);
   U435 : HS65_LH_FA1X4 port map( A0 => n567, B0 => n1320, CI => n1352, CO => 
                           n564, S0 => n565);
   U436 : HS65_LH_FA1X4 port map( A0 => n569, B0 => n1288, CI => n584, CO => 
                           n566, S0 => n567);
   U437 : HS65_LH_FA1X4 port map( A0 => n571, B0 => n1256, CI => n586, CO => 
                           n568, S0 => n569);
   U438 : HS65_LH_FA1X4 port map( A0 => n573, B0 => n590, CI => n588, CO => 
                           n570, S0 => n571);
   U439 : HS65_LH_FA1X4 port map( A0 => n575, B0 => n1192, CI => n1224, CO => 
                           n572, S0 => n573);
   U440 : HS65_LH_FA1X4 port map( A0 => n577, B0 => n594, CI => n592, CO => 
                           n574, S0 => n575);
   U441 : HS65_LH_FA1X4 port map( A0 => n579, B0 => n1128, CI => n1160, CO => 
                           n576, S0 => n577);
   U442 : HS65_LH_FA1X4 port map( A0 => n581, B0 => n1096, CI => n596, CO => 
                           n578, S0 => n579);
   U443 : HS65_LH_FA1X4 port map( A0 => n1064, B0 => a(2), CI => n598, CO => 
                           n580, S0 => n581);
   U444 : HS65_LH_FA1X4 port map( A0 => n585, B0 => n602, CI => n1353, CO => 
                           n582, S0 => n583);
   U445 : HS65_LH_FA1X4 port map( A0 => n587, B0 => n604, CI => n1321, CO => 
                           n584, S0 => n585);
   U446 : HS65_LH_FA1X4 port map( A0 => n589, B0 => n606, CI => n1289, CO => 
                           n586, S0 => n587);
   U447 : HS65_LH_FA1X4 port map( A0 => n591, B0 => n608, CI => n1257, CO => 
                           n588, S0 => n589);
   U448 : HS65_LH_FA1X4 port map( A0 => n593, B0 => n610, CI => n1225, CO => 
                           n590, S0 => n591);
   U449 : HS65_LH_FA1X4 port map( A0 => n595, B0 => n612, CI => n1193, CO => 
                           n592, S0 => n593);
   U450 : HS65_LH_FA1X4 port map( A0 => n597, B0 => n614, CI => n1161, CO => 
                           n594, S0 => n595);
   U451 : HS65_LH_FA1X4 port map( A0 => n599, B0 => n616, CI => n1129, CO => 
                           n596, S0 => n597);
   U452 : HS65_LH_FA1X4 port map( A0 => n1065, B0 => a(2), CI => n1097, CO => 
                           n598, S0 => n599);
   U453 : HS65_LH_FA1X4 port map( A0 => n1354, B0 => n603, CI => n618, CO => 
                           n600, S0 => n601);
   U454 : HS65_LH_FA1X4 port map( A0 => n1322, B0 => n605, CI => n620, CO => 
                           n602, S0 => n603);
   U455 : HS65_LH_FA1X4 port map( A0 => n1290, B0 => n607, CI => n622, CO => 
                           n604, S0 => n605);
   U456 : HS65_LH_FA1X4 port map( A0 => n1258, B0 => n609, CI => n624, CO => 
                           n606, S0 => n607);
   U457 : HS65_LH_FA1X4 port map( A0 => n1226, B0 => n611, CI => n626, CO => 
                           n608, S0 => n609);
   U458 : HS65_LH_FA1X4 port map( A0 => n1194, B0 => n613, CI => n628, CO => 
                           n610, S0 => n611);
   U459 : HS65_LH_FA1X4 port map( A0 => n1162, B0 => n615, CI => n630, CO => 
                           n612, S0 => n613);
   U460 : HS65_LH_FA1X4 port map( A0 => n1130, B0 => n617, CI => n632, CO => 
                           n614, S0 => n615);
   U461 : HS65_LH_FA1X4 port map( A0 => n1098, B0 => n1066, CI => n634, CO => 
                           n616, S0 => n617);
   U462 : HS65_LH_FA1X4 port map( A0 => n1355, B0 => n621, CI => n636, CO => 
                           n618, S0 => n619);
   U463 : HS65_LH_FA1X4 port map( A0 => n1323, B0 => n623, CI => n638, CO => 
                           n620, S0 => n621);
   U464 : HS65_LH_FA1X4 port map( A0 => n1291, B0 => n625, CI => n640, CO => 
                           n622, S0 => n623);
   U465 : HS65_LH_FA1X4 port map( A0 => n1259, B0 => n627, CI => n642, CO => 
                           n624, S0 => n625);
   U466 : HS65_LH_FA1X4 port map( A0 => n1227, B0 => n629, CI => n644, CO => 
                           n626, S0 => n627);
   U467 : HS65_LH_FA1X4 port map( A0 => n1195, B0 => n631, CI => n646, CO => 
                           n628, S0 => n629);
   U468 : HS65_LH_FA1X4 port map( A0 => n1163, B0 => n633, CI => n648, CO => 
                           n630, S0 => n631);
   U469 : HS65_LH_FA1X4 port map( A0 => n1131, B0 => n635, CI => n650, CO => 
                           n632, S0 => n633);
   U470 : HS65_LH_FA1X4 port map( A0 => n1099, B0 => n1067, CI => n652, CO => 
                           n634, S0 => n635);
   U471 : HS65_LH_FA1X4 port map( A0 => n1356, B0 => n639, CI => n654, CO => 
                           n636, S0 => n637);
   U472 : HS65_LH_FA1X4 port map( A0 => n1324, B0 => n641, CI => n656, CO => 
                           n638, S0 => n639);
   U473 : HS65_LH_FA1X4 port map( A0 => n1292, B0 => n643, CI => n658, CO => 
                           n640, S0 => n641);
   U474 : HS65_LH_FA1X4 port map( A0 => n1260, B0 => n645, CI => n660, CO => 
                           n642, S0 => n643);
   U475 : HS65_LH_FA1X4 port map( A0 => n1228, B0 => n647, CI => n662, CO => 
                           n644, S0 => n645);
   U476 : HS65_LH_FA1X4 port map( A0 => n1196, B0 => n649, CI => n664, CO => 
                           n646, S0 => n647);
   U477 : HS65_LH_FA1X4 port map( A0 => n1164, B0 => n651, CI => n666, CO => 
                           n648, S0 => n649);
   U478 : HS65_LH_FA1X4 port map( A0 => n1132, B0 => n653, CI => n668, CO => 
                           n650, S0 => n651);
   U479 : HS65_LH_FA1X4 port map( A0 => n1100, B0 => n1068, CI => n670, CO => 
                           n652, S0 => n653);
   U480 : HS65_LH_FA1X4 port map( A0 => n1357, B0 => n657, CI => n672, CO => 
                           n654, S0 => n655);
   U481 : HS65_LH_FA1X4 port map( A0 => n1325, B0 => n659, CI => n674, CO => 
                           n656, S0 => n657);
   U482 : HS65_LH_FA1X4 port map( A0 => n1293, B0 => n661, CI => n676, CO => 
                           n658, S0 => n659);
   U483 : HS65_LH_FA1X4 port map( A0 => n1261, B0 => n663, CI => n678, CO => 
                           n660, S0 => n661);
   U484 : HS65_LH_FA1X4 port map( A0 => n1229, B0 => n665, CI => n680, CO => 
                           n662, S0 => n663);
   U485 : HS65_LH_FA1X4 port map( A0 => n1197, B0 => n667, CI => n682, CO => 
                           n664, S0 => n665);
   U486 : HS65_LH_FA1X4 port map( A0 => n1165, B0 => n669, CI => n684, CO => 
                           n666, S0 => n667);
   U487 : HS65_LH_FA1X4 port map( A0 => n1133, B0 => n671, CI => n686, CO => 
                           n668, S0 => n669);
   U488 : HS65_LH_FA1X4 port map( A0 => n1101, B0 => n1069, CI => n688, CO => 
                           n670, S0 => n671);
   U489 : HS65_LH_FA1X4 port map( A0 => n1358, B0 => n675, CI => n690, CO => 
                           n672, S0 => n673);
   U490 : HS65_LH_FA1X4 port map( A0 => n1326, B0 => n677, CI => n692, CO => 
                           n674, S0 => n675);
   U491 : HS65_LH_FA1X4 port map( A0 => n1294, B0 => n679, CI => n694, CO => 
                           n676, S0 => n677);
   U492 : HS65_LH_FA1X4 port map( A0 => n1262, B0 => n681, CI => n696, CO => 
                           n678, S0 => n679);
   U493 : HS65_LH_FA1X4 port map( A0 => n1230, B0 => n683, CI => n698, CO => 
                           n680, S0 => n681);
   U494 : HS65_LH_FA1X4 port map( A0 => n1198, B0 => n685, CI => n700, CO => 
                           n682, S0 => n683);
   U495 : HS65_LH_FA1X4 port map( A0 => n1166, B0 => n687, CI => n702, CO => 
                           n684, S0 => n685);
   U496 : HS65_LH_FA1X4 port map( A0 => n1134, B0 => n689, CI => n704, CO => 
                           n686, S0 => n687);
   U497 : HS65_LH_HA1X4 port map( A0 => n1102, B0 => n706, CO => n688, S0 => 
                           n689);
   U498 : HS65_LH_FA1X4 port map( A0 => n1359, B0 => n693, CI => n708, CO => 
                           n690, S0 => n691);
   U499 : HS65_LH_FA1X4 port map( A0 => n1327, B0 => n695, CI => n710, CO => 
                           n692, S0 => n693);
   U500 : HS65_LH_FA1X4 port map( A0 => n1295, B0 => n697, CI => n712, CO => 
                           n694, S0 => n695);
   U501 : HS65_LH_FA1X4 port map( A0 => n1263, B0 => n699, CI => n714, CO => 
                           n696, S0 => n697);
   U502 : HS65_LH_FA1X4 port map( A0 => n1231, B0 => n701, CI => n716, CO => 
                           n698, S0 => n699);
   U503 : HS65_LH_FA1X4 port map( A0 => n1199, B0 => n703, CI => n718, CO => 
                           n700, S0 => n701);
   U504 : HS65_LH_FA1X4 port map( A0 => n1167, B0 => n705, CI => n720, CO => 
                           n702, S0 => n703);
   U505 : HS65_LH_FA1X4 port map( A0 => n1135, B0 => n707, CI => n722, CO => 
                           n704, S0 => n705);
   U506 : HS65_LH_HA1X4 port map( A0 => n1103, B0 => n724, CO => n706, S0 => 
                           n707);
   U507 : HS65_LH_FA1X4 port map( A0 => n1360, B0 => n711, CI => n726, CO => 
                           n708, S0 => n709);
   U508 : HS65_LH_FA1X4 port map( A0 => n1328, B0 => n713, CI => n728, CO => 
                           n710, S0 => n711);
   U509 : HS65_LH_FA1X4 port map( A0 => n1296, B0 => n715, CI => n730, CO => 
                           n712, S0 => n713);
   U510 : HS65_LH_FA1X4 port map( A0 => n1264, B0 => n717, CI => n732, CO => 
                           n714, S0 => n715);
   U511 : HS65_LH_FA1X4 port map( A0 => n1232, B0 => n719, CI => n734, CO => 
                           n716, S0 => n717);
   U512 : HS65_LH_FA1X4 port map( A0 => n1200, B0 => n721, CI => n736, CO => 
                           n718, S0 => n719);
   U513 : HS65_LH_FA1X4 port map( A0 => n1168, B0 => n723, CI => n738, CO => 
                           n720, S0 => n721);
   U514 : HS65_LH_FA1X4 port map( A0 => n1136, B0 => n725, CI => n740, CO => 
                           n722, S0 => n723);
   U515 : HS65_LH_HA1X4 port map( A0 => n2645, B0 => n1104, CO => n724, S0 => 
                           n725);
   U516 : HS65_LH_FA1X4 port map( A0 => n1361, B0 => n729, CI => n742, CO => 
                           n726, S0 => n727);
   U517 : HS65_LH_FA1X4 port map( A0 => n1329, B0 => n731, CI => n744, CO => 
                           n728, S0 => n729);
   U518 : HS65_LH_FA1X4 port map( A0 => n1297, B0 => n733, CI => n746, CO => 
                           n730, S0 => n731);
   U519 : HS65_LH_FA1X4 port map( A0 => n1265, B0 => n735, CI => n748, CO => 
                           n732, S0 => n733);
   U520 : HS65_LH_FA1X4 port map( A0 => n1233, B0 => n737, CI => n750, CO => 
                           n734, S0 => n735);
   U521 : HS65_LH_FA1X4 port map( A0 => n1201, B0 => n739, CI => n752, CO => 
                           n736, S0 => n737);
   U522 : HS65_LH_FA1X4 port map( A0 => n1169, B0 => n741, CI => n754, CO => 
                           n738, S0 => n739);
   U523 : HS65_LH_HA1X4 port map( A0 => n1137, B0 => n756, CO => n740, S0 => 
                           n741);
   U524 : HS65_LH_FA1X4 port map( A0 => n1362, B0 => n745, CI => n758, CO => 
                           n742, S0 => n743);
   U525 : HS65_LH_FA1X4 port map( A0 => n1330, B0 => n747, CI => n760, CO => 
                           n744, S0 => n745);
   U526 : HS65_LH_FA1X4 port map( A0 => n1298, B0 => n749, CI => n762, CO => 
                           n746, S0 => n747);
   U527 : HS65_LH_FA1X4 port map( A0 => n1266, B0 => n751, CI => n764, CO => 
                           n748, S0 => n749);
   U528 : HS65_LH_FA1X4 port map( A0 => n1234, B0 => n753, CI => n766, CO => 
                           n750, S0 => n751);
   U529 : HS65_LH_FA1X4 port map( A0 => n1202, B0 => n755, CI => n768, CO => 
                           n752, S0 => n753);
   U530 : HS65_LH_FA1X4 port map( A0 => n1170, B0 => n757, CI => n770, CO => 
                           n754, S0 => n755);
   U531 : HS65_LH_HA1X4 port map( A0 => n1138, B0 => n772, CO => n756, S0 => 
                           n757);
   U532 : HS65_LH_FA1X4 port map( A0 => n1363, B0 => n761, CI => n774, CO => 
                           n758, S0 => n759);
   U533 : HS65_LH_FA1X4 port map( A0 => n1331, B0 => n763, CI => n776, CO => 
                           n760, S0 => n761);
   U534 : HS65_LH_FA1X4 port map( A0 => n1299, B0 => n765, CI => n778, CO => 
                           n762, S0 => n763);
   U535 : HS65_LH_FA1X4 port map( A0 => n1267, B0 => n767, CI => n780, CO => 
                           n764, S0 => n765);
   U536 : HS65_LH_FA1X4 port map( A0 => n1235, B0 => n769, CI => n782, CO => 
                           n766, S0 => n767);
   U537 : HS65_LH_FA1X4 port map( A0 => n1203, B0 => n771, CI => n784, CO => 
                           n768, S0 => n769);
   U538 : HS65_LH_FA1X4 port map( A0 => n1171, B0 => n773, CI => n786, CO => 
                           n770, S0 => n771);
   U539 : HS65_LH_HA1X4 port map( A0 => a(26), B0 => n1139, CO => n772, S0 => 
                           n773);
   U540 : HS65_LH_FA1X4 port map( A0 => n1364, B0 => n777, CI => n788, CO => 
                           n774, S0 => n775);
   U541 : HS65_LH_FA1X4 port map( A0 => n1332, B0 => n779, CI => n790, CO => 
                           n776, S0 => n777);
   U542 : HS65_LH_FA1X4 port map( A0 => n1300, B0 => n781, CI => n792, CO => 
                           n778, S0 => n779);
   U543 : HS65_LH_FA1X4 port map( A0 => n1268, B0 => n783, CI => n794, CO => 
                           n780, S0 => n781);
   U544 : HS65_LH_FA1X4 port map( A0 => n1236, B0 => n785, CI => n796, CO => 
                           n782, S0 => n783);
   U545 : HS65_LH_FA1X4 port map( A0 => n1204, B0 => n787, CI => n798, CO => 
                           n784, S0 => n785);
   U546 : HS65_LH_HA1X4 port map( A0 => n1172, B0 => n800, CO => n786, S0 => 
                           n787);
   U547 : HS65_LH_FA1X4 port map( A0 => n1365, B0 => n791, CI => n802, CO => 
                           n788, S0 => n789);
   U548 : HS65_LH_FA1X4 port map( A0 => n1333, B0 => n793, CI => n804, CO => 
                           n790, S0 => n791);
   U549 : HS65_LH_FA1X4 port map( A0 => n1301, B0 => n795, CI => n806, CO => 
                           n792, S0 => n793);
   U550 : HS65_LH_FA1X4 port map( A0 => n1269, B0 => n797, CI => n808, CO => 
                           n794, S0 => n795);
   U551 : HS65_LH_FA1X4 port map( A0 => n1237, B0 => n799, CI => n810, CO => 
                           n796, S0 => n797);
   U552 : HS65_LH_FA1X4 port map( A0 => n1205, B0 => n801, CI => n812, CO => 
                           n798, S0 => n799);
   U553 : HS65_LH_HA1X4 port map( A0 => n1173, B0 => n814, CO => n800, S0 => 
                           n801);
   U554 : HS65_LH_FA1X4 port map( A0 => n1366, B0 => n805, CI => n816, CO => 
                           n802, S0 => n803);
   U555 : HS65_LH_FA1X4 port map( A0 => n1334, B0 => n807, CI => n818, CO => 
                           n804, S0 => n805);
   U556 : HS65_LH_FA1X4 port map( A0 => n1302, B0 => n809, CI => n820, CO => 
                           n806, S0 => n807);
   U557 : HS65_LH_FA1X4 port map( A0 => n1270, B0 => n811, CI => n822, CO => 
                           n808, S0 => n809);
   U558 : HS65_LH_FA1X4 port map( A0 => n1238, B0 => n813, CI => n824, CO => 
                           n810, S0 => n811);
   U559 : HS65_LH_FA1X4 port map( A0 => n1206, B0 => n815, CI => n826, CO => 
                           n812, S0 => n813);
   U560 : HS65_LH_HA1X4 port map( A0 => a(23), B0 => n1174, CO => n814, S0 => 
                           n815);
   U561 : HS65_LH_FA1X4 port map( A0 => n1367, B0 => n819, CI => n828, CO => 
                           n816, S0 => n817);
   U562 : HS65_LH_FA1X4 port map( A0 => n1335, B0 => n821, CI => n830, CO => 
                           n818, S0 => n819);
   U563 : HS65_LH_FA1X4 port map( A0 => n1303, B0 => n823, CI => n832, CO => 
                           n820, S0 => n821);
   U564 : HS65_LH_FA1X4 port map( A0 => n1271, B0 => n825, CI => n834, CO => 
                           n822, S0 => n823);
   U565 : HS65_LH_FA1X4 port map( A0 => n1239, B0 => n827, CI => n836, CO => 
                           n824, S0 => n825);
   U566 : HS65_LH_HA1X4 port map( A0 => n1207, B0 => n838, CO => n826, S0 => 
                           n827);
   U567 : HS65_LH_FA1X4 port map( A0 => n1368, B0 => n831, CI => n840, CO => 
                           n828, S0 => n829);
   U568 : HS65_LH_FA1X4 port map( A0 => n1336, B0 => n833, CI => n842, CO => 
                           n830, S0 => n831);
   U569 : HS65_LH_FA1X4 port map( A0 => n1304, B0 => n835, CI => n844, CO => 
                           n832, S0 => n833);
   U570 : HS65_LH_FA1X4 port map( A0 => n1272, B0 => n837, CI => n846, CO => 
                           n834, S0 => n835);
   U571 : HS65_LH_FA1X4 port map( A0 => n1240, B0 => n839, CI => n848, CO => 
                           n836, S0 => n837);
   U572 : HS65_LH_HA1X4 port map( A0 => n1208, B0 => n850, CO => n838, S0 => 
                           n839);
   U573 : HS65_LH_FA1X4 port map( A0 => n1369, B0 => n843, CI => n852, CO => 
                           n840, S0 => n841);
   U574 : HS65_LH_FA1X4 port map( A0 => n1337, B0 => n845, CI => n854, CO => 
                           n842, S0 => n843);
   U575 : HS65_LH_FA1X4 port map( A0 => n1305, B0 => n847, CI => n856, CO => 
                           n844, S0 => n845);
   U576 : HS65_LH_FA1X4 port map( A0 => n1273, B0 => n849, CI => n858, CO => 
                           n846, S0 => n847);
   U577 : HS65_LH_FA1X4 port map( A0 => n1241, B0 => n851, CI => n860, CO => 
                           n848, S0 => n849);
   U578 : HS65_LH_HA1X4 port map( A0 => a(20), B0 => n1209, CO => n850, S0 => 
                           n851);
   U579 : HS65_LH_FA1X4 port map( A0 => n1370, B0 => n855, CI => n862, CO => 
                           n852, S0 => n853);
   U580 : HS65_LH_FA1X4 port map( A0 => n1338, B0 => n857, CI => n864, CO => 
                           n854, S0 => n855);
   U581 : HS65_LH_FA1X4 port map( A0 => n1306, B0 => n859, CI => n866, CO => 
                           n856, S0 => n857);
   U582 : HS65_LH_FA1X4 port map( A0 => n1274, B0 => n861, CI => n868, CO => 
                           n858, S0 => n859);
   U583 : HS65_LH_HA1X4 port map( A0 => n1242, B0 => n870, CO => n860, S0 => 
                           n861);
   U584 : HS65_LH_FA1X4 port map( A0 => n1371, B0 => n865, CI => n872, CO => 
                           n862, S0 => n863);
   U585 : HS65_LH_FA1X4 port map( A0 => n1339, B0 => n867, CI => n874, CO => 
                           n864, S0 => n865);
   U586 : HS65_LH_FA1X4 port map( A0 => n1307, B0 => n869, CI => n876, CO => 
                           n866, S0 => n867);
   U587 : HS65_LH_FA1X4 port map( A0 => n1275, B0 => n871, CI => n878, CO => 
                           n868, S0 => n869);
   U588 : HS65_LH_HA1X4 port map( A0 => n1243, B0 => n880, CO => n870, S0 => 
                           n871);
   U589 : HS65_LH_FA1X4 port map( A0 => n1372, B0 => n875, CI => n882, CO => 
                           n872, S0 => n873);
   U590 : HS65_LH_FA1X4 port map( A0 => n1340, B0 => n877, CI => n884, CO => 
                           n874, S0 => n875);
   U591 : HS65_LH_FA1X4 port map( A0 => n1308, B0 => n879, CI => n886, CO => 
                           n876, S0 => n877);
   U592 : HS65_LH_FA1X4 port map( A0 => n1276, B0 => n881, CI => n888, CO => 
                           n878, S0 => n879);
   U593 : HS65_LH_HA1X4 port map( A0 => a(17), B0 => n1244, CO => n880, S0 => 
                           n881);
   U594 : HS65_LH_FA1X4 port map( A0 => n1373, B0 => n885, CI => n890, CO => 
                           n882, S0 => n883);
   U595 : HS65_LH_FA1X4 port map( A0 => n1341, B0 => n887, CI => n892, CO => 
                           n884, S0 => n885);
   U596 : HS65_LH_FA1X4 port map( A0 => n1309, B0 => n889, CI => n894, CO => 
                           n886, S0 => n887);
   U597 : HS65_LH_HA1X4 port map( A0 => n1277, B0 => n896, CO => n888, S0 => 
                           n889);
   U598 : HS65_LH_FA1X4 port map( A0 => n1374, B0 => n893, CI => n898, CO => 
                           n890, S0 => n891);
   U599 : HS65_LH_FA1X4 port map( A0 => n1342, B0 => n895, CI => n900, CO => 
                           n892, S0 => n893);
   U600 : HS65_LH_FA1X4 port map( A0 => n1310, B0 => n897, CI => n902, CO => 
                           n894, S0 => n895);
   U601 : HS65_LH_HA1X4 port map( A0 => n1278, B0 => n904, CO => n896, S0 => 
                           n897);
   U602 : HS65_LH_FA1X4 port map( A0 => n1375, B0 => n901, CI => n906, CO => 
                           n898, S0 => n899);
   U603 : HS65_LH_FA1X4 port map( A0 => n1343, B0 => n903, CI => n908, CO => 
                           n900, S0 => n901);
   U604 : HS65_LH_FA1X4 port map( A0 => n1311, B0 => n905, CI => n910, CO => 
                           n902, S0 => n903);
   U605 : HS65_LH_HA1X4 port map( A0 => a(14), B0 => n1279, CO => n904, S0 => 
                           n905);
   U606 : HS65_LH_FA1X4 port map( A0 => n1376, B0 => n909, CI => n912, CO => 
                           n906, S0 => n907);
   U607 : HS65_LH_FA1X4 port map( A0 => n1344, B0 => n911, CI => n914, CO => 
                           n908, S0 => n909);
   U608 : HS65_LH_HA1X4 port map( A0 => n1312, B0 => n916, CO => n910, S0 => 
                           n911);
   U609 : HS65_LH_FA1X4 port map( A0 => n1377, B0 => n915, CI => n918, CO => 
                           n912, S0 => n913);
   U610 : HS65_LH_FA1X4 port map( A0 => n1345, B0 => n917, CI => n920, CO => 
                           n914, S0 => n915);
   U611 : HS65_LH_HA1X4 port map( A0 => n1313, B0 => n922, CO => n916, S0 => 
                           n917);
   U612 : HS65_LH_FA1X4 port map( A0 => n1378, B0 => n921, CI => n924, CO => 
                           n918, S0 => n919);
   U613 : HS65_LH_FA1X4 port map( A0 => n1346, B0 => n923, CI => n926, CO => 
                           n920, S0 => n921);
   U614 : HS65_LH_HA1X4 port map( A0 => a(11), B0 => n1314, CO => n922, S0 => 
                           n923);
   U615 : HS65_LH_FA1X4 port map( A0 => n1379, B0 => n927, CI => n928, CO => 
                           n924, S0 => n925);
   U616 : HS65_LH_HA1X4 port map( A0 => n1347, B0 => n930, CO => n926, S0 => 
                           n927);
   U617 : HS65_LH_FA1X4 port map( A0 => n1380, B0 => n931, CI => n932, CO => 
                           n928, S0 => n929);
   U618 : HS65_LH_HA1X4 port map( A0 => n1348, B0 => n934, CO => n930, S0 => 
                           n931);
   U619 : HS65_LH_FA1X4 port map( A0 => n1381, B0 => n935, CI => n936, CO => 
                           n932, S0 => n933);
   U620 : HS65_LH_HA1X4 port map( A0 => a(8), B0 => n1349, CO => n934, S0 => 
                           n935);
   U621 : HS65_LH_HA1X4 port map( A0 => n1382, B0 => n938, CO => n936, S0 => 
                           n937);
   U622 : HS65_LH_HA1X4 port map( A0 => n1383, B0 => n940, CO => n938, S0 => 
                           n939);
   U623 : HS65_LH_HA1X4 port map( A0 => a(5), B0 => n1384, CO => n940, S0 => 
                           n941);
   U1907 : HS65_LH_HA1X4 port map( A0 => n2626, B0 => n975, CO => n1006, S0 => 
                           n1007);
   U1908 : HS65_LH_FA1X4 port map( A0 => n2624, B0 => n2626, CI => n976, CO => 
                           n975, S0 => n1008);
   U1909 : HS65_LH_FA1X4 port map( A0 => n2622, B0 => n2624, CI => n977, CO => 
                           n976, S0 => n1009);
   U1910 : HS65_LH_FA1X4 port map( A0 => n2620, B0 => n2622, CI => n978, CO => 
                           n977, S0 => n1010);
   U1911 : HS65_LH_FA1X4 port map( A0 => n2618, B0 => n2620, CI => n979, CO => 
                           n978, S0 => n1011);
   U1912 : HS65_LH_FA1X4 port map( A0 => n2616, B0 => n2618, CI => n980, CO => 
                           n979, S0 => n1012);
   U1913 : HS65_LH_FA1X4 port map( A0 => n2614, B0 => n2616, CI => n981, CO => 
                           n980, S0 => n1013);
   U1914 : HS65_LH_FA1X4 port map( A0 => n2612, B0 => n2614, CI => n982, CO => 
                           n981, S0 => n1014);
   U1915 : HS65_LH_FA1X4 port map( A0 => n2610, B0 => n2612, CI => n983, CO => 
                           n982, S0 => n1015);
   U1916 : HS65_LH_FA1X4 port map( A0 => n2608, B0 => n2610, CI => n984, CO => 
                           n983, S0 => n1016);
   U1917 : HS65_LH_FA1X4 port map( A0 => n2606, B0 => n2608, CI => n985, CO => 
                           n984, S0 => n1017);
   U1918 : HS65_LH_FA1X4 port map( A0 => n2604, B0 => n2606, CI => n986, CO => 
                           n985, S0 => n1018);
   U1919 : HS65_LH_FA1X4 port map( A0 => n2602, B0 => n2604, CI => n987, CO => 
                           n986, S0 => n1019);
   U1920 : HS65_LH_FA1X4 port map( A0 => n2600, B0 => n2602, CI => n988, CO => 
                           n987, S0 => n1020);
   U1921 : HS65_LH_FA1X4 port map( A0 => n2598, B0 => n2600, CI => n989, CO => 
                           n988, S0 => n1021);
   U1922 : HS65_LH_FA1X4 port map( A0 => n2596, B0 => n2598, CI => n990, CO => 
                           n989, S0 => n1022);
   U1923 : HS65_LH_FA1X4 port map( A0 => n2594, B0 => n2596, CI => n991, CO => 
                           n990, S0 => n1023);
   U1924 : HS65_LH_FA1X4 port map( A0 => n2592, B0 => n2594, CI => n992, CO => 
                           n991, S0 => n1024);
   U1925 : HS65_LH_FA1X4 port map( A0 => n2590, B0 => n2592, CI => n993, CO => 
                           n992, S0 => n1025);
   U1926 : HS65_LH_FA1X4 port map( A0 => n2588, B0 => n2590, CI => n994, CO => 
                           n993, S0 => n1026);
   U1927 : HS65_LH_FA1X4 port map( A0 => n2586, B0 => n2588, CI => n995, CO => 
                           n994, S0 => n1027);
   U1928 : HS65_LH_FA1X4 port map( A0 => n2584, B0 => n2586, CI => n996, CO => 
                           n995, S0 => n1028);
   U1929 : HS65_LH_FA1X4 port map( A0 => n2582, B0 => n2584, CI => n997, CO => 
                           n996, S0 => n1029);
   U1930 : HS65_LH_FA1X4 port map( A0 => n2580, B0 => n2582, CI => n998, CO => 
                           n997, S0 => n1030);
   U1931 : HS65_LH_FA1X4 port map( A0 => n2578, B0 => n2580, CI => n999, CO => 
                           n998, S0 => n1031);
   U1932 : HS65_LH_FA1X4 port map( A0 => n2576, B0 => n2578, CI => n1000, CO =>
                           n999, S0 => n1032);
   U1933 : HS65_LH_FA1X4 port map( A0 => n2574, B0 => n2576, CI => n1001, CO =>
                           n1000, S0 => n1033);
   U1934 : HS65_LH_FA1X4 port map( A0 => n2572, B0 => n2574, CI => n1002, CO =>
                           n1001, S0 => n1034);
   U1935 : HS65_LH_FA1X4 port map( A0 => n2570, B0 => n2572, CI => n1003, CO =>
                           n1002, S0 => n1035);
   U1936 : HS65_LH_FA1X4 port map( A0 => n2568, B0 => n2570, CI => n1004, CO =>
                           n1003, S0 => n1036);
   U1937 : HS65_LH_FA1X4 port map( A0 => n2566, B0 => n2568, CI => n1005, CO =>
                           n1004, S0 => n1037);
   U1941 : HS65_LH_IVX9 port map( A => a(2), Z => n2628);
   U1942 : HS65_LH_IVX9 port map( A => n1007, Z => n2657);
   U1943 : HS65_LH_IVX9 port map( A => n419, Z => n2654);
   U1944 : HS65_LH_IVX9 port map( A => n352, Z => n2653);
   U1945 : HS65_LH_IVX9 port map( A => n309, Z => n2652);
   U1946 : HS65_LH_IVX9 port map( A => n510, Z => n2651);
   U1947 : HS65_LH_IVX9 port map( A => n462, Z => n2650);
   U1948 : HS65_LH_IVX9 port map( A => n383, Z => n2649);
   U1949 : HS65_LH_IVX9 port map( A => n328, Z => n2648);
   U1950 : HS65_LH_IVX9 port map( A => n297, Z => n2647);
   U1951 : HS65_LH_HA1X4 port map( A0 => n2566, B0 => n2563, CO => n1005, S0 =>
                           n1038);
   U1952 : HS65_LH_BFX9 port map( A => b(27), Z => n2618);
   U1953 : HS65_LH_BFX9 port map( A => b(3), Z => n2570);
   U1954 : HS65_LH_BFX9 port map( A => b(2), Z => n2568);
   U1955 : HS65_LH_BFX9 port map( A => b(20), Z => n2604);
   U1956 : HS65_LH_BFX9 port map( A => b(11), Z => n2586);
   U1957 : HS65_LH_BFX9 port map( A => b(4), Z => n2572);
   U1958 : HS65_LH_BFX9 port map( A => b(28), Z => n2620);
   U1959 : HS65_LH_BFX9 port map( A => n2655, Z => n2418);
   U1960 : HS65_LH_BFX9 port map( A => n2655, Z => n2417);
   U1961 : HS65_LH_BFX9 port map( A => n2656, Z => n2421);
   U1962 : HS65_LH_BFX9 port map( A => n2656, Z => n2420);
   U1963 : HS65_LH_BFX9 port map( A => b(31), Z => n2626);
   U1964 : HS65_LH_BFX9 port map( A => n2655, Z => n2419);
   U1965 : HS65_LH_BFX9 port map( A => n2656, Z => n2422);
   U1966 : HS65_LH_BFX9 port map( A => n2562, Z => n2563);
   U1967 : HS65_LH_BFX9 port map( A => n2562, Z => n2564);
   U1968 : HS65_LH_BFX9 port map( A => b(27), Z => n2619);
   U1969 : HS65_LH_BFX9 port map( A => b(2), Z => n2569);
   U1970 : HS65_LH_BFX9 port map( A => b(3), Z => n2571);
   U1971 : HS65_LH_BFX9 port map( A => n2445, Z => n2446);
   U1972 : HS65_LH_BFX9 port map( A => n2458, Z => n2459);
   U1973 : HS65_LH_BFX9 port map( A => n2484, Z => n2485);
   U1974 : HS65_LH_BFX9 port map( A => n2497, Z => n2498);
   U1975 : HS65_LH_BFX9 port map( A => n2510, Z => n2511);
   U1976 : HS65_LH_BFX9 port map( A => n2536, Z => n2537);
   U1977 : HS65_LH_BFX9 port map( A => n2549, Z => n2550);
   U1978 : HS65_LH_BFX9 port map( A => b(20), Z => n2605);
   U1979 : HS65_LH_BFX9 port map( A => b(11), Z => n2587);
   U1980 : HS65_LH_BFX9 port map( A => b(4), Z => n2573);
   U1981 : HS65_LH_BFX9 port map( A => b(28), Z => n2621);
   U1982 : HS65_LH_BFX9 port map( A => n2471, Z => n2472);
   U1983 : HS65_LH_BFX9 port map( A => n2523, Z => n2524);
   U1984 : HS65_LH_BFX9 port map( A => n2433, Z => n2430);
   U1985 : HS65_LH_BFX9 port map( A => n2433, Z => n2431);
   U1986 : HS65_LH_BFX9 port map( A => b(31), Z => n2627);
   U1987 : HS65_LH_BFX9 port map( A => n2523, Z => n2525);
   U1988 : HS65_LH_BFX9 port map( A => n2471, Z => n2473);
   U1989 : HS65_LH_BFX9 port map( A => n2535, Z => n2533);
   U1990 : HS65_LH_BFX9 port map( A => n2531, Z => n2529);
   U1991 : HS65_LH_BFX9 port map( A => n2453, Z => n2451);
   U1992 : HS65_LH_BFX9 port map( A => n2466, Z => n2464);
   U1993 : HS65_LH_BFX9 port map( A => n2479, Z => n2477);
   U1994 : HS65_LH_BFX9 port map( A => n2492, Z => n2490);
   U1995 : HS65_LH_BFX9 port map( A => n2505, Z => n2503);
   U1996 : HS65_LH_BFX9 port map( A => n2518, Z => n2516);
   U1997 : HS65_LH_BFX9 port map( A => n2544, Z => n2542);
   U1998 : HS65_LH_BFX9 port map( A => n2557, Z => n2555);
   U1999 : HS65_LH_BFX9 port map( A => n2445, Z => n2447);
   U2000 : HS65_LH_BFX9 port map( A => n2458, Z => n2460);
   U2001 : HS65_LH_BFX9 port map( A => n2484, Z => n2486);
   U2002 : HS65_LH_BFX9 port map( A => n2497, Z => n2499);
   U2003 : HS65_LH_BFX9 port map( A => n2510, Z => n2512);
   U2004 : HS65_LH_BFX9 port map( A => n2536, Z => n2538);
   U2005 : HS65_LH_BFX9 port map( A => n2549, Z => n2551);
   U2006 : HS65_LH_BFX9 port map( A => n2457, Z => n2454);
   U2007 : HS65_LH_BFX9 port map( A => n2561, Z => n2558);
   U2008 : HS65_LH_BFX9 port map( A => n2470, Z => n2467);
   U2009 : HS65_LH_BFX9 port map( A => n2496, Z => n2493);
   U2010 : HS65_LH_BFX9 port map( A => n2509, Z => n2506);
   U2011 : HS65_LH_BFX9 port map( A => n2522, Z => n2519);
   U2012 : HS65_LH_BFX9 port map( A => n2548, Z => n2545);
   U2013 : HS65_LH_BFX9 port map( A => n2457, Z => n2455);
   U2014 : HS65_LH_BFX9 port map( A => n2470, Z => n2468);
   U2015 : HS65_LH_BFX9 port map( A => n2496, Z => n2494);
   U2016 : HS65_LH_BFX9 port map( A => n2509, Z => n2507);
   U2017 : HS65_LH_BFX9 port map( A => n2522, Z => n2520);
   U2018 : HS65_LH_BFX9 port map( A => n2548, Z => n2546);
   U2019 : HS65_LH_BFX9 port map( A => n2561, Z => n2559);
   U2020 : HS65_LH_BFX9 port map( A => n2483, Z => n2480);
   U2021 : HS65_LH_BFX9 port map( A => n2535, Z => n2532);
   U2022 : HS65_LH_BFX9 port map( A => n2479, Z => n2476);
   U2023 : HS65_LH_BFX9 port map( A => n2531, Z => n2528);
   U2024 : HS65_LH_BFX9 port map( A => n2453, Z => n2450);
   U2025 : HS65_LH_BFX9 port map( A => n2466, Z => n2463);
   U2026 : HS65_LH_BFX9 port map( A => n2492, Z => n2489);
   U2027 : HS65_LH_BFX9 port map( A => n2505, Z => n2502);
   U2028 : HS65_LH_BFX9 port map( A => n2518, Z => n2515);
   U2029 : HS65_LH_BFX9 port map( A => n2544, Z => n2541);
   U2030 : HS65_LH_BFX9 port map( A => n2557, Z => n2554);
   U2031 : HS65_LH_BFX9 port map( A => n2483, Z => n2481);
   U2032 : HS65_LH_IVX9 port map( A => n2632, Z => n2631);
   U2033 : HS65_LH_IVX9 port map( A => n2636, Z => n2635);
   U2034 : HS65_LH_IVX9 port map( A => a(8), Z => n2632);
   U2035 : HS65_LH_IVX9 port map( A => a(14), Z => n2636);
   U2036 : HS65_LH_BFX9 port map( A => n2562, Z => n2565);
   U2037 : HS65_LH_IVX9 port map( A => n2640, Z => n2639);
   U2038 : HS65_LH_IVX9 port map( A => a(20), Z => n2640);
   U2039 : HS65_LH_IVX9 port map( A => n2634, Z => n2633);
   U2040 : HS65_LH_IVX9 port map( A => a(11), Z => n2634);
   U2041 : HS65_LH_IVX9 port map( A => n2644, Z => n2643);
   U2042 : HS65_LH_IVX9 port map( A => a(26), Z => n2644);
   U2043 : HS65_LH_IVX9 port map( A => n2630, Z => n2629);
   U2044 : HS65_LH_IVX9 port map( A => n2638, Z => n2637);
   U2045 : HS65_LH_IVX9 port map( A => a(5), Z => n2630);
   U2046 : HS65_LH_IVX9 port map( A => a(17), Z => n2638);
   U2047 : HS65_LH_IVX9 port map( A => n2646, Z => n2645);
   U2048 : HS65_LH_IVX9 port map( A => a(29), Z => n2646);
   U2049 : HS65_LH_BFX9 port map( A => n2433, Z => n2432);
   U2050 : HS65_LH_BFX9 port map( A => n2457, Z => n2456);
   U2051 : HS65_LH_BFX9 port map( A => n2470, Z => n2469);
   U2052 : HS65_LH_BFX9 port map( A => n2496, Z => n2495);
   U2053 : HS65_LH_BFX9 port map( A => n2509, Z => n2508);
   U2054 : HS65_LH_BFX9 port map( A => n2522, Z => n2521);
   U2055 : HS65_LH_BFX9 port map( A => n2548, Z => n2547);
   U2056 : HS65_LH_BFX9 port map( A => n2561, Z => n2560);
   U2057 : HS65_LH_BFX9 port map( A => n2483, Z => n2482);
   U2058 : HS65_LH_BFX9 port map( A => n2535, Z => n2534);
   U2059 : HS65_LH_BFX9 port map( A => n2531, Z => n2530);
   U2060 : HS65_LH_BFX9 port map( A => n2453, Z => n2452);
   U2061 : HS65_LH_BFX9 port map( A => n2466, Z => n2465);
   U2062 : HS65_LH_BFX9 port map( A => n2479, Z => n2478);
   U2063 : HS65_LH_BFX9 port map( A => n2492, Z => n2491);
   U2064 : HS65_LH_BFX9 port map( A => n2505, Z => n2504);
   U2065 : HS65_LH_BFX9 port map( A => n2518, Z => n2517);
   U2066 : HS65_LH_BFX9 port map( A => n2544, Z => n2543);
   U2067 : HS65_LH_BFX9 port map( A => n2557, Z => n2556);
   U2068 : HS65_LH_IVX9 port map( A => n2642, Z => n2641);
   U2069 : HS65_LH_IVX9 port map( A => a(23), Z => n2642);
   U2070 : HS65_LH_IVX9 port map( A => n2449, Z => n2448);
   U2071 : HS65_LH_IVX9 port map( A => n2462, Z => n2461);
   U2072 : HS65_LH_IVX9 port map( A => n2475, Z => n2474);
   U2073 : HS65_LH_IVX9 port map( A => n2488, Z => n2487);
   U2074 : HS65_LH_IVX9 port map( A => n2501, Z => n2500);
   U2075 : HS65_LH_IVX9 port map( A => n2514, Z => n2513);
   U2076 : HS65_LH_IVX9 port map( A => n2527, Z => n2526);
   U2077 : HS65_LH_IVX9 port map( A => n2540, Z => n2539);
   U2078 : HS65_LH_IVX9 port map( A => n2553, Z => n2552);
   U2079 : HS65_LH_IVX9 port map( A => n2662, Z => n2655);
   U2080 : HS65_LH_IVX9 port map( A => n2702, Z => n2656);
   U2081 : HS65_LH_BFX9 port map( A => n2712, Z => n2457);
   U2082 : HS65_LH_BFX9 port map( A => n3056, Z => n2561);
   U2083 : HS65_LH_BFX9 port map( A => n2755, Z => n2470);
   U2084 : HS65_LH_BFX9 port map( A => n2798, Z => n2483);
   U2085 : HS65_LH_BFX9 port map( A => n2841, Z => n2496);
   U2086 : HS65_LH_BFX9 port map( A => n2884, Z => n2509);
   U2087 : HS65_LH_BFX9 port map( A => n2927, Z => n2522);
   U2088 : HS65_LH_BFX9 port map( A => n2970, Z => n2535);
   U2089 : HS65_LH_BFX9 port map( A => n3013, Z => n2548);
   U2090 : HS65_LH_BFX9 port map( A => n2710, Z => n2453);
   U2091 : HS65_LH_BFX9 port map( A => n2753, Z => n2466);
   U2092 : HS65_LH_BFX9 port map( A => n2839, Z => n2492);
   U2093 : HS65_LH_BFX9 port map( A => n2882, Z => n2505);
   U2094 : HS65_LH_BFX9 port map( A => n2925, Z => n2518);
   U2095 : HS65_LH_BFX9 port map( A => n2968, Z => n2531);
   U2096 : HS65_LH_BFX9 port map( A => n3011, Z => n2544);
   U2097 : HS65_LH_BFX9 port map( A => n3054, Z => n2557);
   U2098 : HS65_LH_BFX9 port map( A => n2796, Z => n2479);
   U2099 : HS65_LH_BFX9 port map( A => n2661, Z => n2433);
   U2100 : HS65_LH_IVX9 port map( A => n2708, Z => n2449);
   U2101 : HS65_LH_IVX9 port map( A => n2751, Z => n2462);
   U2102 : HS65_LH_IVX9 port map( A => n2794, Z => n2475);
   U2103 : HS65_LH_IVX9 port map( A => n2837, Z => n2488);
   U2104 : HS65_LH_IVX9 port map( A => n2880, Z => n2501);
   U2105 : HS65_LH_IVX9 port map( A => n2923, Z => n2514);
   U2106 : HS65_LH_IVX9 port map( A => n2966, Z => n2527);
   U2107 : HS65_LH_IVX9 port map( A => n3009, Z => n2540);
   U2108 : HS65_LH_IVX9 port map( A => n3052, Z => n2553);
   U2109 : HS65_LH_BFX9 port map( A => b(0), Z => n2562);
   U2110 : HS65_LH_BFX9 port map( A => n2707, Z => n2445);
   U2111 : HS65_LH_BFX9 port map( A => n2793, Z => n2471);
   U2112 : HS65_LH_BFX9 port map( A => n2750, Z => n2458);
   U2113 : HS65_LH_BFX9 port map( A => n2836, Z => n2484);
   U2114 : HS65_LH_BFX9 port map( A => n2879, Z => n2497);
   U2115 : HS65_LH_BFX9 port map( A => n2922, Z => n2510);
   U2116 : HS65_LH_BFX9 port map( A => n2965, Z => n2523);
   U2117 : HS65_LH_BFX9 port map( A => n3008, Z => n2536);
   U2118 : HS65_LH_BFX9 port map( A => n3051, Z => n2549);
   U2119 : HS65_LH_BFX9 port map( A => b(1), Z => n2566);
   U2120 : HS65_LH_BFX9 port map( A => b(19), Z => n2602);
   U2121 : HS65_LH_BFX9 port map( A => b(23), Z => n2610);
   U2122 : HS65_LH_BFX9 port map( A => b(25), Z => n2614);
   U2123 : HS65_LH_BFX9 port map( A => b(12), Z => n2588);
   U2124 : HS65_LH_BFX9 port map( A => b(13), Z => n2590);
   U2125 : HS65_LH_BFX9 port map( A => b(24), Z => n2612);
   U2126 : HS65_LH_BFX9 port map( A => b(26), Z => n2616);
   U2127 : HS65_LH_BFX9 port map( A => b(18), Z => n2600);
   U2128 : HS65_LH_BFX9 port map( A => b(5), Z => n2574);
   U2129 : HS65_LH_BFX9 port map( A => b(7), Z => n2578);
   U2130 : HS65_LH_BFX9 port map( A => b(15), Z => n2594);
   U2131 : HS65_LH_BFX9 port map( A => b(9), Z => n2582);
   U2132 : HS65_LH_BFX9 port map( A => b(17), Z => n2598);
   U2133 : HS65_LH_BFX9 port map( A => b(22), Z => n2608);
   U2134 : HS65_LH_BFX9 port map( A => b(21), Z => n2606);
   U2135 : HS65_LH_BFX9 port map( A => b(29), Z => n2622);
   U2136 : HS65_LH_BFX9 port map( A => b(30), Z => n2624);
   U2137 : HS65_LH_BFX9 port map( A => b(16), Z => n2596);
   U2138 : HS65_LH_BFX9 port map( A => b(6), Z => n2576);
   U2139 : HS65_LH_BFX9 port map( A => b(14), Z => n2592);
   U2140 : HS65_LH_BFX9 port map( A => b(8), Z => n2580);
   U2141 : HS65_LH_BFX9 port map( A => b(10), Z => n2584);
   U2142 : HS65_LH_BFX9 port map( A => n2425, Z => n2423);
   U2143 : HS65_LH_BFX9 port map( A => b(19), Z => n2603);
   U2144 : HS65_LH_BFX9 port map( A => n2425, Z => n2424);
   U2145 : HS65_LH_BFX9 port map( A => b(23), Z => n2611);
   U2146 : HS65_LH_BFX9 port map( A => n2436, Z => n2434);
   U2147 : HS65_LH_BFX9 port map( A => n2440, Z => n2437);
   U2148 : HS65_LH_BFX9 port map( A => b(25), Z => n2615);
   U2149 : HS65_LH_BFX9 port map( A => b(12), Z => n2589);
   U2150 : HS65_LH_BFX9 port map( A => b(13), Z => n2591);
   U2151 : HS65_LH_BFX9 port map( A => n2440, Z => n2438);
   U2152 : HS65_LH_BFX9 port map( A => b(24), Z => n2613);
   U2153 : HS65_LH_BFX9 port map( A => b(26), Z => n2617);
   U2154 : HS65_LH_BFX9 port map( A => b(18), Z => n2601);
   U2155 : HS65_LH_BFX9 port map( A => b(5), Z => n2575);
   U2156 : HS65_LH_BFX9 port map( A => b(7), Z => n2579);
   U2157 : HS65_LH_BFX9 port map( A => b(15), Z => n2595);
   U2158 : HS65_LH_BFX9 port map( A => b(9), Z => n2583);
   U2159 : HS65_LH_BFX9 port map( A => b(21), Z => n2607);
   U2160 : HS65_LH_BFX9 port map( A => b(17), Z => n2599);
   U2161 : HS65_LH_BFX9 port map( A => b(22), Z => n2609);
   U2162 : HS65_LH_BFX9 port map( A => b(29), Z => n2623);
   U2163 : HS65_LH_BFX9 port map( A => n2436, Z => n2435);
   U2164 : HS65_LH_BFX9 port map( A => b(1), Z => n2567);
   U2165 : HS65_LH_BFX9 port map( A => b(30), Z => n2625);
   U2166 : HS65_LH_BFX9 port map( A => b(14), Z => n2593);
   U2167 : HS65_LH_BFX9 port map( A => b(6), Z => n2577);
   U2168 : HS65_LH_BFX9 port map( A => b(8), Z => n2581);
   U2169 : HS65_LH_BFX9 port map( A => b(10), Z => n2585);
   U2170 : HS65_LH_BFX9 port map( A => b(16), Z => n2597);
   U2171 : HS65_LH_BFX9 port map( A => n2444, Z => n2441);
   U2172 : HS65_LH_BFX9 port map( A => n2444, Z => n2442);
   U2173 : HS65_LH_BFX9 port map( A => n2429, Z => n2426);
   U2174 : HS65_LH_BFX9 port map( A => n2429, Z => n2427);
   U2175 : HS65_LH_BFX9 port map( A => n2444, Z => n2443);
   U2176 : HS65_LH_BFX9 port map( A => n2429, Z => n2428);
   U2177 : HS65_LH_BFX9 port map( A => n2440, Z => n2439);
   U2178 : HS65_LH_BFX9 port map( A => n2670, Z => n2444);
   U2179 : HS65_LH_BFX9 port map( A => n2659, Z => n2425);
   U2180 : HS65_LH_BFX9 port map( A => n2668, Z => n2440);
   U2181 : HS65_LH_BFX9 port map( A => n2660, Z => n2429);
   U2182 : HS65_LH_BFX9 port map( A => n2666, Z => n2436);
   U2183 : HS65_LHS_XOR3X2 port map( A => n292, B => n227, C => n2658, Z => 
                           product(63));
   U2184 : HS65_LH_AO22X4 port map( A => n2627, B => n2423, C => n2419, D => 
                           n1006, Z => n2658);
   U2185 : HS65_LH_MX41X4 port map( D0 => n1025, S0 => n2419, D1 => n2593, S1 
                           => n2427, D2 => n2591, S2 => n2431, D3 => n2589, S3 
                           => n2423, Z => n419);
   U2186 : HS65_LH_MX41X4 port map( D0 => n1019, S0 => n2419, D1 => n2601, S1 
                           => n2423, D2 => n2603, S2 => n2430, D3 => n2605, S3 
                           => n2426, Z => n352);
   U2187 : HS65_LH_MX41X4 port map( D0 => n1013, S0 => n2419, D1 => n2613, S1 
                           => n2423, D2 => n2615, S2 => n2430, D3 => n2617, S3 
                           => n2426, Z => n309);
   U2188 : HS65_LH_OA12X4 port map( A => n2662, B => n2657, C => n2663, Z => 
                           n292);
   U2189 : HS65_LH_OAI22X1 port map( A => n2625, B => n2664, C => n2423, D => 
                           n2664, Z => n2663);
   U2190 : HS65_LH_AND2X4 port map( A => n2626, B => n2430, Z => n2664);
   U2191 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2665, Z => n1419);
   U2192 : HS65_LH_AO22X4 port map( A => n2565, B => n2434, C => n2422, D => 
                           n2564, Z => n2665);
   U2193 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2667, Z => n1418);
   U2194 : HS65_LH_AO222X4 port map( A => n2564, B => n2437, C => n2434, D => 
                           n2566, E => n2422, F => n1038, Z => n2667);
   U2195 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2669, Z => n1417);
   U2196 : HS65_LH_MX41X4 port map( D0 => n1037, S0 => n2422, D1 => n2442, S1 
                           => n2564, D2 => n2439, S2 => n2566, D3 => n2569, S3 
                           => n2434, Z => n2669);
   U2197 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2671, Z => n1416);
   U2198 : HS65_LH_MX41X4 port map( D0 => n1036, S0 => n2421, D1 => n2443, S1 
                           => n2567, D2 => n2569, S2 => n2437, D3 => n2571, S3 
                           => n2434, Z => n2671);
   U2199 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2672, Z => n1415);
   U2200 : HS65_LH_MX41X4 port map( D0 => n1035, S0 => n2422, D1 => n2443, S1 
                           => n2569, D2 => n2571, S2 => n2437, D3 => n2573, S3 
                           => n2434, Z => n2672);
   U2201 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2673, Z => n1414);
   U2202 : HS65_LH_MX41X4 port map( D0 => n1034, S0 => n2422, D1 => n2571, S1 
                           => n2441, D2 => n2573, S2 => n2437, D3 => n2575, S3 
                           => n2434, Z => n2673);
   U2203 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2674, Z => n1413);
   U2204 : HS65_LH_MX41X4 port map( D0 => n1033, S0 => n2421, D1 => n2573, S1 
                           => n2441, D2 => n2575, S2 => n2437, D3 => n2577, S3 
                           => n2434, Z => n2674);
   U2205 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2675, Z => n1412);
   U2206 : HS65_LH_MX41X4 port map( D0 => n1032, S0 => n2421, D1 => n2575, S1 
                           => n2441, D2 => n2577, S2 => n2437, D3 => n2579, S3 
                           => n2434, Z => n2675);
   U2207 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2676, Z => n1411);
   U2208 : HS65_LH_MX41X4 port map( D0 => n1031, S0 => n2421, D1 => n2577, S1 
                           => n2441, D2 => n2579, S2 => n2437, D3 => n2581, S3 
                           => n2434, Z => n2676);
   U2209 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2677, Z => n1410);
   U2210 : HS65_LH_MX41X4 port map( D0 => n1030, S0 => n2421, D1 => n2579, S1 
                           => n2441, D2 => n2581, S2 => n2437, D3 => n2583, S3 
                           => n2434, Z => n2677);
   U2211 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2678, Z => n1409);
   U2212 : HS65_LH_MX41X4 port map( D0 => n1029, S0 => n2421, D1 => n2581, S1 
                           => n2441, D2 => n2583, S2 => n2437, D3 => n2585, S3 
                           => n2434, Z => n2678);
   U2213 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2679, Z => n1408);
   U2214 : HS65_LH_MX41X4 port map( D0 => n1028, S0 => n2421, D1 => n2583, S1 
                           => n2441, D2 => n2585, S2 => n2437, D3 => n2587, S3 
                           => n2434, Z => n2679);
   U2215 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2680, Z => n1407);
   U2216 : HS65_LH_MX41X4 port map( D0 => n1027, S0 => n2421, D1 => n2585, S1 
                           => n2441, D2 => n2587, S2 => n2437, D3 => n2435, S3 
                           => n2589, Z => n2680);
   U2217 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2681, Z => n1406);
   U2218 : HS65_LH_MX41X4 port map( D0 => n1026, S0 => n2421, D1 => n2587, S1 
                           => n2441, D2 => n2438, S2 => n2588, D3 => n2435, S3 
                           => n2591, Z => n2681);
   U2219 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2682, Z => n1405);
   U2220 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1025, D1 => n2442, S1 
                           => n2589, D2 => n2438, S2 => n2590, D3 => n2435, S3 
                           => n2593, Z => n2682);
   U2221 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2683, Z => n1404);
   U2222 : HS65_LH_MX41X4 port map( D0 => n1024, S0 => n2421, D1 => n2442, S1 
                           => n2591, D2 => n2438, S2 => n2592, D3 => n2595, S3 
                           => n2434, Z => n2683);
   U2223 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2684, Z => n1403);
   U2224 : HS65_LH_MX41X4 port map( D0 => n1023, S0 => n2421, D1 => n2442, S1 
                           => n2593, D2 => n2595, S2 => n2437, D3 => n2597, S3 
                           => n2434, Z => n2684);
   U2225 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2685, Z => n1402);
   U2226 : HS65_LH_MX41X4 port map( D0 => n1022, S0 => n2420, D1 => n2595, S1 
                           => n2441, D2 => n2597, S2 => n2437, D3 => n2599, S3 
                           => n2434, Z => n2685);
   U2227 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2686, Z => n1401);
   U2228 : HS65_LH_MX41X4 port map( D0 => n1021, S0 => n2420, D1 => n2597, S1 
                           => n2441, D2 => n2599, S2 => n2437, D3 => n2435, S3 
                           => n2601, Z => n2686);
   U2229 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2687, Z => n1400);
   U2230 : HS65_LH_MX41X4 port map( D0 => n1020, S0 => n2420, D1 => n2599, S1 
                           => n2441, D2 => n2438, S2 => n2600, D3 => n2435, S3 
                           => n2603, Z => n2687);
   U2231 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2688, Z => n1399);
   U2232 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1019, D1 => n2442, S1 
                           => n2601, D2 => n2438, S2 => n2602, D3 => n2435, S3 
                           => n2605, Z => n2688);
   U2233 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2689, Z => n1398);
   U2234 : HS65_LH_MX41X4 port map( D0 => n1018, S0 => n2420, D1 => n2442, S1 
                           => n2603, D2 => n2438, S2 => n2604, D3 => n2607, S3 
                           => n2435, Z => n2689);
   U2235 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2690, Z => n1397);
   U2236 : HS65_LH_MX41X4 port map( D0 => n1017, S0 => n2420, D1 => n2442, S1 
                           => n2605, D2 => n2607, S2 => n2438, D3 => n2609, S3 
                           => n2434, Z => n2690);
   U2237 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2691, Z => n1396);
   U2238 : HS65_LH_MX41X4 port map( D0 => n1016, S0 => n2420, D1 => n2607, S1 
                           => n2442, D2 => n2609, S2 => n2438, D3 => n2611, S3 
                           => n2435, Z => n2691);
   U2239 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2692, Z => n1395);
   U2240 : HS65_LH_MX41X4 port map( D0 => n1015, S0 => n2421, D1 => n2609, S1 
                           => n2442, D2 => n2611, S2 => n2438, D3 => n2435, S3 
                           => n2613, Z => n2692);
   U2241 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2693, Z => n1394);
   U2242 : HS65_LH_MX41X4 port map( D0 => n1014, S0 => n2420, D1 => n2611, S1 
                           => n2442, D2 => n2439, S2 => n2612, D3 => n2435, S3 
                           => n2615, Z => n2693);
   U2243 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2694, Z => n1393);
   U2244 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1013, D1 => n2443, S1 
                           => n2613, D2 => n2438, S2 => n2614, D3 => n2435, S3 
                           => n2617, Z => n2694);
   U2245 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2695, Z => n1392);
   U2246 : HS65_LH_MX41X4 port map( D0 => n1012, S0 => n2420, D1 => n2443, S1 
                           => n2615, D2 => n2439, S2 => n2616, D3 => n2619, S3 
                           => n2435, Z => n2695);
   U2247 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2696, Z => n1391);
   U2248 : HS65_LH_MX41X4 port map( D0 => n1011, S0 => n2420, D1 => n2443, S1 
                           => n2617, D2 => n2619, S2 => n2438, D3 => n2621, S3 
                           => n2435, Z => n2696);
   U2249 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2697, Z => n1390);
   U2250 : HS65_LH_MX41X4 port map( D0 => n1010, S0 => n2420, D1 => n2619, S1 
                           => n2442, D2 => n2621, S2 => n2438, D3 => n2623, S3 
                           => n2435, Z => n2697);
   U2251 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2698, Z => n1389);
   U2252 : HS65_LH_MX41X4 port map( D0 => n1009, S0 => n2420, D1 => n2621, S1 
                           => n2442, D2 => n2623, S2 => n2438, D3 => n2625, S3 
                           => n2435, Z => n2698);
   U2253 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2699, Z => n1388);
   U2254 : HS65_LH_MX41X4 port map( D0 => n1008, S0 => n2420, D1 => n2623, S1 
                           => n2442, D2 => n2625, S2 => n2438, D3 => n2435, S3 
                           => n2627, Z => n2699);
   U2255 : HS65_LH_NOR2AX3 port map( A => a(0), B => n2700, Z => n2666);
   U2256 : HS65_LHS_XOR2X3 port map( A => a(2), B => n2701, Z => n1387);
   U2257 : HS65_LH_OAI12X2 port map( A => n2657, B => n2702, C => n2703, Z => 
                           n2701);
   U2258 : HS65_LH_OAI22X1 port map( A => n2625, B => n2704, C => n2441, D => 
                           n2704, Z => n2703);
   U2259 : HS65_LH_AND2X4 port map( A => n2438, B => n2626, Z => n2704);
   U2260 : HS65_LH_NOR2AX3 port map( A => a(1), B => a(0), Z => n2668);
   U2261 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2705, Z => n1386);
   U2262 : HS65_LH_AOI22X1 port map( A => n2422, B => n1006, C => n2443, D => 
                           n2627, Z => n2705);
   U2263 : HS65_LH_NOR3AX2 port map( A => n2700, B => a(0), C => a(1), Z => 
                           n2670);
   U2264 : HS65_LH_NAND2X2 port map( A => a(0), B => n2700, Z => n2702);
   U2265 : HS65_LHS_XOR2X3 port map( A => a(2), B => a(1), Z => n2700);
   U2266 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2706, Z => n1384);
   U2267 : HS65_LH_AO22X4 port map( A => n2565, B => n2446, C => n2564, D => 
                           n2708, Z => n2706);
   U2268 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2709, Z => n1383);
   U2269 : HS65_LH_AO222X4 port map( A => n2567, B => n2446, C => n2563, D => 
                           n2450, E => n1038, F => n2708, Z => n2709);
   U2270 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2711, Z => n1382);
   U2271 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1037, D1 => n2455, S1 
                           => n2564, D2 => n2450, S2 => n2566, D3 => n2446, S3 
                           => n2569, Z => n2711);
   U2272 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2713, Z => n1381);
   U2273 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1036, D1 => n2454, S1 
                           => n2567, D2 => n2450, S2 => n2568, D3 => n2446, S3 
                           => n2571, Z => n2713);
   U2274 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2714, Z => n1380);
   U2275 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1035, D1 => n2454, S1 
                           => n2569, D2 => n2450, S2 => n2570, D3 => n2446, S3 
                           => n2573, Z => n2714);
   U2276 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2715, Z => n1379);
   U2277 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1034, D1 => n2454, S1 
                           => n2571, D2 => n2450, S2 => n2572, D3 => n2446, S3 
                           => n2575, Z => n2715);
   U2278 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2716, Z => n1378);
   U2279 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1033, D1 => n2454, S1 
                           => n2573, D2 => n2450, S2 => n2574, D3 => n2446, S3 
                           => n2577, Z => n2716);
   U2280 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2717, Z => n1377);
   U2281 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1032, D1 => n2454, S1 
                           => n2575, D2 => n2450, S2 => n2576, D3 => n2446, S3 
                           => n2579, Z => n2717);
   U2282 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2718, Z => n1376);
   U2283 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1031, D1 => n2454, S1 
                           => n2577, D2 => n2450, S2 => n2578, D3 => n2446, S3 
                           => n2581, Z => n2718);
   U2284 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2719, Z => n1375);
   U2285 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1030, D1 => n2454, S1 
                           => n2579, D2 => n2451, S2 => n2580, D3 => n2446, S3 
                           => n2583, Z => n2719);
   U2286 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2720, Z => n1374);
   U2287 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1029, D1 => n2454, S1 
                           => n2581, D2 => n2450, S2 => n2582, D3 => n2446, S3 
                           => n2585, Z => n2720);
   U2288 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2721, Z => n1373);
   U2289 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1028, D1 => n2454, S1 
                           => n2583, D2 => n2450, S2 => n2584, D3 => n2446, S3 
                           => n2587, Z => n2721);
   U2290 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2722, Z => n1372);
   U2291 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1027, D1 => n2454, S1 
                           => n2585, D2 => n2450, S2 => n2586, D3 => n2446, S3 
                           => n2589, Z => n2722);
   U2292 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2723, Z => n1371);
   U2293 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1026, D1 => n2454, S1 
                           => n2587, D2 => n2451, S2 => n2588, D3 => n2446, S3 
                           => n2591, Z => n2723);
   U2294 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2724, Z => n1370);
   U2295 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1025, D1 => n2454, S1 
                           => n2589, D2 => n2451, S2 => n2590, D3 => n2446, S3 
                           => n2592, Z => n2724);
   U2296 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2725, Z => n1369);
   U2297 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1024, D1 => n2455, S1 
                           => n2591, D2 => n2451, S2 => n2592, D3 => n2446, S3 
                           => n2595, Z => n2725);
   U2298 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2726, Z => n1368);
   U2299 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1023, D1 => n2455, S1 
                           => n2593, D2 => n2451, S2 => n2594, D3 => n2446, S3 
                           => n2597, Z => n2726);
   U2300 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2727, Z => n1367);
   U2301 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1022, D1 => n2455, S1 
                           => n2595, D2 => n2451, S2 => n2596, D3 => n2447, S3 
                           => n2599, Z => n2727);
   U2302 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2728, Z => n1366);
   U2303 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1021, D1 => n2455, S1 
                           => n2597, D2 => n2451, S2 => n2598, D3 => n2447, S3 
                           => n2600, Z => n2728);
   U2304 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2729, Z => n1365);
   U2305 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1020, D1 => n2455, S1 
                           => n2599, D2 => n2451, S2 => n2600, D3 => n2447, S3 
                           => n2602, Z => n2729);
   U2306 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2730, Z => n1364);
   U2307 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1019, D1 => n2455, S1 
                           => n2601, D2 => n2451, S2 => n2602, D3 => n2447, S3 
                           => n2604, Z => n2730);
   U2308 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2731, Z => n1363);
   U2309 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1018, D1 => n2455, S1 
                           => n2603, D2 => n2451, S2 => n2604, D3 => n2447, S3 
                           => n2607, Z => n2731);
   U2310 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2732, Z => n1362);
   U2311 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1017, D1 => n2455, S1 
                           => n2605, D2 => n2451, S2 => n2606, D3 => n2447, S3 
                           => n2609, Z => n2732);
   U2312 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2733, Z => n1361);
   U2313 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1016, D1 => n2455, S1 
                           => n2607, D2 => n2451, S2 => n2608, D3 => n2447, S3 
                           => n2611, Z => n2733);
   U2314 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2734, Z => n1360);
   U2315 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1015, D1 => n2455, S1 
                           => n2609, D2 => n2451, S2 => n2610, D3 => n2447, S3 
                           => n2612, Z => n2734);
   U2316 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2735, Z => n1359);
   U2317 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1014, D1 => n2455, S1 
                           => n2611, D2 => n2451, S2 => n2612, D3 => n2447, S3 
                           => n2614, Z => n2735);
   U2318 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2736, Z => n1358);
   U2319 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1013, D1 => n2455, S1 
                           => n2613, D2 => n2452, S2 => n2614, D3 => n2447, S3 
                           => n2616, Z => n2736);
   U2320 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2737, Z => n1357);
   U2321 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1012, D1 => n2456, S1 
                           => n2615, D2 => n2452, S2 => n2616, D3 => n2447, S3 
                           => n2619, Z => n2737);
   U2322 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2738, Z => n1356);
   U2323 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1011, D1 => n2456, S1 
                           => n2617, D2 => n2452, S2 => n2618, D3 => n2447, S3 
                           => n2621, Z => n2738);
   U2324 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2739, Z => n1355);
   U2325 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1010, D1 => n2456, S1 
                           => n2619, D2 => n2452, S2 => n2620, D3 => n2447, S3 
                           => n2623, Z => n2739);
   U2326 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2740, Z => n1354);
   U2327 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1009, D1 => n2456, S1 
                           => n2621, D2 => n2452, S2 => n2622, D3 => n2447, S3 
                           => n2624, Z => n2740);
   U2328 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2741, Z => n1353);
   U2329 : HS65_LH_MX41X4 port map( D0 => n2708, S0 => n1008, D1 => n2456, S1 
                           => n2623, D2 => n2450, S2 => n2624, D3 => n2447, S3 
                           => n2627, Z => n2741);
   U2330 : HS65_LH_AND2X4 port map( A => n2742, B => n2743, Z => n2707);
   U2331 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2744, Z => n1352);
   U2332 : HS65_LH_OAI12X2 port map( A => n2657, B => n2449, C => n2745, Z => 
                           n2744);
   U2333 : HS65_LH_OAI22X1 port map( A => n2625, B => n2746, C => n2454, D => 
                           n2746, Z => n2745);
   U2334 : HS65_LH_AND2X4 port map( A => n2450, B => n2626, Z => n2746);
   U2335 : HS65_LH_NOR2X2 port map( A => n2742, B => n2747, Z => n2710);
   U2336 : HS65_LHS_XOR2X3 port map( A => n2630, B => n2748, Z => n1351);
   U2337 : HS65_LH_AOI22X1 port map( A => n2708, B => n1006, C => n2456, D => 
                           n2627, Z => n2748);
   U2338 : HS65_LH_NOR3AX2 port map( A => n2747, B => n2743, C => n2742, Z => 
                           n2712);
   U2339 : HS65_LHS_XNOR2X3 port map( A => a(4), B => a(3), Z => n2747);
   U2340 : HS65_LH_NOR2AX3 port map( A => n2742, B => n2743, Z => n2708);
   U2341 : HS65_LHS_XNOR2X3 port map( A => n2629, B => a(4), Z => n2743);
   U2342 : HS65_LHS_XOR2X3 port map( A => a(2), B => a(3), Z => n2742);
   U2343 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2749, Z => n1349);
   U2344 : HS65_LH_AO22X4 port map( A => n2565, B => n2459, C => n2564, D => 
                           n2751, Z => n2749);
   U2345 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2752, Z => n1348);
   U2346 : HS65_LH_AO222X4 port map( A => n2567, B => n2459, C => n2563, D => 
                           n2463, E => n1038, F => n2751, Z => n2752);
   U2347 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2754, Z => n1347);
   U2348 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1037, D1 => n2468, S1 
                           => n2564, D2 => n2463, S2 => n2566, D3 => n2459, S3 
                           => n2569, Z => n2754);
   U2349 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2756, Z => n1346);
   U2350 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1036, D1 => n2467, S1 
                           => n2566, D2 => n2463, S2 => n2568, D3 => n2459, S3 
                           => n2571, Z => n2756);
   U2351 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2757, Z => n1345);
   U2352 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1035, D1 => n2467, S1 
                           => n2569, D2 => n2463, S2 => n2570, D3 => n2459, S3 
                           => n2573, Z => n2757);
   U2353 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2758, Z => n1344);
   U2354 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1034, D1 => n2467, S1 
                           => n2571, D2 => n2463, S2 => n2572, D3 => n2459, S3 
                           => n2575, Z => n2758);
   U2355 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2759, Z => n1343);
   U2356 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1033, D1 => n2467, S1 
                           => n2573, D2 => n2463, S2 => n2574, D3 => n2459, S3 
                           => n2577, Z => n2759);
   U2357 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2760, Z => n1342);
   U2358 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1032, D1 => n2467, S1 
                           => n2575, D2 => n2463, S2 => n2576, D3 => n2459, S3 
                           => n2579, Z => n2760);
   U2359 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2761, Z => n1341);
   U2360 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1031, D1 => n2467, S1 
                           => n2577, D2 => n2463, S2 => n2578, D3 => n2459, S3 
                           => n2581, Z => n2761);
   U2361 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2762, Z => n1340);
   U2362 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1030, D1 => n2467, S1 
                           => n2579, D2 => n2464, S2 => n2580, D3 => n2459, S3 
                           => n2583, Z => n2762);
   U2363 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2763, Z => n1339);
   U2364 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1029, D1 => n2467, S1 
                           => n2581, D2 => n2463, S2 => n2582, D3 => n2459, S3 
                           => n2585, Z => n2763);
   U2365 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2764, Z => n1338);
   U2366 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1028, D1 => n2467, S1 
                           => n2583, D2 => n2463, S2 => n2584, D3 => n2459, S3 
                           => n2587, Z => n2764);
   U2367 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2765, Z => n1337);
   U2368 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1027, D1 => n2467, S1 
                           => n2585, D2 => n2463, S2 => n2586, D3 => n2459, S3 
                           => n2589, Z => n2765);
   U2369 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2766, Z => n1336);
   U2370 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1026, D1 => n2467, S1 
                           => n2587, D2 => n2464, S2 => n2588, D3 => n2459, S3 
                           => n2591, Z => n2766);
   U2371 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2767, Z => n1335);
   U2372 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1025, D1 => n2467, S1 
                           => n2589, D2 => n2464, S2 => n2590, D3 => n2459, S3 
                           => n2593, Z => n2767);
   U2373 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2768, Z => n1334);
   U2374 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1024, D1 => n2468, S1 
                           => n2591, D2 => n2464, S2 => n2592, D3 => n2459, S3 
                           => n2595, Z => n2768);
   U2375 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2769, Z => n1333);
   U2376 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1023, D1 => n2468, S1 
                           => n2593, D2 => n2464, S2 => n2594, D3 => n2459, S3 
                           => n2597, Z => n2769);
   U2377 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2770, Z => n1332);
   U2378 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1022, D1 => n2468, S1 
                           => n2595, D2 => n2464, S2 => n2596, D3 => n2460, S3 
                           => n2599, Z => n2770);
   U2379 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2771, Z => n1331);
   U2380 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1021, D1 => n2468, S1 
                           => n2597, D2 => n2464, S2 => n2598, D3 => n2460, S3 
                           => n2601, Z => n2771);
   U2381 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2772, Z => n1330);
   U2382 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1020, D1 => n2468, S1 
                           => n2599, D2 => n2464, S2 => n2600, D3 => n2460, S3 
                           => n2603, Z => n2772);
   U2383 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2773, Z => n1329);
   U2384 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1019, D1 => n2468, S1 
                           => n2601, D2 => n2464, S2 => n2602, D3 => n2460, S3 
                           => n2605, Z => n2773);
   U2385 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2774, Z => n1328);
   U2386 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1018, D1 => n2468, S1 
                           => n2603, D2 => n2464, S2 => n2604, D3 => n2460, S3 
                           => n2607, Z => n2774);
   U2387 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2775, Z => n1327);
   U2388 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1017, D1 => n2468, S1 
                           => n2605, D2 => n2464, S2 => n2606, D3 => n2460, S3 
                           => n2609, Z => n2775);
   U2389 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2776, Z => n1326);
   U2390 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1016, D1 => n2468, S1 
                           => n2607, D2 => n2464, S2 => n2608, D3 => n2460, S3 
                           => n2611, Z => n2776);
   U2391 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2777, Z => n1325);
   U2392 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1015, D1 => n2468, S1 
                           => n2609, D2 => n2464, S2 => n2610, D3 => n2460, S3 
                           => n2613, Z => n2777);
   U2393 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2778, Z => n1324);
   U2394 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1014, D1 => n2468, S1 
                           => n2611, D2 => n2464, S2 => n2612, D3 => n2460, S3 
                           => n2615, Z => n2778);
   U2395 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2779, Z => n1323);
   U2396 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1013, D1 => n2468, S1 
                           => n2613, D2 => n2465, S2 => n2614, D3 => n2460, S3 
                           => n2617, Z => n2779);
   U2397 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2780, Z => n1322);
   U2398 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1012, D1 => n2469, S1 
                           => n2615, D2 => n2465, S2 => n2616, D3 => n2460, S3 
                           => n2619, Z => n2780);
   U2399 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2781, Z => n1321);
   U2400 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1011, D1 => n2469, S1 
                           => n2617, D2 => n2465, S2 => n2618, D3 => n2460, S3 
                           => n2621, Z => n2781);
   U2401 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2782, Z => n1320);
   U2402 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1010, D1 => n2469, S1 
                           => n2619, D2 => n2465, S2 => n2620, D3 => n2460, S3 
                           => n2623, Z => n2782);
   U2403 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2783, Z => n1319);
   U2404 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1009, D1 => n2469, S1 
                           => n2621, D2 => n2465, S2 => n2622, D3 => n2460, S3 
                           => n2624, Z => n2783);
   U2405 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2784, Z => n1318);
   U2406 : HS65_LH_MX41X4 port map( D0 => n2751, S0 => n1008, D1 => n2469, S1 
                           => n2623, D2 => n2463, S2 => n2624, D3 => n2460, S3 
                           => n2627, Z => n2784);
   U2407 : HS65_LH_AND2X4 port map( A => n2785, B => n2786, Z => n2750);
   U2408 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2787, Z => n1317);
   U2409 : HS65_LH_OAI12X2 port map( A => n2657, B => n2462, C => n2788, Z => 
                           n2787);
   U2410 : HS65_LH_OAI22X1 port map( A => n2625, B => n2789, C => n2467, D => 
                           n2789, Z => n2788);
   U2411 : HS65_LH_AND2X4 port map( A => n2463, B => n2626, Z => n2789);
   U2412 : HS65_LH_NOR2X2 port map( A => n2785, B => n2790, Z => n2753);
   U2413 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2791, Z => n1316);
   U2414 : HS65_LH_AOI22X1 port map( A => n2751, B => n1006, C => n2469, D => 
                           n2627, Z => n2791);
   U2415 : HS65_LH_NOR3AX2 port map( A => n2790, B => n2786, C => n2785, Z => 
                           n2755);
   U2416 : HS65_LHS_XNOR2X3 port map( A => a(7), B => a(6), Z => n2790);
   U2417 : HS65_LH_NOR2AX3 port map( A => n2785, B => n2786, Z => n2751);
   U2418 : HS65_LHS_XNOR2X3 port map( A => n2631, B => a(7), Z => n2786);
   U2419 : HS65_LHS_XOR2X3 port map( A => n2629, B => a(6), Z => n2785);
   U2420 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2792, Z => n1314);
   U2421 : HS65_LH_AO22X4 port map( A => n2565, B => n2472, C => n2564, D => 
                           n2794, Z => n2792);
   U2422 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2795, Z => n1313);
   U2423 : HS65_LH_AO222X4 port map( A => n2567, B => n2472, C => n2563, D => 
                           n2476, E => n1038, F => n2794, Z => n2795);
   U2424 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2797, Z => n1312);
   U2425 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1037, D1 => n2472, S1 
                           => n2569, D2 => n2477, S2 => n2566, D3 => n2481, S3 
                           => n2564, Z => n2797);
   U2426 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2799, Z => n1311);
   U2427 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1036, D1 => n2472, S1 
                           => n2571, D2 => n2476, S2 => n2568, D3 => n2480, S3 
                           => n2566, Z => n2799);
   U2428 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2800, Z => n1310);
   U2429 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1035, D1 => n2472, S1 
                           => n2573, D2 => n2476, S2 => n2570, D3 => n2480, S3 
                           => n2569, Z => n2800);
   U2430 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2801, Z => n1309);
   U2431 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1034, D1 => n2472, S1 
                           => n2575, D2 => n2476, S2 => n2572, D3 => n2480, S3 
                           => n2571, Z => n2801);
   U2432 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2802, Z => n1308);
   U2433 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1033, D1 => n2472, S1 
                           => n2577, D2 => n2476, S2 => n2574, D3 => n2480, S3 
                           => n2573, Z => n2802);
   U2434 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2803, Z => n1307);
   U2435 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1032, D1 => n2472, S1 
                           => n2579, D2 => n2476, S2 => n2576, D3 => n2480, S3 
                           => n2575, Z => n2803);
   U2436 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2804, Z => n1306);
   U2437 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1031, D1 => n2472, S1 
                           => n2581, D2 => n2476, S2 => n2578, D3 => n2480, S3 
                           => n2577, Z => n2804);
   U2438 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2805, Z => n1305);
   U2439 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1030, D1 => n2472, S1 
                           => n2583, D2 => n2477, S2 => n2580, D3 => n2480, S3 
                           => n2579, Z => n2805);
   U2440 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2806, Z => n1304);
   U2441 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1029, D1 => n2472, S1 
                           => n2585, D2 => n2476, S2 => n2582, D3 => n2480, S3 
                           => n2581, Z => n2806);
   U2442 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2807, Z => n1303);
   U2443 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1028, D1 => n2472, S1 
                           => n2587, D2 => n2477, S2 => n2584, D3 => n2480, S3 
                           => n2583, Z => n2807);
   U2444 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2808, Z => n1302);
   U2445 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1027, D1 => n2472, S1 
                           => n2589, D2 => n2477, S2 => n2586, D3 => n2480, S3 
                           => n2585, Z => n2808);
   U2446 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2809, Z => n1301);
   U2447 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1026, D1 => n2472, S1 
                           => n2591, D2 => n2477, S2 => n2588, D3 => n2480, S3 
                           => n2587, Z => n2809);
   U2448 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2810, Z => n1300);
   U2449 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1025, D1 => n2472, S1 
                           => n2593, D2 => n2477, S2 => n2590, D3 => n2480, S3 
                           => n2589, Z => n2810);
   U2450 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2811, Z => n1299);
   U2451 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1024, D1 => n2476, S1 
                           => n2593, D2 => n2473, S2 => n2594, D3 => n2481, S3 
                           => n2591, Z => n2811);
   U2452 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2812, Z => n1298);
   U2453 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1023, D1 => n2476, S1 
                           => n2595, D2 => n2473, S2 => n2596, D3 => n2481, S3 
                           => n2593, Z => n2812);
   U2454 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2813, Z => n1297);
   U2455 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1022, D1 => n2473, S1 
                           => n2599, D2 => n2477, S2 => n2596, D3 => n2481, S3 
                           => n2595, Z => n2813);
   U2456 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2814, Z => n1296);
   U2457 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1021, D1 => n2473, S1 
                           => n2601, D2 => n2477, S2 => n2598, D3 => n2481, S3 
                           => n2597, Z => n2814);
   U2458 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2815, Z => n1295);
   U2459 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1020, D1 => n2472, S1 
                           => n2603, D2 => n2477, S2 => n2600, D3 => n2481, S3 
                           => n2599, Z => n2815);
   U2460 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2816, Z => n1294);
   U2461 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1019, D1 => n2473, S1 
                           => n2605, D2 => n2477, S2 => n2602, D3 => n2481, S3 
                           => n2601, Z => n2816);
   U2462 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2817, Z => n1293);
   U2463 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1018, D1 => n2473, S1 
                           => n2607, D2 => n2477, S2 => n2604, D3 => n2481, S3 
                           => n2603, Z => n2817);
   U2464 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2818, Z => n1292);
   U2465 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1017, D1 => n2473, S1 
                           => n2609, D2 => n2477, S2 => n2606, D3 => n2481, S3 
                           => n2605, Z => n2818);
   U2466 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2819, Z => n1291);
   U2467 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1016, D1 => n2473, S1 
                           => n2611, D2 => n2477, S2 => n2608, D3 => n2481, S3 
                           => n2607, Z => n2819);
   U2468 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2820, Z => n1290);
   U2469 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1015, D1 => n2473, S1 
                           => n2613, D2 => n2477, S2 => n2610, D3 => n2481, S3 
                           => n2609, Z => n2820);
   U2470 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2821, Z => n1289);
   U2471 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1014, D1 => n2473, S1 
                           => n2615, D2 => n2478, S2 => n2612, D3 => n2481, S3 
                           => n2611, Z => n2821);
   U2472 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2822, Z => n1288);
   U2473 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1013, D1 => n2473, S1 
                           => n2617, D2 => n2478, S2 => n2614, D3 => n2481, S3 
                           => n2613, Z => n2822);
   U2474 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2823, Z => n1287);
   U2475 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1012, D1 => n2473, S1 
                           => n2619, D2 => n2478, S2 => n2616, D3 => n2482, S3 
                           => n2615, Z => n2823);
   U2476 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2824, Z => n1286);
   U2477 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1011, D1 => n2473, S1 
                           => n2621, D2 => n2478, S2 => n2618, D3 => n2482, S3 
                           => n2617, Z => n2824);
   U2478 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2825, Z => n1285);
   U2479 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1010, D1 => n2473, S1 
                           => n2623, D2 => n2478, S2 => n2620, D3 => n2482, S3 
                           => n2619, Z => n2825);
   U2480 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2826, Z => n1284);
   U2481 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1009, D1 => n2473, S1 
                           => n2624, D2 => n2476, S2 => n2622, D3 => n2482, S3 
                           => n2621, Z => n2826);
   U2482 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2827, Z => n1283);
   U2483 : HS65_LH_MX41X4 port map( D0 => n2794, S0 => n1008, D1 => n2476, S1 
                           => n2624, D2 => n2473, S2 => n2626, D3 => n2482, S3 
                           => n2623, Z => n2827);
   U2484 : HS65_LH_AND2X4 port map( A => n2828, B => n2829, Z => n2793);
   U2485 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2830, Z => n1282);
   U2486 : HS65_LH_OAI12X2 port map( A => n2657, B => n2475, C => n2831, Z => 
                           n2830);
   U2487 : HS65_LH_OAI22X1 port map( A => n2625, B => n2832, C => n2480, D => 
                           n2832, Z => n2831);
   U2488 : HS65_LH_AND2X4 port map( A => n2476, B => n2626, Z => n2832);
   U2489 : HS65_LH_NOR2X2 port map( A => n2828, B => n2833, Z => n2796);
   U2490 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2834, Z => n1281);
   U2491 : HS65_LH_AOI22X1 port map( A => n2794, B => n1006, C => n2482, D => 
                           n2627, Z => n2834);
   U2492 : HS65_LH_NOR3AX2 port map( A => n2833, B => n2829, C => n2828, Z => 
                           n2798);
   U2493 : HS65_LHS_XNOR2X3 port map( A => a(9), B => a(10), Z => n2833);
   U2494 : HS65_LH_NOR2AX3 port map( A => n2828, B => n2829, Z => n2794);
   U2495 : HS65_LHS_XNOR2X3 port map( A => n2633, B => a(10), Z => n2829);
   U2496 : HS65_LHS_XOR2X3 port map( A => n2631, B => a(9), Z => n2828);
   U2497 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2835, Z => n1279);
   U2498 : HS65_LH_AO22X4 port map( A => n2565, B => n2485, C => n2564, D => 
                           n2837, Z => n2835);
   U2499 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2838, Z => n1278);
   U2500 : HS65_LH_AO222X4 port map( A => n2567, B => n2485, C => n2563, D => 
                           n2489, E => n1038, F => n2837, Z => n2838);
   U2501 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2840, Z => n1277);
   U2502 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1037, D1 => n2494, S1 
                           => n2563, D2 => n2489, S2 => n2566, D3 => n2485, S3 
                           => n2569, Z => n2840);
   U2503 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2842, Z => n1276);
   U2504 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1036, D1 => n2493, S1 
                           => n2566, D2 => n2489, S2 => n2568, D3 => n2485, S3 
                           => n2571, Z => n2842);
   U2505 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2843, Z => n1275);
   U2506 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1035, D1 => n2493, S1 
                           => n2569, D2 => n2489, S2 => n2570, D3 => n2485, S3 
                           => n2573, Z => n2843);
   U2507 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2844, Z => n1274);
   U2508 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1034, D1 => n2493, S1 
                           => n2571, D2 => n2489, S2 => n2572, D3 => n2485, S3 
                           => n2575, Z => n2844);
   U2509 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2845, Z => n1273);
   U2510 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1033, D1 => n2493, S1 
                           => n2573, D2 => n2489, S2 => n2574, D3 => n2485, S3 
                           => n2577, Z => n2845);
   U2511 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2846, Z => n1272);
   U2512 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1032, D1 => n2493, S1 
                           => n2575, D2 => n2489, S2 => n2576, D3 => n2485, S3 
                           => n2579, Z => n2846);
   U2513 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2847, Z => n1271);
   U2514 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1031, D1 => n2493, S1 
                           => n2577, D2 => n2489, S2 => n2578, D3 => n2485, S3 
                           => n2581, Z => n2847);
   U2515 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2848, Z => n1270);
   U2516 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1030, D1 => n2493, S1 
                           => n2579, D2 => n2490, S2 => n2580, D3 => n2485, S3 
                           => n2583, Z => n2848);
   U2517 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2849, Z => n1269);
   U2518 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1029, D1 => n2493, S1 
                           => n2581, D2 => n2489, S2 => n2582, D3 => n2485, S3 
                           => n2585, Z => n2849);
   U2519 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2850, Z => n1268);
   U2520 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1028, D1 => n2493, S1 
                           => n2583, D2 => n2489, S2 => n2584, D3 => n2485, S3 
                           => n2587, Z => n2850);
   U2521 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2851, Z => n1267);
   U2522 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1027, D1 => n2493, S1 
                           => n2585, D2 => n2489, S2 => n2586, D3 => n2485, S3 
                           => n2589, Z => n2851);
   U2523 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2852, Z => n1266);
   U2524 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1026, D1 => n2493, S1 
                           => n2587, D2 => n2490, S2 => n2588, D3 => n2485, S3 
                           => n2591, Z => n2852);
   U2525 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2853, Z => n1265);
   U2526 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1025, D1 => n2493, S1 
                           => n2589, D2 => n2490, S2 => n2590, D3 => n2485, S3 
                           => n2593, Z => n2853);
   U2527 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2854, Z => n1264);
   U2528 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1024, D1 => n2494, S1 
                           => n2591, D2 => n2490, S2 => n2592, D3 => n2485, S3 
                           => n2595, Z => n2854);
   U2529 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2855, Z => n1263);
   U2530 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1023, D1 => n2494, S1 
                           => n2593, D2 => n2490, S2 => n2594, D3 => n2485, S3 
                           => n2597, Z => n2855);
   U2531 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2856, Z => n1262);
   U2532 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1022, D1 => n2494, S1 
                           => n2595, D2 => n2490, S2 => n2596, D3 => n2486, S3 
                           => n2599, Z => n2856);
   U2533 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2857, Z => n1261);
   U2534 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1021, D1 => n2494, S1 
                           => n2597, D2 => n2490, S2 => n2598, D3 => n2486, S3 
                           => n2601, Z => n2857);
   U2535 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2858, Z => n1260);
   U2536 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1020, D1 => n2494, S1 
                           => n2599, D2 => n2490, S2 => n2600, D3 => n2486, S3 
                           => n2603, Z => n2858);
   U2537 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2859, Z => n1259);
   U2538 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1019, D1 => n2494, S1 
                           => n2601, D2 => n2490, S2 => n2602, D3 => n2486, S3 
                           => n2605, Z => n2859);
   U2539 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2860, Z => n1258);
   U2540 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1018, D1 => n2494, S1 
                           => n2603, D2 => n2490, S2 => n2604, D3 => n2486, S3 
                           => n2607, Z => n2860);
   U2541 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2861, Z => n1257);
   U2542 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1017, D1 => n2494, S1 
                           => n2605, D2 => n2490, S2 => n2606, D3 => n2486, S3 
                           => n2609, Z => n2861);
   U2543 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2862, Z => n1256);
   U2544 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1016, D1 => n2494, S1 
                           => n2607, D2 => n2490, S2 => n2608, D3 => n2486, S3 
                           => n2611, Z => n2862);
   U2545 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2863, Z => n1255);
   U2546 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1015, D1 => n2494, S1 
                           => n2609, D2 => n2490, S2 => n2610, D3 => n2486, S3 
                           => n2613, Z => n2863);
   U2547 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2864, Z => n1254);
   U2548 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1014, D1 => n2494, S1 
                           => n2611, D2 => n2490, S2 => n2612, D3 => n2486, S3 
                           => n2615, Z => n2864);
   U2549 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2865, Z => n1253);
   U2550 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1013, D1 => n2494, S1 
                           => n2613, D2 => n2491, S2 => n2614, D3 => n2486, S3 
                           => n2617, Z => n2865);
   U2551 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2866, Z => n1252);
   U2552 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1012, D1 => n2495, S1 
                           => n2615, D2 => n2491, S2 => n2616, D3 => n2486, S3 
                           => n2619, Z => n2866);
   U2553 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2867, Z => n1251);
   U2554 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1011, D1 => n2495, S1 
                           => n2617, D2 => n2491, S2 => n2618, D3 => n2486, S3 
                           => n2621, Z => n2867);
   U2555 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2868, Z => n1250);
   U2556 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1010, D1 => n2495, S1 
                           => n2619, D2 => n2491, S2 => n2620, D3 => n2486, S3 
                           => n2623, Z => n2868);
   U2557 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2869, Z => n1249);
   U2558 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1009, D1 => n2495, S1 
                           => n2621, D2 => n2491, S2 => n2622, D3 => n2486, S3 
                           => n2624, Z => n2869);
   U2559 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2870, Z => n1248);
   U2560 : HS65_LH_MX41X4 port map( D0 => n2837, S0 => n1008, D1 => n2495, S1 
                           => n2623, D2 => n2489, S2 => n2624, D3 => n2486, S3 
                           => n2627, Z => n2870);
   U2561 : HS65_LH_AND2X4 port map( A => n2871, B => n2872, Z => n2836);
   U2562 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2873, Z => n1247);
   U2563 : HS65_LH_OAI12X2 port map( A => n2657, B => n2488, C => n2874, Z => 
                           n2873);
   U2564 : HS65_LH_OAI22X1 port map( A => n2625, B => n2875, C => n2493, D => 
                           n2875, Z => n2874);
   U2565 : HS65_LH_AND2X4 port map( A => n2489, B => n2626, Z => n2875);
   U2566 : HS65_LH_NOR2X2 port map( A => n2871, B => n2876, Z => n2839);
   U2567 : HS65_LHS_XOR2X3 port map( A => n2636, B => n2877, Z => n1246);
   U2568 : HS65_LH_AOI22X1 port map( A => n2837, B => n1006, C => n2495, D => 
                           n2627, Z => n2877);
   U2569 : HS65_LH_NOR3AX2 port map( A => n2876, B => n2872, C => n2871, Z => 
                           n2841);
   U2570 : HS65_LHS_XNOR2X3 port map( A => a(13), B => a(12), Z => n2876);
   U2571 : HS65_LH_NOR2AX3 port map( A => n2871, B => n2872, Z => n2837);
   U2572 : HS65_LHS_XNOR2X3 port map( A => n2635, B => a(13), Z => n2872);
   U2573 : HS65_LHS_XOR2X3 port map( A => n2633, B => a(12), Z => n2871);
   U2574 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2878, Z => n1244);
   U2575 : HS65_LH_AO22X4 port map( A => n2564, B => n2498, C => n2564, D => 
                           n2880, Z => n2878);
   U2576 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2881, Z => n1243);
   U2577 : HS65_LH_AO222X4 port map( A => n2567, B => n2498, C => n2563, D => 
                           n2502, E => n1038, F => n2880, Z => n2881);
   U2578 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2883, Z => n1242);
   U2579 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1037, D1 => n2507, S1 
                           => n2563, D2 => n2502, S2 => n2566, D3 => n2498, S3 
                           => n2569, Z => n2883);
   U2580 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2885, Z => n1241);
   U2581 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1036, D1 => n2506, S1 
                           => n2566, D2 => n2502, S2 => n2568, D3 => n2498, S3 
                           => n2571, Z => n2885);
   U2582 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2886, Z => n1240);
   U2583 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1035, D1 => n2506, S1 
                           => n2568, D2 => n2502, S2 => n2570, D3 => n2498, S3 
                           => n2573, Z => n2886);
   U2584 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2887, Z => n1239);
   U2585 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1034, D1 => n2506, S1 
                           => n2570, D2 => n2502, S2 => n2572, D3 => n2498, S3 
                           => n2575, Z => n2887);
   U2586 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2888, Z => n1238);
   U2587 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1033, D1 => n2506, S1 
                           => n2572, D2 => n2502, S2 => n2574, D3 => n2498, S3 
                           => n2577, Z => n2888);
   U2588 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2889, Z => n1237);
   U2589 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1032, D1 => n2506, S1 
                           => n2574, D2 => n2502, S2 => n2576, D3 => n2498, S3 
                           => n2579, Z => n2889);
   U2590 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2890, Z => n1236);
   U2591 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1031, D1 => n2506, S1 
                           => n2576, D2 => n2502, S2 => n2578, D3 => n2498, S3 
                           => n2581, Z => n2890);
   U2592 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2891, Z => n1235);
   U2593 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1030, D1 => n2506, S1 
                           => n2578, D2 => n2503, S2 => n2580, D3 => n2498, S3 
                           => n2583, Z => n2891);
   U2594 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2892, Z => n1234);
   U2595 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1029, D1 => n2506, S1 
                           => n2580, D2 => n2502, S2 => n2582, D3 => n2498, S3 
                           => n2585, Z => n2892);
   U2596 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2893, Z => n1233);
   U2597 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1028, D1 => n2506, S1 
                           => n2582, D2 => n2502, S2 => n2584, D3 => n2498, S3 
                           => n2587, Z => n2893);
   U2598 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2894, Z => n1232);
   U2599 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1027, D1 => n2506, S1 
                           => n2584, D2 => n2502, S2 => n2586, D3 => n2498, S3 
                           => n2589, Z => n2894);
   U2600 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2895, Z => n1231);
   U2601 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1026, D1 => n2506, S1 
                           => n2586, D2 => n2503, S2 => n2588, D3 => n2498, S3 
                           => n2591, Z => n2895);
   U2602 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2896, Z => n1230);
   U2603 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1025, D1 => n2506, S1 
                           => n2589, D2 => n2503, S2 => n2590, D3 => n2498, S3 
                           => n2593, Z => n2896);
   U2604 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2897, Z => n1229);
   U2605 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1024, D1 => n2507, S1 
                           => n2591, D2 => n2503, S2 => n2592, D3 => n2498, S3 
                           => n2595, Z => n2897);
   U2606 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2898, Z => n1228);
   U2607 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1023, D1 => n2507, S1 
                           => n2593, D2 => n2503, S2 => n2594, D3 => n2498, S3 
                           => n2597, Z => n2898);
   U2608 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2899, Z => n1227);
   U2609 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1022, D1 => n2507, S1 
                           => n2594, D2 => n2503, S2 => n2596, D3 => n2499, S3 
                           => n2599, Z => n2899);
   U2610 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2900, Z => n1226);
   U2611 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1021, D1 => n2507, S1 
                           => n2597, D2 => n2503, S2 => n2598, D3 => n2499, S3 
                           => n2601, Z => n2900);
   U2612 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2901, Z => n1225);
   U2613 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1020, D1 => n2507, S1 
                           => n2598, D2 => n2503, S2 => n2600, D3 => n2499, S3 
                           => n2603, Z => n2901);
   U2614 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2902, Z => n1224);
   U2615 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1019, D1 => n2507, S1 
                           => n2601, D2 => n2503, S2 => n2602, D3 => n2499, S3 
                           => n2605, Z => n2902);
   U2616 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2903, Z => n1223);
   U2617 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1018, D1 => n2507, S1 
                           => n2603, D2 => n2503, S2 => n2604, D3 => n2499, S3 
                           => n2607, Z => n2903);
   U2618 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2904, Z => n1222);
   U2619 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1017, D1 => n2507, S1 
                           => n2605, D2 => n2503, S2 => n2606, D3 => n2499, S3 
                           => n2609, Z => n2904);
   U2620 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2905, Z => n1221);
   U2621 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1016, D1 => n2507, S1 
                           => n2606, D2 => n2503, S2 => n2608, D3 => n2499, S3 
                           => n2611, Z => n2905);
   U2622 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2906, Z => n1220);
   U2623 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1015, D1 => n2507, S1 
                           => n2608, D2 => n2503, S2 => n2610, D3 => n2499, S3 
                           => n2613, Z => n2906);
   U2624 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2907, Z => n1219);
   U2625 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1014, D1 => n2507, S1 
                           => n2610, D2 => n2503, S2 => n2612, D3 => n2499, S3 
                           => n2615, Z => n2907);
   U2626 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2908, Z => n1218);
   U2627 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1013, D1 => n2507, S1 
                           => n2613, D2 => n2504, S2 => n2614, D3 => n2499, S3 
                           => n2617, Z => n2908);
   U2628 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2909, Z => n1217);
   U2629 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1012, D1 => n2508, S1 
                           => n2615, D2 => n2504, S2 => n2616, D3 => n2499, S3 
                           => n2619, Z => n2909);
   U2630 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2910, Z => n1216);
   U2631 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1011, D1 => n2508, S1 
                           => n2617, D2 => n2504, S2 => n2618, D3 => n2499, S3 
                           => n2621, Z => n2910);
   U2632 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2911, Z => n1215);
   U2633 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1010, D1 => n2508, S1 
                           => n2618, D2 => n2504, S2 => n2620, D3 => n2499, S3 
                           => n2623, Z => n2911);
   U2634 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2912, Z => n1214);
   U2635 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1009, D1 => n2508, S1 
                           => n2620, D2 => n2504, S2 => n2622, D3 => n2499, S3 
                           => n2624, Z => n2912);
   U2636 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2913, Z => n1213);
   U2637 : HS65_LH_MX41X4 port map( D0 => n2880, S0 => n1008, D1 => n2508, S1 
                           => n2622, D2 => n2502, S2 => n2624, D3 => n2499, S3 
                           => n2626, Z => n2913);
   U2638 : HS65_LH_AND2X4 port map( A => n2914, B => n2915, Z => n2879);
   U2639 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2916, Z => n1212);
   U2640 : HS65_LH_OAI12X2 port map( A => n2657, B => n2501, C => n2917, Z => 
                           n2916);
   U2641 : HS65_LH_OAI22X1 port map( A => n2625, B => n2918, C => n2506, D => 
                           n2918, Z => n2917);
   U2642 : HS65_LH_AND2X4 port map( A => n2502, B => n2626, Z => n2918);
   U2643 : HS65_LH_NOR2X2 port map( A => n2914, B => n2919, Z => n2882);
   U2644 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2920, Z => n1211);
   U2645 : HS65_LH_AOI22X1 port map( A => n2880, B => n1006, C => n2508, D => 
                           n2627, Z => n2920);
   U2646 : HS65_LH_NOR3AX2 port map( A => n2919, B => n2915, C => n2914, Z => 
                           n2884);
   U2647 : HS65_LHS_XNOR2X3 port map( A => a(16), B => a(15), Z => n2919);
   U2648 : HS65_LH_NOR2AX3 port map( A => n2914, B => n2915, Z => n2880);
   U2649 : HS65_LHS_XNOR2X3 port map( A => n2637, B => a(16), Z => n2915);
   U2650 : HS65_LHS_XOR2X3 port map( A => n2635, B => a(15), Z => n2914);
   U2651 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2921, Z => n1209);
   U2652 : HS65_LH_AO22X4 port map( A => n2565, B => n2511, C => n2564, D => 
                           n2923, Z => n2921);
   U2653 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2924, Z => n1208);
   U2654 : HS65_LH_AO222X4 port map( A => n2567, B => n2511, C => n2563, D => 
                           n2515, E => n1038, F => n2923, Z => n2924);
   U2655 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2926, Z => n1207);
   U2656 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1037, D1 => n2520, S1 
                           => n2564, D2 => n2515, S2 => n2566, D3 => n2511, S3 
                           => n2568, Z => n2926);
   U2657 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2928, Z => n1206);
   U2658 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1036, D1 => n2519, S1 
                           => n2566, D2 => n2515, S2 => n2568, D3 => n2511, S3 
                           => n2570, Z => n2928);
   U2659 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2929, Z => n1205);
   U2660 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1035, D1 => n2519, S1 
                           => n2568, D2 => n2515, S2 => n2570, D3 => n2511, S3 
                           => n2572, Z => n2929);
   U2661 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2930, Z => n1204);
   U2662 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1034, D1 => n2519, S1 
                           => n2570, D2 => n2515, S2 => n2572, D3 => n2511, S3 
                           => n2574, Z => n2930);
   U2663 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2931, Z => n1203);
   U2664 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1033, D1 => n2519, S1 
                           => n2572, D2 => n2515, S2 => n2574, D3 => n2511, S3 
                           => n2576, Z => n2931);
   U2665 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2932, Z => n1202);
   U2666 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1032, D1 => n2519, S1 
                           => n2574, D2 => n2515, S2 => n2576, D3 => n2511, S3 
                           => n2578, Z => n2932);
   U2667 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2933, Z => n1201);
   U2668 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1031, D1 => n2519, S1 
                           => n2576, D2 => n2515, S2 => n2578, D3 => n2511, S3 
                           => n2580, Z => n2933);
   U2669 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2934, Z => n1200);
   U2670 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1030, D1 => n2519, S1 
                           => n2578, D2 => n2516, S2 => n2580, D3 => n2511, S3 
                           => n2582, Z => n2934);
   U2671 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2935, Z => n1199);
   U2672 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1029, D1 => n2519, S1 
                           => n2580, D2 => n2515, S2 => n2582, D3 => n2511, S3 
                           => n2584, Z => n2935);
   U2673 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2936, Z => n1198);
   U2674 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1028, D1 => n2519, S1 
                           => n2582, D2 => n2515, S2 => n2584, D3 => n2511, S3 
                           => n2586, Z => n2936);
   U2675 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2937, Z => n1197);
   U2676 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1027, D1 => n2519, S1 
                           => n2584, D2 => n2515, S2 => n2586, D3 => n2511, S3 
                           => n2589, Z => n2937);
   U2677 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2938, Z => n1196);
   U2678 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1026, D1 => n2519, S1 
                           => n2586, D2 => n2516, S2 => n2588, D3 => n2511, S3 
                           => n2591, Z => n2938);
   U2679 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2939, Z => n1195);
   U2680 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1025, D1 => n2519, S1 
                           => n2588, D2 => n2516, S2 => n2590, D3 => n2511, S3 
                           => n2592, Z => n2939);
   U2681 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2940, Z => n1194);
   U2682 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1024, D1 => n2520, S1 
                           => n2590, D2 => n2516, S2 => n2592, D3 => n2511, S3 
                           => n2594, Z => n2940);
   U2683 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2941, Z => n1193);
   U2684 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1023, D1 => n2520, S1 
                           => n2592, D2 => n2516, S2 => n2594, D3 => n2511, S3 
                           => n2596, Z => n2941);
   U2685 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2942, Z => n1192);
   U2686 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1022, D1 => n2520, S1 
                           => n2594, D2 => n2516, S2 => n2596, D3 => n2512, S3 
                           => n2598, Z => n2942);
   U2687 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2943, Z => n1191);
   U2688 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1021, D1 => n2520, S1 
                           => n2596, D2 => n2516, S2 => n2598, D3 => n2512, S3 
                           => n2601, Z => n2943);
   U2689 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2944, Z => n1190);
   U2690 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1020, D1 => n2520, S1 
                           => n2598, D2 => n2516, S2 => n2600, D3 => n2512, S3 
                           => n2603, Z => n2944);
   U2691 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2945, Z => n1189);
   U2692 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1019, D1 => n2520, S1 
                           => n2600, D2 => n2516, S2 => n2602, D3 => n2512, S3 
                           => n2605, Z => n2945);
   U2693 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2946, Z => n1188);
   U2694 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1018, D1 => n2520, S1 
                           => n2602, D2 => n2516, S2 => n2604, D3 => n2512, S3 
                           => n2606, Z => n2946);
   U2695 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2947, Z => n1187);
   U2696 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1017, D1 => n2520, S1 
                           => n2604, D2 => n2516, S2 => n2606, D3 => n2512, S3 
                           => n2608, Z => n2947);
   U2697 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2948, Z => n1186);
   U2698 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1016, D1 => n2520, S1 
                           => n2606, D2 => n2516, S2 => n2608, D3 => n2512, S3 
                           => n2610, Z => n2948);
   U2699 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2949, Z => n1185);
   U2700 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1015, D1 => n2520, S1 
                           => n2608, D2 => n2516, S2 => n2610, D3 => n2512, S3 
                           => n2613, Z => n2949);
   U2701 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2950, Z => n1184);
   U2702 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1014, D1 => n2520, S1 
                           => n2610, D2 => n2516, S2 => n2612, D3 => n2512, S3 
                           => n2615, Z => n2950);
   U2703 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2951, Z => n1183);
   U2704 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1013, D1 => n2520, S1 
                           => n2612, D2 => n2517, S2 => n2614, D3 => n2512, S3 
                           => n2617, Z => n2951);
   U2705 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2952, Z => n1182);
   U2706 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1012, D1 => n2521, S1 
                           => n2614, D2 => n2517, S2 => n2616, D3 => n2512, S3 
                           => n2618, Z => n2952);
   U2707 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2953, Z => n1181);
   U2708 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1011, D1 => n2521, S1 
                           => n2616, D2 => n2517, S2 => n2618, D3 => n2512, S3 
                           => n2620, Z => n2953);
   U2709 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2954, Z => n1180);
   U2710 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1010, D1 => n2521, S1 
                           => n2618, D2 => n2517, S2 => n2620, D3 => n2512, S3 
                           => n2622, Z => n2954);
   U2711 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2955, Z => n1179);
   U2712 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1009, D1 => n2521, S1 
                           => n2620, D2 => n2517, S2 => n2622, D3 => n2512, S3 
                           => n2624, Z => n2955);
   U2713 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2956, Z => n1178);
   U2714 : HS65_LH_MX41X4 port map( D0 => n2923, S0 => n1008, D1 => n2521, S1 
                           => n2622, D2 => n2515, S2 => n2624, D3 => n2512, S3 
                           => n2626, Z => n2956);
   U2715 : HS65_LH_AND2X4 port map( A => n2957, B => n2958, Z => n2922);
   U2716 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2959, Z => n1177);
   U2717 : HS65_LH_OAI12X2 port map( A => n2657, B => n2514, C => n2960, Z => 
                           n2959);
   U2718 : HS65_LH_OAI22X1 port map( A => n2625, B => n2961, C => n2519, D => 
                           n2961, Z => n2960);
   U2719 : HS65_LH_AND2X4 port map( A => n2515, B => n2626, Z => n2961);
   U2720 : HS65_LH_NOR2X2 port map( A => n2957, B => n2962, Z => n2925);
   U2721 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2963, Z => n1176);
   U2722 : HS65_LH_AOI22X1 port map( A => n2923, B => n1006, C => n2521, D => 
                           n2627, Z => n2963);
   U2723 : HS65_LH_NOR3AX2 port map( A => n2962, B => n2958, C => n2957, Z => 
                           n2927);
   U2724 : HS65_LHS_XNOR2X3 port map( A => a(19), B => a(18), Z => n2962);
   U2725 : HS65_LH_NOR2AX3 port map( A => n2957, B => n2958, Z => n2923);
   U2726 : HS65_LHS_XNOR2X3 port map( A => n2639, B => a(19), Z => n2958);
   U2727 : HS65_LHS_XOR2X3 port map( A => n2637, B => a(18), Z => n2957);
   U2728 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2964, Z => n1174);
   U2729 : HS65_LH_AO22X4 port map( A => n2565, B => n2524, C => n2564, D => 
                           n2966, Z => n2964);
   U2730 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2967, Z => n1173);
   U2731 : HS65_LH_AO222X4 port map( A => n2567, B => n2524, C => n2563, D => 
                           n2528, E => n1038, F => n2966, Z => n2967);
   U2732 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2969, Z => n1172);
   U2733 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1037, D1 => n2524, S1 
                           => n2568, D2 => n2533, S2 => n2563, D3 => n2528, S3 
                           => n2566, Z => n2969);
   U2734 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2971, Z => n1171);
   U2735 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1036, D1 => n2524, S1 
                           => n2570, D2 => n2532, S2 => n2566, D3 => n2528, S3 
                           => n2568, Z => n2971);
   U2736 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2972, Z => n1170);
   U2737 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1035, D1 => n2524, S1 
                           => n2572, D2 => n2532, S2 => n2568, D3 => n2528, S3 
                           => n2570, Z => n2972);
   U2738 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2973, Z => n1169);
   U2739 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1034, D1 => n2524, S1 
                           => n2574, D2 => n2532, S2 => n2570, D3 => n2528, S3 
                           => n2572, Z => n2973);
   U2740 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2974, Z => n1168);
   U2741 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1033, D1 => n2524, S1 
                           => n2576, D2 => n2532, S2 => n2572, D3 => n2528, S3 
                           => n2574, Z => n2974);
   U2742 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2975, Z => n1167);
   U2743 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1032, D1 => n2524, S1 
                           => n2578, D2 => n2532, S2 => n2574, D3 => n2528, S3 
                           => n2576, Z => n2975);
   U2744 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2976, Z => n1166);
   U2745 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1031, D1 => n2524, S1 
                           => n2580, D2 => n2532, S2 => n2576, D3 => n2528, S3 
                           => n2578, Z => n2976);
   U2746 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2977, Z => n1165);
   U2747 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1030, D1 => n2524, S1 
                           => n2582, D2 => n2532, S2 => n2578, D3 => n2529, S3 
                           => n2580, Z => n2977);
   U2748 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2978, Z => n1164);
   U2749 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1029, D1 => n2524, S1 
                           => n2584, D2 => n2532, S2 => n2580, D3 => n2528, S3 
                           => n2582, Z => n2978);
   U2750 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2979, Z => n1163);
   U2751 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1028, D1 => n2524, S1 
                           => n2586, D2 => n2532, S2 => n2582, D3 => n2528, S3 
                           => n2584, Z => n2979);
   U2752 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2980, Z => n1162);
   U2753 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1027, D1 => n2524, S1 
                           => n2588, D2 => n2532, S2 => n2584, D3 => n2528, S3 
                           => n2586, Z => n2980);
   U2754 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2981, Z => n1161);
   U2755 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1026, D1 => n2524, S1 
                           => n2590, D2 => n2532, S2 => n2586, D3 => n2529, S3 
                           => n2588, Z => n2981);
   U2756 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2982, Z => n1160);
   U2757 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1025, D1 => n2524, S1 
                           => n2592, D2 => n2532, S2 => n2588, D3 => n2529, S3 
                           => n2590, Z => n2982);
   U2758 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2983, Z => n1159);
   U2759 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1024, D1 => n2524, S1 
                           => n2594, D2 => n2533, S2 => n2590, D3 => n2529, S3 
                           => n2592, Z => n2983);
   U2760 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2984, Z => n1158);
   U2761 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1023, D1 => n2525, S1 
                           => n2596, D2 => n2533, S2 => n2592, D3 => n2529, S3 
                           => n2594, Z => n2984);
   U2762 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2985, Z => n1157);
   U2763 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1022, D1 => n2525, S1 
                           => n2598, D2 => n2533, S2 => n2594, D3 => n2529, S3 
                           => n2596, Z => n2985);
   U2764 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2986, Z => n1156);
   U2765 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1021, D1 => n2525, S1 
                           => n2600, D2 => n2533, S2 => n2596, D3 => n2529, S3 
                           => n2598, Z => n2986);
   U2766 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2987, Z => n1155);
   U2767 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1020, D1 => n2525, S1 
                           => n2602, D2 => n2533, S2 => n2598, D3 => n2529, S3 
                           => n2600, Z => n2987);
   U2768 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2988, Z => n1154);
   U2769 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1019, D1 => n2525, S1 
                           => n2604, D2 => n2533, S2 => n2600, D3 => n2529, S3 
                           => n2602, Z => n2988);
   U2770 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2989, Z => n1153);
   U2771 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1018, D1 => n2525, S1 
                           => n2606, D2 => n2533, S2 => n2602, D3 => n2529, S3 
                           => n2604, Z => n2989);
   U2772 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2990, Z => n1152);
   U2773 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1017, D1 => n2525, S1 
                           => n2608, D2 => n2533, S2 => n2604, D3 => n2529, S3 
                           => n2606, Z => n2990);
   U2774 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2991, Z => n1151);
   U2775 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1016, D1 => n2525, S1 
                           => n2610, D2 => n2533, S2 => n2606, D3 => n2529, S3 
                           => n2608, Z => n2991);
   U2776 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2992, Z => n1150);
   U2777 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1015, D1 => n2525, S1 
                           => n2612, D2 => n2533, S2 => n2608, D3 => n2529, S3 
                           => n2610, Z => n2992);
   U2778 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2993, Z => n1149);
   U2779 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1014, D1 => n2525, S1 
                           => n2614, D2 => n2533, S2 => n2610, D3 => n2529, S3 
                           => n2612, Z => n2993);
   U2780 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2994, Z => n1148);
   U2781 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1013, D1 => n2525, S1 
                           => n2616, D2 => n2533, S2 => n2612, D3 => n2530, S3 
                           => n2614, Z => n2994);
   U2782 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2995, Z => n1147);
   U2783 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1012, D1 => n2525, S1 
                           => n2618, D2 => n2533, S2 => n2614, D3 => n2530, S3 
                           => n2616, Z => n2995);
   U2784 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2996, Z => n1146);
   U2785 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1011, D1 => n2525, S1 
                           => n2620, D2 => n2534, S2 => n2616, D3 => n2530, S3 
                           => n2618, Z => n2996);
   U2786 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2997, Z => n1145);
   U2787 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1010, D1 => n2525, S1 
                           => n2622, D2 => n2534, S2 => n2618, D3 => n2530, S3 
                           => n2620, Z => n2997);
   U2788 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2998, Z => n1144);
   U2789 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1009, D1 => n2525, S1 
                           => n2624, D2 => n2534, S2 => n2620, D3 => n2530, S3 
                           => n2622, Z => n2998);
   U2790 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2999, Z => n1143);
   U2791 : HS65_LH_MX41X4 port map( D0 => n2966, S0 => n1008, D1 => n2525, S1 
                           => n2626, D2 => n2534, S2 => n2622, D3 => n2528, S3 
                           => n2624, Z => n2999);
   U2792 : HS65_LH_AND2X4 port map( A => n3000, B => n3001, Z => n2965);
   U2793 : HS65_LHS_XOR2X3 port map( A => a(23), B => n3002, Z => n1142);
   U2794 : HS65_LH_OAI12X2 port map( A => n2657, B => n2527, C => n3003, Z => 
                           n3002);
   U2795 : HS65_LH_OAI22X1 port map( A => n2625, B => n3004, C => n2532, D => 
                           n3004, Z => n3003);
   U2796 : HS65_LH_AND2X4 port map( A => n2528, B => n2626, Z => n3004);
   U2797 : HS65_LH_NOR2X2 port map( A => n3000, B => n3005, Z => n2968);
   U2798 : HS65_LHS_XOR2X3 port map( A => n2642, B => n3006, Z => n1141);
   U2799 : HS65_LH_AOI22X1 port map( A => n2966, B => n1006, C => n2534, D => 
                           n2627, Z => n3006);
   U2800 : HS65_LH_NOR3AX2 port map( A => n3005, B => n3001, C => n3000, Z => 
                           n2970);
   U2801 : HS65_LHS_XNOR2X3 port map( A => a(22), B => a(21), Z => n3005);
   U2802 : HS65_LH_NOR2AX3 port map( A => n3000, B => n3001, Z => n2966);
   U2803 : HS65_LHS_XNOR2X3 port map( A => n2641, B => a(22), Z => n3001);
   U2804 : HS65_LHS_XOR2X3 port map( A => n2639, B => a(21), Z => n3000);
   U2805 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3007, Z => n1139);
   U2806 : HS65_LH_AO22X4 port map( A => n2565, B => n2537, C => n2564, D => 
                           n3009, Z => n3007);
   U2807 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3010, Z => n1138);
   U2808 : HS65_LH_AO222X4 port map( A => n2567, B => n2537, C => n2563, D => 
                           n2541, E => n1038, F => n3009, Z => n3010);
   U2809 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3012, Z => n1137);
   U2810 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1037, D1 => n2546, S1 
                           => n2563, D2 => n2541, S2 => n2566, D3 => n2537, S3 
                           => n2568, Z => n3012);
   U2811 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3014, Z => n1136);
   U2812 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1036, D1 => n2545, S1 
                           => n2567, D2 => n2541, S2 => n2568, D3 => n2537, S3 
                           => n2570, Z => n3014);
   U2813 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3015, Z => n1135);
   U2814 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1035, D1 => n2545, S1 
                           => n2568, D2 => n2541, S2 => n2570, D3 => n2537, S3 
                           => n2572, Z => n3015);
   U2815 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3016, Z => n1134);
   U2816 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1034, D1 => n2545, S1 
                           => n2570, D2 => n2541, S2 => n2572, D3 => n2537, S3 
                           => n2574, Z => n3016);
   U2817 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3017, Z => n1133);
   U2818 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1033, D1 => n2545, S1 
                           => n2572, D2 => n2541, S2 => n2574, D3 => n2537, S3 
                           => n2576, Z => n3017);
   U2819 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3018, Z => n1132);
   U2820 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1032, D1 => n2545, S1 
                           => n2574, D2 => n2541, S2 => n2576, D3 => n2537, S3 
                           => n2578, Z => n3018);
   U2821 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3019, Z => n1131);
   U2822 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1031, D1 => n2545, S1 
                           => n2576, D2 => n2541, S2 => n2578, D3 => n2537, S3 
                           => n2580, Z => n3019);
   U2823 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3020, Z => n1130);
   U2824 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1030, D1 => n2545, S1 
                           => n2578, D2 => n2542, S2 => n2580, D3 => n2537, S3 
                           => n2582, Z => n3020);
   U2825 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3021, Z => n1129);
   U2826 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1029, D1 => n2545, S1 
                           => n2580, D2 => n2541, S2 => n2582, D3 => n2537, S3 
                           => n2584, Z => n3021);
   U2827 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3022, Z => n1128);
   U2828 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1028, D1 => n2545, S1 
                           => n2582, D2 => n2541, S2 => n2584, D3 => n2537, S3 
                           => n2586, Z => n3022);
   U2829 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3023, Z => n1127);
   U2830 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1027, D1 => n2545, S1 
                           => n2584, D2 => n2541, S2 => n2586, D3 => n2537, S3 
                           => n2588, Z => n3023);
   U2831 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3024, Z => n1126);
   U2832 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1026, D1 => n2545, S1 
                           => n2586, D2 => n2542, S2 => n2588, D3 => n2537, S3 
                           => n2590, Z => n3024);
   U2833 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3025, Z => n1125);
   U2834 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1025, D1 => n2545, S1 
                           => n2588, D2 => n2542, S2 => n2590, D3 => n2537, S3 
                           => n2592, Z => n3025);
   U2835 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3026, Z => n1124);
   U2836 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1024, D1 => n2546, S1 
                           => n2590, D2 => n2542, S2 => n2592, D3 => n2537, S3 
                           => n2594, Z => n3026);
   U2837 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3027, Z => n1123);
   U2838 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1023, D1 => n2546, S1 
                           => n2592, D2 => n2542, S2 => n2594, D3 => n2537, S3 
                           => n2596, Z => n3027);
   U2839 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3028, Z => n1122);
   U2840 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1022, D1 => n2546, S1 
                           => n2594, D2 => n2542, S2 => n2596, D3 => n2538, S3 
                           => n2598, Z => n3028);
   U2841 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3029, Z => n1121);
   U2842 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1021, D1 => n2546, S1 
                           => n2596, D2 => n2542, S2 => n2598, D3 => n2538, S3 
                           => n2600, Z => n3029);
   U2843 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3030, Z => n1120);
   U2844 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1020, D1 => n2546, S1 
                           => n2598, D2 => n2542, S2 => n2600, D3 => n2538, S3 
                           => n2602, Z => n3030);
   U2845 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3031, Z => n1119);
   U2846 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1019, D1 => n2546, S1 
                           => n2600, D2 => n2542, S2 => n2602, D3 => n2538, S3 
                           => n2604, Z => n3031);
   U2847 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3032, Z => n1118);
   U2848 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1018, D1 => n2546, S1 
                           => n2602, D2 => n2542, S2 => n2604, D3 => n2538, S3 
                           => n2606, Z => n3032);
   U2849 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3033, Z => n1117);
   U2850 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1017, D1 => n2546, S1 
                           => n2604, D2 => n2542, S2 => n2606, D3 => n2538, S3 
                           => n2608, Z => n3033);
   U2851 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3034, Z => n1116);
   U2852 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1016, D1 => n2546, S1 
                           => n2606, D2 => n2542, S2 => n2608, D3 => n2538, S3 
                           => n2610, Z => n3034);
   U2853 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3035, Z => n1115);
   U2854 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1015, D1 => n2546, S1 
                           => n2608, D2 => n2542, S2 => n2610, D3 => n2538, S3 
                           => n2612, Z => n3035);
   U2855 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3036, Z => n1114);
   U2856 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1014, D1 => n2546, S1 
                           => n2610, D2 => n2542, S2 => n2612, D3 => n2538, S3 
                           => n2614, Z => n3036);
   U2857 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3037, Z => n1113);
   U2858 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1013, D1 => n2546, S1 
                           => n2612, D2 => n2543, S2 => n2614, D3 => n2538, S3 
                           => n2616, Z => n3037);
   U2859 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3038, Z => n1112);
   U2860 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1012, D1 => n2547, S1 
                           => n2614, D2 => n2543, S2 => n2616, D3 => n2538, S3 
                           => n2618, Z => n3038);
   U2861 : HS65_LHS_XOR2X3 port map( A => n2643, B => n3039, Z => n1111);
   U2862 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1011, D1 => n2547, S1 
                           => n2616, D2 => n2543, S2 => n2618, D3 => n2538, S3 
                           => n2620, Z => n3039);
   U2863 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3040, Z => n1110);
   U2864 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1010, D1 => n2547, S1 
                           => n2618, D2 => n2543, S2 => n2620, D3 => n2538, S3 
                           => n2622, Z => n3040);
   U2865 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3041, Z => n1109);
   U2866 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1009, D1 => n2547, S1 
                           => n2620, D2 => n2543, S2 => n2622, D3 => n2538, S3 
                           => n2624, Z => n3041);
   U2867 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3042, Z => n1108);
   U2868 : HS65_LH_MX41X4 port map( D0 => n3009, S0 => n1008, D1 => n2547, S1 
                           => n2622, D2 => n2541, S2 => n2624, D3 => n2538, S3 
                           => n2626, Z => n3042);
   U2869 : HS65_LH_AND2X4 port map( A => n3043, B => n3044, Z => n3008);
   U2870 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3045, Z => n1107);
   U2871 : HS65_LH_OAI12X2 port map( A => n2657, B => n2540, C => n3046, Z => 
                           n3045);
   U2872 : HS65_LH_OAI22X1 port map( A => n2625, B => n3047, C => n2545, D => 
                           n3047, Z => n3046);
   U2873 : HS65_LH_AND2X4 port map( A => n2541, B => n2626, Z => n3047);
   U2874 : HS65_LH_NOR2X2 port map( A => n3043, B => n3048, Z => n3011);
   U2875 : HS65_LHS_XOR2X3 port map( A => n2644, B => n3049, Z => n1106);
   U2876 : HS65_LH_AOI22X1 port map( A => n3009, B => n1006, C => n2547, D => 
                           n2627, Z => n3049);
   U2877 : HS65_LH_NOR3AX2 port map( A => n3048, B => n3044, C => n3043, Z => 
                           n3013);
   U2878 : HS65_LHS_XNOR2X3 port map( A => a(25), B => a(24), Z => n3048);
   U2879 : HS65_LH_NOR2AX3 port map( A => n3043, B => n3044, Z => n3009);
   U2880 : HS65_LHS_XNOR2X3 port map( A => n2643, B => a(25), Z => n3044);
   U2881 : HS65_LHS_XOR2X3 port map( A => n2641, B => a(24), Z => n3043);
   U2882 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3050, Z => n1104);
   U2883 : HS65_LH_AO22X4 port map( A => n2565, B => n2550, C => n2564, D => 
                           n3052, Z => n3050);
   U2884 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3053, Z => n1103);
   U2885 : HS65_LH_AO222X4 port map( A => n2567, B => n2550, C => n2563, D => 
                           n2554, E => n1038, F => n3052, Z => n3053);
   U2886 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3055, Z => n1102);
   U2887 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1037, D1 => n2559, S1 
                           => n2563, D2 => n2554, S2 => n2566, D3 => n2550, S3 
                           => n2568, Z => n3055);
   U2888 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3057, Z => n1101);
   U2889 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1036, D1 => n2558, S1 
                           => n2567, D2 => n2554, S2 => n2568, D3 => n2550, S3 
                           => n2570, Z => n3057);
   U2890 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3058, Z => n1100);
   U2891 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1035, D1 => n2558, S1 
                           => n2568, D2 => n2554, S2 => n2570, D3 => n2550, S3 
                           => n2572, Z => n3058);
   U2892 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3059, Z => n1099);
   U2893 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1034, D1 => n2558, S1 
                           => n2570, D2 => n2554, S2 => n2572, D3 => n2550, S3 
                           => n2574, Z => n3059);
   U2894 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3060, Z => n1098);
   U2895 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1033, D1 => n2558, S1 
                           => n2572, D2 => n2554, S2 => n2574, D3 => n2550, S3 
                           => n2576, Z => n3060);
   U2896 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3061, Z => n1097);
   U2897 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1032, D1 => n2558, S1 
                           => n2574, D2 => n2554, S2 => n2576, D3 => n2550, S3 
                           => n2578, Z => n3061);
   U2898 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3062, Z => n1096);
   U2899 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1031, D1 => n2558, S1 
                           => n2576, D2 => n2554, S2 => n2578, D3 => n2550, S3 
                           => n2580, Z => n3062);
   U2900 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3063, Z => n1095);
   U2901 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1030, D1 => n2558, S1 
                           => n2578, D2 => n2555, S2 => n2580, D3 => n2550, S3 
                           => n2582, Z => n3063);
   U2902 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3064, Z => n1094);
   U2903 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1029, D1 => n2558, S1 
                           => n2580, D2 => n2554, S2 => n2582, D3 => n2550, S3 
                           => n2584, Z => n3064);
   U2904 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3065, Z => n1093);
   U2905 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1028, D1 => n2558, S1 
                           => n2582, D2 => n2554, S2 => n2584, D3 => n2550, S3 
                           => n2586, Z => n3065);
   U2906 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3066, Z => n1092);
   U2907 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1027, D1 => n2558, S1 
                           => n2584, D2 => n2554, S2 => n2586, D3 => n2550, S3 
                           => n2588, Z => n3066);
   U2908 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3067, Z => n1091);
   U2909 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1026, D1 => n2558, S1 
                           => n2586, D2 => n2555, S2 => n2588, D3 => n2550, S3 
                           => n2590, Z => n3067);
   U2910 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3068, Z => n1090);
   U2911 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1025, D1 => n2558, S1 
                           => n2588, D2 => n2555, S2 => n2590, D3 => n2550, S3 
                           => n2592, Z => n3068);
   U2912 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3069, Z => n1089);
   U2913 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1024, D1 => n2559, S1 
                           => n2590, D2 => n2555, S2 => n2592, D3 => n2550, S3 
                           => n2594, Z => n3069);
   U2914 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3070, Z => n1088);
   U2915 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1023, D1 => n2559, S1 
                           => n2592, D2 => n2555, S2 => n2594, D3 => n2550, S3 
                           => n2596, Z => n3070);
   U2916 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3071, Z => n1087);
   U2917 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1022, D1 => n2559, S1 
                           => n2594, D2 => n2555, S2 => n2596, D3 => n2551, S3 
                           => n2598, Z => n3071);
   U2918 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3072, Z => n1086);
   U2919 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1021, D1 => n2559, S1 
                           => n2596, D2 => n2555, S2 => n2598, D3 => n2551, S3 
                           => n2600, Z => n3072);
   U2920 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3073, Z => n1085);
   U2921 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1020, D1 => n2559, S1 
                           => n2598, D2 => n2555, S2 => n2600, D3 => n2551, S3 
                           => n2602, Z => n3073);
   U2922 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3074, Z => n1084);
   U2923 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1019, D1 => n2559, S1 
                           => n2600, D2 => n2555, S2 => n2602, D3 => n2551, S3 
                           => n2604, Z => n3074);
   U2924 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3075, Z => n1083);
   U2925 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1018, D1 => n2559, S1 
                           => n2602, D2 => n2555, S2 => n2604, D3 => n2551, S3 
                           => n2606, Z => n3075);
   U2926 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3076, Z => n1082);
   U2927 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1017, D1 => n2559, S1 
                           => n2604, D2 => n2555, S2 => n2606, D3 => n2551, S3 
                           => n2608, Z => n3076);
   U2928 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3077, Z => n1081);
   U2929 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1016, D1 => n2559, S1 
                           => n2606, D2 => n2555, S2 => n2608, D3 => n2551, S3 
                           => n2610, Z => n3077);
   U2930 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3078, Z => n1080);
   U2931 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1015, D1 => n2559, S1 
                           => n2608, D2 => n2555, S2 => n2610, D3 => n2551, S3 
                           => n2612, Z => n3078);
   U2932 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3079, Z => n1079);
   U2933 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1014, D1 => n2559, S1 
                           => n2610, D2 => n2555, S2 => n2612, D3 => n2551, S3 
                           => n2614, Z => n3079);
   U2934 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3080, Z => n1078);
   U2935 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1013, D1 => n2559, S1 
                           => n2612, D2 => n2556, S2 => n2614, D3 => n2551, S3 
                           => n2616, Z => n3080);
   U2936 : HS65_LHS_XOR2X3 port map( A => n2645, B => n3081, Z => n1077);
   U2937 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1012, D1 => n2560, S1 
                           => n2614, D2 => n2556, S2 => n2616, D3 => n2551, S3 
                           => n2618, Z => n3081);
   U2938 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3082, Z => n1076);
   U2939 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1011, D1 => n2560, S1 
                           => n2616, D2 => n2556, S2 => n2618, D3 => n2551, S3 
                           => n2620, Z => n3082);
   U2940 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3083, Z => n1075);
   U2941 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1010, D1 => n2560, S1 
                           => n2618, D2 => n2556, S2 => n2620, D3 => n2551, S3 
                           => n2622, Z => n3083);
   U2942 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3084, Z => n1074);
   U2943 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1009, D1 => n2560, S1 
                           => n2620, D2 => n2556, S2 => n2622, D3 => n2551, S3 
                           => n2624, Z => n3084);
   U2944 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3085, Z => n1073);
   U2945 : HS65_LH_MX41X4 port map( D0 => n3052, S0 => n1008, D1 => n2560, S1 
                           => n2622, D2 => n2554, S2 => n2624, D3 => n2551, S3 
                           => n2626, Z => n3085);
   U2946 : HS65_LH_AND2X4 port map( A => n3086, B => n3087, Z => n3051);
   U2947 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3088, Z => n1072);
   U2948 : HS65_LH_OAI12X2 port map( A => n2657, B => n2553, C => n3089, Z => 
                           n3088);
   U2949 : HS65_LH_OAI22X1 port map( A => n2625, B => n3090, C => n2558, D => 
                           n3090, Z => n3089);
   U2950 : HS65_LH_AND2X4 port map( A => n2554, B => n2626, Z => n3090);
   U2951 : HS65_LH_NOR2X2 port map( A => n3086, B => n3091, Z => n3054);
   U2952 : HS65_LHS_XOR2X3 port map( A => n2646, B => n3092, Z => n1071);
   U2953 : HS65_LH_AOI22X1 port map( A => n3052, B => n1006, C => n2560, D => 
                           n2627, Z => n3092);
   U2954 : HS65_LH_NOR3AX2 port map( A => n3091, B => n3087, C => n3086, Z => 
                           n3056);
   U2955 : HS65_LHS_XNOR2X3 port map( A => a(28), B => a(27), Z => n3091);
   U2956 : HS65_LH_NOR2AX3 port map( A => n3086, B => n3087, Z => n3052);
   U2957 : HS65_LHS_XNOR2X3 port map( A => a(29), B => a(28), Z => n3087);
   U2958 : HS65_LHS_XOR2X3 port map( A => n2643, B => a(27), Z => n3086);
   U2959 : HS65_LH_AO22X4 port map( A => n2428, B => n2563, C => n2419, D => 
                           n2564, Z => n1069);
   U2960 : HS65_LH_AO222X4 port map( A => n2428, B => n2566, C => n2432, D => 
                           n2563, E => n2419, F => n1038, Z => n1068);
   U2961 : HS65_LH_MX41X4 port map( D0 => n1037, S0 => n2419, D1 => n2569, S1 
                           => n2426, D2 => n2567, S2 => n2430, D3 => n2564, S3 
                           => n2423, Z => n1067);
   U2962 : HS65_LH_MX41X4 port map( D0 => n1036, S0 => n2419, D1 => n2571, S1 
                           => n2426, D2 => n2569, S2 => n2430, D3 => n2567, S3 
                           => n2423, Z => n1066);
   U2963 : HS65_LH_MX41X4 port map( D0 => n1035, S0 => n2419, D1 => n2573, S1 
                           => n2426, D2 => n2571, S2 => n2430, D3 => n2569, S3 
                           => n2423, Z => n1065);
   U2964 : HS65_LH_MX41X4 port map( D0 => n1034, S0 => n2418, D1 => n2575, S1 
                           => n2426, D2 => n2573, S2 => n2430, D3 => n2571, S3 
                           => n2423, Z => n1064);
   U2965 : HS65_LH_MX41X4 port map( D0 => n1033, S0 => n2418, D1 => n2577, S1 
                           => n2426, D2 => n2575, S2 => n2430, D3 => n2573, S3 
                           => n2423, Z => n1063);
   U2966 : HS65_LH_MX41X4 port map( D0 => n1032, S0 => n2418, D1 => n2579, S1 
                           => n2426, D2 => n2577, S2 => n2430, D3 => n2575, S3 
                           => n2423, Z => n1062);
   U2967 : HS65_LH_MX41X4 port map( D0 => n1031, S0 => n2418, D1 => n2581, S1 
                           => n2426, D2 => n2579, S2 => n2430, D3 => n2577, S3 
                           => n2423, Z => n1061);
   U2968 : HS65_LH_MX41X4 port map( D0 => n1030, S0 => n2418, D1 => n2583, S1 
                           => n2426, D2 => n2581, S2 => n2430, D3 => n2579, S3 
                           => n2423, Z => n1060);
   U2969 : HS65_LH_MX41X4 port map( D0 => n1029, S0 => n2418, D1 => n2585, S1 
                           => n2426, D2 => n2583, S2 => n2430, D3 => n2581, S3 
                           => n2423, Z => n1059);
   U2970 : HS65_LH_MX41X4 port map( D0 => n1028, S0 => n2418, D1 => n2587, S1 
                           => n2426, D2 => n2585, S2 => n2431, D3 => n2583, S3 
                           => n2424, Z => n1058);
   U2971 : HS65_LH_MX41X4 port map( D0 => n1027, S0 => n2418, D1 => n2428, S1 
                           => n2588, D2 => n2587, S2 => n2431, D3 => n2585, S3 
                           => n2424, Z => n1057);
   U2972 : HS65_LH_MX41X4 port map( D0 => n1026, S0 => n2418, D1 => n2428, S1 
                           => n2590, D2 => n2589, S2 => n2431, D3 => n2587, S3 
                           => n2424, Z => n1056);
   U2973 : HS65_LH_MX41X4 port map( D0 => n1024, S0 => n2418, D1 => n2593, S1 
                           => n2432, D2 => n2591, S2 => n2423, D3 => n2595, S3 
                           => n2426, Z => n1055);
   U2974 : HS65_LH_MX41X4 port map( D0 => n1023, S0 => n2418, D1 => n2593, S1 
                           => n2424, D2 => n2595, S2 => n2431, D3 => n2597, S3 
                           => n2427, Z => n1054);
   U2975 : HS65_LH_MX41X4 port map( D0 => n1022, S0 => n2417, D1 => n2595, S1 
                           => n2424, D2 => n2597, S2 => n2431, D3 => n2599, S3 
                           => n2427, Z => n1053);
   U2976 : HS65_LH_MX41X4 port map( D0 => n1021, S0 => n2417, D1 => n2597, S1 
                           => n2424, D2 => n2599, S2 => n2431, D3 => n2601, S3 
                           => n2427, Z => n1052);
   U2977 : HS65_LH_MX41X4 port map( D0 => n1020, S0 => n2417, D1 => n2599, S1 
                           => n2424, D2 => n2601, S2 => n2431, D3 => n2603, S3 
                           => n2427, Z => n1051);
   U2978 : HS65_LH_MX41X4 port map( D0 => n1018, S0 => n2417, D1 => n2603, S1 
                           => n2424, D2 => n2605, S2 => n2431, D3 => n2607, S3 
                           => n2427, Z => n1050);
   U2979 : HS65_LH_MX41X4 port map( D0 => n1017, S0 => n2417, D1 => n2605, S1 
                           => n2424, D2 => n2607, S2 => n2431, D3 => n2609, S3 
                           => n2427, Z => n1049);
   U2980 : HS65_LH_MX41X4 port map( D0 => n1016, S0 => n2417, D1 => n2607, S1 
                           => n2424, D2 => n2609, S2 => n2431, D3 => n2611, S3 
                           => n2427, Z => n1048);
   U2981 : HS65_LH_MX41X4 port map( D0 => n1015, S0 => n2417, D1 => n2609, S1 
                           => n2424, D2 => n2611, S2 => n2431, D3 => n2613, S3 
                           => n2427, Z => n1047);
   U2982 : HS65_LH_MX41X4 port map( D0 => n1014, S0 => n2417, D1 => n2611, S1 
                           => n2424, D2 => n2613, S2 => n2432, D3 => n2615, S3 
                           => n2427, Z => n1046);
   U2983 : HS65_LH_MX41X4 port map( D0 => n1012, S0 => n2417, D1 => n2615, S1 
                           => n2424, D2 => n2617, S2 => n2432, D3 => n2619, S3 
                           => n2427, Z => n1045);
   U2984 : HS65_LH_MX41X4 port map( D0 => n1011, S0 => n2417, D1 => n2617, S1 
                           => n2424, D2 => n2619, S2 => n2432, D3 => n2621, S3 
                           => n2427, Z => n1044);
   U2985 : HS65_LH_MX41X4 port map( D0 => n1010, S0 => n2417, D1 => n2619, S1 
                           => n2424, D2 => n2621, S2 => n2432, D3 => n2623, S3 
                           => n2427, Z => n1043);
   U2986 : HS65_LH_MX41X4 port map( D0 => n1009, S0 => n2417, D1 => n2621, S1 
                           => n2423, D2 => n2623, S2 => n2431, D3 => n2625, S3 
                           => n2428, Z => n1042);
   U2987 : HS65_LH_MX41X4 port map( D0 => n1008, S0 => n2418, D1 => n2623, S1 
                           => n2424, D2 => n2625, S2 => n2430, D3 => n2428, S3 
                           => n2626, Z => n1041);
   U2988 : HS65_LH_NOR2AX3 port map( A => n3093, B => a(31), Z => n2660);
   U2989 : HS65_LH_NOR2AX3 port map( A => n3094, B => n3093, Z => n2661);
   U2990 : HS65_LH_NOR3AX2 port map( A => a(31), B => n3094, C => n3093, Z => 
                           n2659);
   U2991 : HS65_LHS_XOR2X3 port map( A => a(31), B => a(30), Z => n3094);
   U2992 : HS65_LH_NAND2X2 port map( A => a(31), B => n3093, Z => n2662);
   U2993 : HS65_LHS_XOR2X3 port map( A => n2645, B => a(30), Z => n3093);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_add_0;

architecture SYN_rpl of alu_DW01_add_0 is

   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1 : std_logic;

begin
   
   U1_31 : HS65_LHS_XOR3X2 port map( A => A(31), B => B(31), C => carry_31_port
                           , Z => SUM(31));
   U1_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => B(30), CI => 
                           carry_30_port, CO => carry_31_port, S0 => SUM(30));
   U1_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => B(28), CI => 
                           carry_28_port, CO => carry_29_port, S0 => SUM(28));
   U1_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => B(27), CI => 
                           carry_27_port, CO => carry_28_port, S0 => SUM(27));
   U1_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => B(25), CI => 
                           carry_25_port, CO => carry_26_port, S0 => SUM(25));
   U1_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => B(24), CI => 
                           carry_24_port, CO => carry_25_port, S0 => SUM(24));
   U1_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => B(22), CI => 
                           carry_22_port, CO => carry_23_port, S0 => SUM(22));
   U1_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => B(21), CI => 
                           carry_21_port, CO => carry_22_port, S0 => SUM(21));
   U1_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => B(19), CI => 
                           carry_19_port, CO => carry_20_port, S0 => SUM(19));
   U1_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => B(18), CI => 
                           carry_18_port, CO => carry_19_port, S0 => SUM(18));
   U1_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => B(16), CI => 
                           carry_16_port, CO => carry_17_port, S0 => SUM(16));
   U1_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => B(3), CI => carry_3_port, 
                           CO => carry_4_port, S0 => SUM(3));
   U1_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => B(1), CI => n1, CO => 
                           carry_2_port, S0 => SUM(1));
   U1_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => B(15), CI => 
                           carry_15_port, CO => carry_16_port, S0 => SUM(15));
   U1_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => B(13), CI => 
                           carry_13_port, CO => carry_14_port, S0 => SUM(13));
   U1_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => B(12), CI => 
                           carry_12_port, CO => carry_13_port, S0 => SUM(12));
   U1_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => B(10), CI => 
                           carry_10_port, CO => carry_11_port, S0 => SUM(10));
   U1_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => B(9), CI => carry_9_port, 
                           CO => carry_10_port, S0 => SUM(9));
   U1_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => B(7), CI => carry_7_port, 
                           CO => carry_8_port, S0 => SUM(7));
   U1_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => B(6), CI => carry_6_port, 
                           CO => carry_7_port, S0 => SUM(6));
   U1_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => B(4), CI => carry_4_port, 
                           CO => carry_5_port, S0 => SUM(4));
   U1_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => B(23), CI => 
                           carry_23_port, CO => carry_24_port, S0 => SUM(23));
   U1_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => B(2), CI => carry_2_port, 
                           CO => carry_3_port, S0 => SUM(2));
   U1_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => B(29), CI => 
                           carry_29_port, CO => carry_30_port, S0 => SUM(29));
   U1_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => B(26), CI => 
                           carry_26_port, CO => carry_27_port, S0 => SUM(26));
   U1_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => B(20), CI => 
                           carry_20_port, CO => carry_21_port, S0 => SUM(20));
   U1_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => B(17), CI => 
                           carry_17_port, CO => carry_18_port, S0 => SUM(17));
   U1_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => B(11), CI => 
                           carry_11_port, CO => carry_12_port, S0 => SUM(11));
   U1_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => B(5), CI => carry_5_port, 
                           CO => carry_6_port, S0 => SUM(5));
   U1_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => B(14), CI => 
                           carry_14_port, CO => carry_15_port, S0 => SUM(14));
   U1_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => B(8), CI => carry_8_port, 
                           CO => carry_9_port, S0 => SUM(8));
   U1 : HS65_LH_AND2X4 port map( A => A(0), B => B(0), Z => n1);
   U2 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => SUM(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end alu_DW01_cmp6_0;

architecture SYN_rpl of alu_DW01_cmp6_0 is

   component HS65_LH_NAND2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2AX4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND4X3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal LT_port, EQ_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115 : std_logic;

begin
   LT <= LT_port;
   EQ <= EQ_port;
   
   U1 : HS65_LH_IVX9 port map( A => n54, Z => n35);
   U2 : HS65_LH_IVX9 port map( A => EQ_port, Z => NE);
   U3 : HS65_LH_IVX9 port map( A => n115, Z => n40);
   U4 : HS65_LH_IVX9 port map( A => A(14), Z => n21);
   U5 : HS65_LH_IVX9 port map( A => A(26), Z => n22);
   U6 : HS65_LH_IVX9 port map( A => B(2), Z => n1);
   U7 : HS65_LH_IVX9 port map( A => B(3), Z => n2);
   U8 : HS65_LH_IVX9 port map( A => B(27), Z => n16);
   U9 : HS65_LH_IVX9 port map( A => B(20), Z => n12);
   U10 : HS65_LH_IVX9 port map( A => B(11), Z => n6);
   U11 : HS65_LH_IVX9 port map( A => A(8), Z => n20);
   U12 : HS65_LH_IVX9 port map( A => B(28), Z => n17);
   U13 : HS65_LH_IVX9 port map( A => B(31), Z => n19);
   U14 : HS65_LH_IVX9 port map( A => n102, Z => n38);
   U15 : HS65_LH_IVX9 port map( A => n67, Z => n27);
   U16 : HS65_LH_OR2X9 port map( A => B(26), B => n22, Z => n66);
   U17 : HS65_LH_OR2X9 port map( A => B(14), B => n21, Z => n50);
   U18 : HS65_LH_IVX9 port map( A => B(23), Z => n14);
   U19 : HS65_LH_IVX9 port map( A => B(19), Z => n11);
   U20 : HS65_LH_IVX9 port map( A => B(25), Z => n15);
   U21 : HS65_LH_IVX9 port map( A => B(12), Z => n7);
   U22 : HS65_LH_IVX9 port map( A => B(13), Z => n8);
   U23 : HS65_LH_IVX9 port map( A => B(21), Z => n13);
   U24 : HS65_LH_IVX9 port map( A => B(15), Z => n9);
   U25 : HS65_LH_IVX9 port map( A => B(7), Z => n4);
   U26 : HS65_LH_IVX9 port map( A => B(5), Z => n3);
   U27 : HS65_LH_IVX9 port map( A => B(29), Z => n18);
   U28 : HS65_LH_IVX9 port map( A => B(9), Z => n5);
   U29 : HS65_LH_IVX9 port map( A => B(17), Z => n10);
   U30 : HS65_LH_IVX9 port map( A => n76, Z => n24);
   U31 : HS65_LH_IVX9 port map( A => n60, Z => n25);
   U32 : HS65_LH_IVX9 port map( A => n64, Z => n28);
   U33 : HS65_LH_IVX9 port map( A => n51, Z => n37);
   U34 : HS65_LH_IVX9 port map( A => A(22), Z => n30);
   U35 : HS65_LH_IVX9 port map( A => A(6), Z => n39);
   U36 : HS65_LH_IVX9 port map( A => n71, Z => n33);
   U37 : HS65_LH_IVX9 port map( A => n70, Z => n31);
   U38 : HS65_LH_IVX9 port map( A => A(1), Z => n42);
   U39 : HS65_LH_IVX9 port map( A => A(18), Z => n32);
   U40 : HS65_LH_IVX9 port map( A => A(4), Z => n41);
   U41 : HS65_LH_IVX9 port map( A => A(16), Z => n34);
   U42 : HS65_LH_IVX9 port map( A => A(24), Z => n29);
   U43 : HS65_LH_IVX9 port map( A => A(30), Z => n26);
   U44 : HS65_LH_IVX9 port map( A => A(10), Z => n36);
   U45 : HS65_LH_NOR4ABX2 port map( A => n43, B => n44, C => n45, D => n46, Z 
                           => EQ_port);
   U46 : HS65_LH_NAND4X4 port map( A => n47, B => n48, C => n49, D => n50, Z =>
                           n46);
   U47 : HS65_LH_NAND4ABX3 port map( A => n51, B => n35, C => n52, D => n53, Z 
                           => n45);
   U48 : HS65_LH_NOR4ABX2 port map( A => n55, B => n56, C => n57, D => n58, Z 
                           => n44);
   U49 : HS65_LH_NAND4ABX3 port map( A => n59, B => n60, C => n61, D => n62, Z 
                           => n58);
   U50 : HS65_LH_AOI22X1 port map( A => n42, B => n63, C => n63, D => B(1), Z 
                           => n59);
   U51 : HS65_LH_NAND2AX4 port map( A => B(0), B => A(0), Z => n63);
   U52 : HS65_LH_NAND4ABX3 port map( A => n64, B => n27, C => n65, D => n66, Z 
                           => n57);
   U53 : HS65_LH_NOR4ABX2 port map( A => n68, B => n69, C => n70, D => n71, Z 
                           => n56);
   U54 : HS65_LH_AND4X3 port map( A => n72, B => n73, C => n74, D => n75, Z => 
                           n55);
   U55 : HS65_LH_NOR4ABX2 port map( A => n76, B => n77, C => n78, D => LT_port,
                           Z => n43);
   U56 : HS65_LH_OAI22X1 port map( A => A(31), B => n19, C => n24, D => n79, Z 
                           => LT_port);
   U57 : HS65_LH_AOI32X3 port map( A => n62, B => n25, C => n80, D => B(30), E 
                           => n26, Z => n79);
   U58 : HS65_LH_OAI212X3 port map( A => A(28), B => n17, C => A(29), D => n18,
                           E => n81, Z => n80);
   U59 : HS65_LH_NAND3X2 port map( A => n61, B => n67, C => n82, Z => n81);
   U60 : HS65_LH_OAI12X2 port map( A => A(27), B => n16, C => n83, Z => n82);
   U61 : HS65_LH_AOI32X3 port map( A => n66, B => n65, C => n84, D => B(26), E 
                           => n22, Z => n83);
   U62 : HS65_LH_OAI12X2 port map( A => A(25), B => n15, C => n85, Z => n84);
   U63 : HS65_LH_AOI32X3 port map( A => n28, B => n72, C => n86, D => B(24), E 
                           => n29, Z => n85);
   U64 : HS65_LH_OAI12X2 port map( A => A(23), B => n14, C => n87, Z => n86);
   U65 : HS65_LH_AOI32X3 port map( A => n73, B => n75, C => n88, D => B(22), E 
                           => n30, Z => n87);
   U66 : HS65_LH_OAI212X3 port map( A => A(20), B => n12, C => A(21), D => n13,
                           E => n89, Z => n88);
   U67 : HS65_LH_NAND3X2 port map( A => n74, B => n68, C => n90, Z => n89);
   U68 : HS65_LH_OAI12X2 port map( A => A(19), B => n11, C => n91, Z => n90);
   U69 : HS65_LH_AOI32X3 port map( A => n31, B => n69, C => n92, D => B(18), E 
                           => n32, Z => n91);
   U70 : HS65_LH_OAI12X2 port map( A => A(17), B => n10, C => n93, Z => n92);
   U71 : HS65_LH_AOI32X3 port map( A => n33, B => n49, C => n94, D => B(16), E 
                           => n34, Z => n93);
   U72 : HS65_LH_OAI12X2 port map( A => A(15), B => n9, C => n95, Z => n94);
   U73 : HS65_LH_AOI32X3 port map( A => n50, B => n48, C => n96, D => B(14), E 
                           => n21, Z => n95);
   U74 : HS65_LH_OAI212X3 port map( A => A(12), B => n7, C => A(13), D => n8, E
                           => n97, Z => n96);
   U75 : HS65_LH_NAND3X2 port map( A => n47, B => n54, C => n98, Z => n97);
   U76 : HS65_LH_OAI12X2 port map( A => A(11), B => n6, C => n99, Z => n98);
   U77 : HS65_LH_AOI32X3 port map( A => n53, B => n52, C => n100, D => B(10), E
                           => n36, Z => n99);
   U78 : HS65_LH_OAI12X2 port map( A => A(9), B => n5, C => n101, Z => n100);
   U79 : HS65_LH_AOI32X3 port map( A => n37, B => n102, C => n103, D => B(8), E
                           => n20, Z => n101);
   U80 : HS65_LH_OAI12X2 port map( A => A(7), B => n4, C => n104, Z => n103);
   U81 : HS65_LH_AOI32X3 port map( A => n105, B => n106, C => n107, D => B(6), 
                           E => n39, Z => n104);
   U82 : HS65_LH_OAI12X2 port map( A => A(5), B => n3, C => n108, Z => n107);
   U83 : HS65_LH_AOI32X3 port map( A => n40, B => n109, C => n110, D => B(4), E
                           => n41, Z => n108);
   U84 : HS65_LH_OAI212X3 port map( A => A(2), B => n1, C => A(3), D => n2, E 
                           => n111, Z => n110);
   U85 : HS65_LH_OAI212X3 port map( A => B(1), B => n112, C => n113, D => n42, 
                           E => n114, Z => n111);
   U86 : HS65_LH_AND2X4 port map( A => n113, B => n42, Z => n112);
   U87 : HS65_LH_NOR2AX3 port map( A => B(0), B => A(0), Z => n113);
   U88 : HS65_LH_NOR2X2 port map( A => n20, B => B(8), Z => n51);
   U89 : HS65_LH_NAND2X2 port map( A => A(9), B => n5, Z => n52);
   U90 : HS65_LH_NAND2AX4 port map( A => B(10), B => A(10), Z => n53);
   U91 : HS65_LH_NAND2X2 port map( A => A(11), B => n6, Z => n54);
   U92 : HS65_LH_NAND2X2 port map( A => A(12), B => n7, Z => n47);
   U93 : HS65_LH_NAND2X2 port map( A => A(13), B => n8, Z => n48);
   U94 : HS65_LH_NAND2X2 port map( A => A(15), B => n9, Z => n49);
   U95 : HS65_LH_NOR2X2 port map( A => n34, B => B(16), Z => n71);
   U96 : HS65_LH_NAND2X2 port map( A => A(17), B => n10, Z => n69);
   U97 : HS65_LH_NOR2X2 port map( A => B(18), B => n32, Z => n70);
   U98 : HS65_LH_NAND2X2 port map( A => A(19), B => n11, Z => n68);
   U99 : HS65_LH_NAND2X2 port map( A => A(20), B => n12, Z => n74);
   U100 : HS65_LH_NAND2X2 port map( A => A(21), B => n13, Z => n75);
   U101 : HS65_LH_NAND2AX4 port map( A => B(22), B => A(22), Z => n73);
   U102 : HS65_LH_NAND2X2 port map( A => A(23), B => n14, Z => n72);
   U103 : HS65_LH_NOR2X2 port map( A => n29, B => B(24), Z => n64);
   U104 : HS65_LH_NAND2X2 port map( A => A(25), B => n15, Z => n65);
   U105 : HS65_LH_NAND2X2 port map( A => A(27), B => n16, Z => n67);
   U106 : HS65_LH_NAND2X2 port map( A => A(28), B => n17, Z => n61);
   U107 : HS65_LH_NOR2X2 port map( A => n26, B => B(30), Z => n60);
   U108 : HS65_LH_NAND2X2 port map( A => A(29), B => n18, Z => n62);
   U109 : HS65_LH_NAND4ABX3 port map( A => n115, B => n38, C => n106, D => n105
                           , Z => n78);
   U110 : HS65_LH_NAND2AX4 port map( A => B(6), B => A(6), Z => n105);
   U111 : HS65_LH_NAND2X2 port map( A => A(5), B => n3, Z => n106);
   U112 : HS65_LH_NAND2X2 port map( A => A(7), B => n4, Z => n102);
   U113 : HS65_LH_NOR2X2 port map( A => n41, B => B(4), Z => n115);
   U114 : HS65_LH_AND2X4 port map( A => n114, B => n109, Z => n77);
   U115 : HS65_LH_NAND2X2 port map( A => A(3), B => n2, Z => n109);
   U116 : HS65_LH_NAND2X2 port map( A => A(2), B => n1, Z => n114);
   U117 : HS65_LH_NAND2X2 port map( A => A(31), B => n19, Z => n76);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_sub_0;

architecture SYN_rpl of alu_DW01_sub_0 is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33 : 
      std_logic;

begin
   
   U2_31 : HS65_LHS_XOR3X2 port map( A => A(31), B => n33, C => carry_31_port, 
                           Z => DIFF(31));
   U2_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => n32, CI => carry_30_port,
                           CO => carry_31_port, S0 => DIFF(30));
   U2_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => n30, CI => carry_28_port,
                           CO => carry_29_port, S0 => DIFF(28));
   U2_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => n29, CI => carry_27_port,
                           CO => carry_28_port, S0 => DIFF(27));
   U2_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => n27, CI => carry_25_port,
                           CO => carry_26_port, S0 => DIFF(25));
   U2_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => n26, CI => carry_24_port,
                           CO => carry_25_port, S0 => DIFF(24));
   U2_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => n24, CI => carry_22_port,
                           CO => carry_23_port, S0 => DIFF(22));
   U2_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => n23, CI => carry_21_port,
                           CO => carry_22_port, S0 => DIFF(21));
   U2_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => n21, CI => carry_19_port,
                           CO => carry_20_port, S0 => DIFF(19));
   U2_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => n20, CI => carry_18_port,
                           CO => carry_19_port, S0 => DIFF(18));
   U2_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => n18, CI => carry_16_port,
                           CO => carry_17_port, S0 => DIFF(16));
   U2_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => n17, CI => carry_15_port,
                           CO => carry_16_port, S0 => DIFF(15));
   U2_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => n15, CI => carry_13_port,
                           CO => carry_14_port, S0 => DIFF(13));
   U2_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => n14, CI => carry_12_port,
                           CO => carry_13_port, S0 => DIFF(12));
   U2_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => n12, CI => carry_10_port,
                           CO => carry_11_port, S0 => DIFF(10));
   U2_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => n11, CI => carry_9_port, CO
                           => carry_10_port, S0 => DIFF(9));
   U2_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => n9, CI => carry_7_port, CO 
                           => carry_8_port, S0 => DIFF(7));
   U2_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => n8, CI => carry_6_port, CO 
                           => carry_7_port, S0 => DIFF(6));
   U2_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => n6, CI => carry_4_port, CO 
                           => carry_5_port, S0 => DIFF(4));
   U2_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => n5, CI => carry_3_port, CO 
                           => carry_4_port, S0 => DIFF(3));
   U2_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => n3, CI => carry_1_port, CO 
                           => carry_2_port, S0 => DIFF(1));
   U2_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => n25, CI => carry_23_port,
                           CO => carry_24_port, S0 => DIFF(23));
   U2_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => n4, CI => carry_2_port, CO 
                           => carry_3_port, S0 => DIFF(2));
   U2_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => n31, CI => carry_29_port,
                           CO => carry_30_port, S0 => DIFF(29));
   U2_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => n28, CI => carry_26_port,
                           CO => carry_27_port, S0 => DIFF(26));
   U2_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => n22, CI => carry_20_port,
                           CO => carry_21_port, S0 => DIFF(20));
   U2_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => n19, CI => carry_17_port,
                           CO => carry_18_port, S0 => DIFF(17));
   U2_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => n13, CI => carry_11_port,
                           CO => carry_12_port, S0 => DIFF(11));
   U2_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => n7, CI => carry_5_port, CO 
                           => carry_6_port, S0 => DIFF(5));
   U2_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => n16, CI => carry_14_port,
                           CO => carry_15_port, S0 => DIFF(14));
   U2_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => n10, CI => carry_8_port, CO
                           => carry_9_port, S0 => DIFF(8));
   U1 : HS65_LH_IVX9 port map( A => B(8), Z => n10);
   U2 : HS65_LH_IVX9 port map( A => B(14), Z => n16);
   U3 : HS65_LH_IVX9 port map( A => B(5), Z => n7);
   U4 : HS65_LH_IVX9 port map( A => B(11), Z => n13);
   U5 : HS65_LH_IVX9 port map( A => B(17), Z => n19);
   U6 : HS65_LH_IVX9 port map( A => B(20), Z => n22);
   U7 : HS65_LH_IVX9 port map( A => B(26), Z => n28);
   U8 : HS65_LH_IVX9 port map( A => B(29), Z => n31);
   U9 : HS65_LH_IVX9 port map( A => B(2), Z => n4);
   U10 : HS65_LH_IVX9 port map( A => B(23), Z => n25);
   U11 : HS65_LH_IVX9 port map( A => B(0), Z => n2);
   U12 : HS65_LHS_XNOR2X6 port map( A => A(0), B => n2, Z => DIFF(0));
   U13 : HS65_LH_IVX9 port map( A => B(1), Z => n3);
   U14 : HS65_LH_NAND2X7 port map( A => n1, B => B(0), Z => carry_1_port);
   U15 : HS65_LH_IVX9 port map( A => A(0), Z => n1);
   U16 : HS65_LH_IVX9 port map( A => B(3), Z => n5);
   U17 : HS65_LH_IVX9 port map( A => B(4), Z => n6);
   U18 : HS65_LH_IVX9 port map( A => B(6), Z => n8);
   U19 : HS65_LH_IVX9 port map( A => B(7), Z => n9);
   U20 : HS65_LH_IVX9 port map( A => B(9), Z => n11);
   U21 : HS65_LH_IVX9 port map( A => B(10), Z => n12);
   U22 : HS65_LH_IVX9 port map( A => B(12), Z => n14);
   U23 : HS65_LH_IVX9 port map( A => B(13), Z => n15);
   U24 : HS65_LH_IVX9 port map( A => B(15), Z => n17);
   U25 : HS65_LH_IVX9 port map( A => B(16), Z => n18);
   U26 : HS65_LH_IVX9 port map( A => B(18), Z => n20);
   U27 : HS65_LH_IVX9 port map( A => B(19), Z => n21);
   U28 : HS65_LH_IVX9 port map( A => B(21), Z => n23);
   U29 : HS65_LH_IVX9 port map( A => B(22), Z => n24);
   U30 : HS65_LH_IVX9 port map( A => B(24), Z => n26);
   U31 : HS65_LH_IVX9 port map( A => B(25), Z => n27);
   U32 : HS65_LH_IVX9 port map( A => B(27), Z => n29);
   U33 : HS65_LH_IVX9 port map( A => B(28), Z => n30);
   U34 : HS65_LH_IVX9 port map( A => B(30), Z => n32);
   U35 : HS65_LH_IVX9 port map( A => B(31), Z => n33);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_cmp_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in 
         std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);

end alu_DW_cmp_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_cmp_0 is

   component HS65_LH_NAND2AX4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI312X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI112X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X2
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3AX3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X1
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA112X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI32X2
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328 : std_logic;

begin
   
   U157 : HS65_LH_IVX9 port map( A => n305, Z => n256);
   U158 : HS65_LH_OR2X9 port map( A => B(11), B => n241, Z => n327);
   U159 : HS65_LH_IVX9 port map( A => n316, Z => n266);
   U160 : HS65_LH_IVX9 port map( A => B(3), Z => n228);
   U161 : HS65_LH_IVX9 port map( A => B(4), Z => n229);
   U162 : HS65_LH_IVX9 port map( A => A(17), Z => n243);
   U163 : HS65_LH_IVX9 port map( A => A(11), Z => n241);
   U164 : HS65_LH_IVX9 port map( A => B(27), Z => n237);
   U165 : HS65_LH_IVX9 port map( A => B(2), Z => n227);
   U166 : HS65_LH_IVX9 port map( A => A(14), Z => n242);
   U167 : HS65_LH_IVX9 port map( A => A(8), Z => n240);
   U168 : HS65_LH_IVX9 port map( A => A(20), Z => n244);
   U169 : HS65_LH_IVX9 port map( A => A(5), Z => n239);
   U170 : HS65_LH_IVX9 port map( A => A(29), Z => n245);
   U171 : HS65_LH_IVX9 port map( A => n321, Z => n257);
   U172 : HS65_LH_IVX9 port map( A => n306, Z => n260);
   U173 : HS65_LH_IVX9 port map( A => n296, Z => n247);
   U174 : HS65_LH_OR2X9 port map( A => B(17), B => n243, Z => n281);
   U175 : HS65_LH_IVX9 port map( A => n279, Z => n252);
   U176 : HS65_LH_IVX9 port map( A => n297, Z => n246);
   U177 : HS65_LH_IVX9 port map( A => n284, Z => n250);
   U178 : HS65_LH_IVX9 port map( A => n320, Z => n254);
   U179 : HS65_LH_IVX9 port map( A => n308, Z => n263);
   U180 : HS65_LH_IVX9 port map( A => B(1), Z => n226);
   U181 : HS65_LH_IVX9 port map( A => B(23), Z => n233);
   U182 : HS65_LH_IVX9 port map( A => B(19), Z => n231);
   U183 : HS65_LH_IVX9 port map( A => B(26), Z => n236);
   U184 : HS65_LH_IVX9 port map( A => B(22), Z => n232);
   U185 : HS65_LH_IVX9 port map( A => B(18), Z => n230);
   U186 : HS65_LH_IVX9 port map( A => B(24), Z => n234);
   U187 : HS65_LH_IVX9 port map( A => B(30), Z => n238);
   U188 : HS65_LH_IVX9 port map( A => A(15), Z => n255);
   U189 : HS65_LH_IVX9 port map( A => A(7), Z => n264);
   U190 : HS65_LH_IVX9 port map( A => A(1), Z => n268);
   U191 : HS65_LH_IVX9 port map( A => B(25), Z => n235);
   U192 : HS65_LH_AND2X4 port map( A => A(3), B => n228, Z => n318);
   U193 : HS65_LH_IVX9 port map( A => A(9), Z => n262);
   U194 : HS65_LH_IVX9 port map( A => A(31), Z => n248);
   U195 : HS65_LH_IVX9 port map( A => A(21), Z => n251);
   U196 : HS65_LH_IVX9 port map( A => A(16), Z => n253);
   U197 : HS65_LH_IVX9 port map( A => A(13), Z => n258);
   U198 : HS65_LH_IVX9 port map( A => A(12), Z => n259);
   U199 : HS65_LH_IVX9 port map( A => A(28), Z => n249);
   U200 : HS65_LH_IVX9 port map( A => A(6), Z => n265);
   U201 : HS65_LH_IVX9 port map( A => A(10), Z => n261);
   U202 : HS65_LH_IVX9 port map( A => A(4), Z => n267);
   U203 : HS65_LH_OAI12X2 port map( A => n269, B => n270, C => n271, Z => 
                           GE_LT_GT_LE);
   U204 : HS65_LH_OAI32X2 port map( A => n272, B => n273, C => n274, D => n275,
                           E => n272, Z => n271);
   U205 : HS65_LH_AOI212X2 port map( A => n276, B => n277, C => n277, D => n252
                           , E => n278, Z => n274);
   U206 : HS65_LH_OA32X4 port map( A => n230, B => A(18), C => n280, D => A(19)
                           , E => n231, Z => n277);
   U207 : HS65_LH_AOI32X3 port map( A => n281, B => n253, C => B(16), D => 
                           B(17), E => n243, Z => n276);
   U208 : HS65_LH_AOI22X1 port map( A => n282, B => n283, C => n283, D => n250,
                           Z => n273);
   U209 : HS65_LH_OA32X4 port map( A => n232, B => A(22), C => n285, D => A(23)
                           , E => n233, Z => n283);
   U210 : HS65_LH_AOI32X3 port map( A => n286, B => n244, C => B(20), D => 
                           B(21), E => n251, Z => n282);
   U211 : HS65_LH_CBI4I1X3 port map( A => n247, B => n246, C => n287, D => n288
                           , Z => n272);
   U212 : HS65_LH_OAI212X3 port map( A => n289, B => n290, C => n291, D => n289
                           , E => n292, Z => n288);
   U213 : HS65_LH_OAI32X2 port map( A => n234, B => A(24), C => n293, D => 
                           A(25), E => n235, Z => n290);
   U214 : HS65_LH_OAI32X2 port map( A => n236, B => A(26), C => n294, D => 
                           A(27), E => n237, Z => n289);
   U215 : HS65_LH_AOI312X2 port map( A => n295, B => n249, C => B(28), D => 
                           B(29), E => n245, F => n296, Z => n287);
   U216 : HS65_LH_OAI32X2 port map( A => n238, B => A(30), C => n298, D => 
                           B(31), E => n248, Z => n296);
   U217 : HS65_LH_NAND3AX3 port map( A => n278, B => n279, C => n275, Z => n270
                           );
   U218 : HS65_LH_AND3X4 port map( A => n291, B => n292, C => n299, Z => n275);
   U219 : HS65_LH_AOI12X2 port map( A => A(24), B => n234, C => n293, Z => n299
                           );
   U220 : HS65_LH_NOR2AX3 port map( A => A(25), B => B(25), Z => n293);
   U221 : HS65_LH_OA112X4 port map( A => B(28), B => n249, C => n295, D => n297
                           , Z => n292);
   U222 : HS65_LH_AOI12X2 port map( A => n238, B => A(30), C => n298, Z => n297
                           );
   U223 : HS65_LH_AND2X4 port map( A => B(31), B => n248, Z => n298);
   U224 : HS65_LH_OR2X4 port map( A => B(29), B => n245, Z => n295);
   U225 : HS65_LH_AOI12X2 port map( A => n236, B => A(26), C => n294, Z => n291
                           );
   U226 : HS65_LH_AND2X4 port map( A => A(27), B => n237, Z => n294);
   U227 : HS65_LH_AOI12X2 port map( A => n230, B => A(18), C => n280, Z => n279
                           );
   U228 : HS65_LH_AND2X4 port map( A => A(19), B => n231, Z => n280);
   U229 : HS65_LH_OAI112X1 port map( A => B(20), B => n244, C => n286, D => 
                           n284, Z => n278);
   U230 : HS65_LH_AOI12X2 port map( A => n232, B => A(22), C => n285, Z => n284
                           );
   U231 : HS65_LH_AND2X4 port map( A => A(23), B => n233, Z => n285);
   U232 : HS65_LH_OR2X4 port map( A => B(21), B => n251, Z => n286);
   U233 : HS65_LH_OAI212X3 port map( A => n300, B => n301, C => n302, D => n300
                           , E => n303, Z => n269);
   U234 : HS65_LH_OA12X4 port map( A => n253, B => B(16), C => n281, Z => n303)
                           ;
   U235 : HS65_LH_NOR3X1 port map( A => n304, B => n305, C => n306, Z => n302);
   U236 : HS65_LH_OAI12X2 port map( A => B(8), B => n240, C => n307, Z => n304)
                           ;
   U237 : HS65_LH_CBI4I1X3 port map( A => n308, B => n309, C => n310, D => n311
                           , Z => n301);
   U238 : HS65_LH_NAND3AX3 port map( A => n309, B => n312, C => n313, Z => n311
                           );
   U239 : HS65_LH_AOI212X2 port map( A => n314, B => n315, C => A(4), D => n229
                           , E => n316, Z => n313);
   U240 : HS65_LH_AOI22X1 port map( A => B(1), B => n268, C => n317, D => B(0),
                           Z => n314);
   U241 : HS65_LH_AOI12X2 port map( A => A(1), B => n226, C => A(0), Z => n317)
                           ;
   U242 : HS65_LH_CBI4I1X3 port map( A => A(2), B => n227, C => n318, D => n315
                           , Z => n312);
   U243 : HS65_LH_OA32X4 port map( A => n227, B => A(2), C => n318, D => A(3), 
                           E => n228, Z => n315);
   U244 : HS65_LH_AOI312X2 port map( A => n266, B => n267, C => B(4), D => B(5)
                           , E => n239, F => n263, Z => n310);
   U245 : HS65_LH_NOR2X2 port map( A => n239, B => B(5), Z => n316);
   U246 : HS65_LH_OAI12X2 port map( A => B(6), B => n265, C => n319, Z => n309)
                           ;
   U247 : HS65_LH_AOI32X3 port map( A => B(6), B => n265, C => n319, D => n264,
                           E => B(7), Z => n308);
   U248 : HS65_LH_NAND2AX4 port map( A => B(7), B => A(7), Z => n319);
   U249 : HS65_LH_CBI4I1X3 port map( A => n320, B => n321, C => n322, D => n323
                           , Z => n300);
   U250 : HS65_LH_OAI212X3 port map( A => n324, B => n325, C => n260, D => n324
                           , E => n256, Z => n323);
   U251 : HS65_LH_OAI112X1 port map( A => B(12), B => n259, C => n326, D => 
                           n257, Z => n305);
   U252 : HS65_LH_OAI12X2 port map( A => B(10), B => n261, C => n327, Z => n306
                           );
   U253 : HS65_LH_AO32X4 port map( A => B(8), B => n240, C => n307, D => n262, 
                           E => B(9), Z => n325);
   U254 : HS65_LH_NAND2AX4 port map( A => B(9), B => A(9), Z => n307);
   U255 : HS65_LH_AO32X4 port map( A => B(10), B => n261, C => n327, D => n241,
                           E => B(11), Z => n324);
   U256 : HS65_LH_AOI312X2 port map( A => n326, B => n259, C => B(12), D => 
                           B(13), E => n258, F => n254, Z => n322);
   U257 : HS65_LH_OR2X4 port map( A => B(13), B => n258, Z => n326);
   U258 : HS65_LH_OAI12X2 port map( A => B(14), B => n242, C => n328, Z => n321
                           );
   U259 : HS65_LH_AOI32X3 port map( A => B(14), B => n242, C => n328, D => n255
                           , E => B(15), Z => n320);
   U260 : HS65_LH_NAND2AX4 port map( A => B(15), B => A(15), Z => n328);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu is

   port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 0);
         alu_o : out std_logic_vector (32 downto 0));

end alu;

architecture SYN_behavioral of alu is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO112X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI222X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I6X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI211X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component alu_DW_mult_uns_0
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component alu_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component alu_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW_cmp_0
      port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in
            std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal HI_LO_c_HI_31_port, HI_LO_c_HI_30_port, HI_LO_c_HI_29_port, 
      HI_LO_c_HI_28_port, HI_LO_c_HI_27_port, HI_LO_c_HI_26_port, 
      HI_LO_c_HI_25_port, HI_LO_c_HI_24_port, HI_LO_c_HI_23_port, 
      HI_LO_c_HI_22_port, HI_LO_c_HI_21_port, HI_LO_c_HI_20_port, 
      HI_LO_c_HI_19_port, HI_LO_c_HI_18_port, HI_LO_c_HI_17_port, 
      HI_LO_c_HI_16_port, HI_LO_c_HI_15_port, HI_LO_c_HI_14_port, 
      HI_LO_c_HI_13_port, HI_LO_c_HI_12_port, HI_LO_c_HI_11_port, 
      HI_LO_c_HI_10_port, HI_LO_c_HI_9_port, HI_LO_c_HI_8_port, 
      HI_LO_c_HI_7_port, HI_LO_c_HI_6_port, HI_LO_c_HI_5_port, 
      HI_LO_c_HI_4_port, HI_LO_c_HI_3_port, HI_LO_c_HI_2_port, 
      HI_LO_c_HI_1_port, HI_LO_c_HI_0_port, HI_LO_c_LO_31_port, 
      HI_LO_c_LO_30_port, HI_LO_c_LO_29_port, HI_LO_c_LO_28_port, 
      HI_LO_c_LO_27_port, HI_LO_c_LO_26_port, HI_LO_c_LO_25_port, 
      HI_LO_c_LO_24_port, HI_LO_c_LO_23_port, HI_LO_c_LO_22_port, 
      HI_LO_c_LO_21_port, HI_LO_c_LO_20_port, HI_LO_c_LO_19_port, 
      HI_LO_c_LO_18_port, HI_LO_c_LO_17_port, HI_LO_c_LO_16_port, 
      HI_LO_c_LO_15_port, HI_LO_c_LO_14_port, HI_LO_c_LO_13_port, 
      HI_LO_c_LO_12_port, HI_LO_c_LO_11_port, HI_LO_c_LO_10_port, 
      HI_LO_c_LO_9_port, HI_LO_c_LO_8_port, HI_LO_c_LO_7_port, 
      HI_LO_c_LO_6_port, HI_LO_c_LO_5_port, HI_LO_c_LO_4_port, 
      HI_LO_c_LO_3_port, HI_LO_c_LO_2_port, HI_LO_c_LO_1_port, 
      HI_LO_c_LO_0_port, N99, N100, N101, N102, N103, N104, N105, N106, N107, 
      N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, 
      N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, 
      N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, 
      N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, 
      N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, 
      N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, 
      N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, 
      N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, 
      N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, 
      N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N648, 
      N649, N714, N715, n1, n2, n3, n4, n5, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114_port, n115_port, n116_port, 
      n117_port, n118_port, n119_port, n120_port, n121_port, n122_port, 
      n123_port, n124_port, n125_port, n126_port, n127_port, n128_port, 
      n129_port, n130_port, n131_port, n132_port, n133_port, n134_port, 
      n135_port, n136_port, n137_port, n138_port, n139_port, n140_port, 
      n141_port, n142_port, n143_port, n144_port, n145_port, n146_port, 
      n147_port, n148_port, n149_port, n150_port, n151_port, n152_port, 
      n153_port, n154_port, n155_port, n156_port, n157_port, n158_port, 
      n159_port, n160_port, n161_port, n162_port, n163_port, n164_port, 
      n165_port, n166_port, n167_port, n168_port, n169_port, n170_port, 
      n171_port, n172_port, n173_port, n174_port, n175_port, n176_port, 
      n177_port, n178_port, n179_port, n180_port, n181_port, n182_port, 
      n183_port, n184_port, n185_port, n186_port, n187_port, n188_port, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204_port, n205_port, n206_port, 
      n207_port, n208_port, n209_port, n210_port, n211_port, n212_port, 
      n213_port, n214_port, n215_port, n216_port, n217_port, n218_port, 
      n219_port, n220_port, n221_port, n222_port, n223_port, n224_port, 
      n225_port, n226_port, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n300, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017 : std_logic;

begin
   
   n1 <= '1';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   HI_LO_c_reg_HI_31_inst : HS65_LH_DFPRQX9 port map( D => n516, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_31_port);
   HI_LO_c_reg_HI_30_inst : HS65_LH_DFPRQX9 port map( D => n515, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_30_port);
   HI_LO_c_reg_HI_29_inst : HS65_LH_DFPRQX9 port map( D => n514, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_29_port);
   HI_LO_c_reg_HI_28_inst : HS65_LH_DFPRQX9 port map( D => n513, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_28_port);
   HI_LO_c_reg_HI_27_inst : HS65_LH_DFPRQX9 port map( D => n512, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_27_port);
   HI_LO_c_reg_HI_26_inst : HS65_LH_DFPRQX9 port map( D => n511, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_26_port);
   HI_LO_c_reg_HI_25_inst : HS65_LH_DFPRQX9 port map( D => n510, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_25_port);
   HI_LO_c_reg_HI_24_inst : HS65_LH_DFPRQX9 port map( D => n509, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_24_port);
   HI_LO_c_reg_HI_23_inst : HS65_LH_DFPRQX9 port map( D => n508, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_23_port);
   HI_LO_c_reg_HI_22_inst : HS65_LH_DFPRQX9 port map( D => n507, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_22_port);
   HI_LO_c_reg_HI_21_inst : HS65_LH_DFPRQX9 port map( D => n506, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_21_port);
   HI_LO_c_reg_HI_20_inst : HS65_LH_DFPRQX9 port map( D => n505, CP => clk, RN 
                           => n538, Q => HI_LO_c_HI_20_port);
   HI_LO_c_reg_HI_19_inst : HS65_LH_DFPRQX9 port map( D => n504, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_19_port);
   HI_LO_c_reg_HI_18_inst : HS65_LH_DFPRQX9 port map( D => n503, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_18_port);
   HI_LO_c_reg_HI_17_inst : HS65_LH_DFPRQX9 port map( D => n502, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_17_port);
   HI_LO_c_reg_HI_16_inst : HS65_LH_DFPRQX9 port map( D => n501, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_16_port);
   HI_LO_c_reg_HI_15_inst : HS65_LH_DFPRQX9 port map( D => n500, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_15_port);
   HI_LO_c_reg_HI_14_inst : HS65_LH_DFPRQX9 port map( D => n499, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_14_port);
   HI_LO_c_reg_HI_13_inst : HS65_LH_DFPRQX9 port map( D => n498, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_13_port);
   HI_LO_c_reg_HI_12_inst : HS65_LH_DFPRQX9 port map( D => n497, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_12_port);
   HI_LO_c_reg_HI_11_inst : HS65_LH_DFPRQX9 port map( D => n496, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_11_port);
   HI_LO_c_reg_HI_10_inst : HS65_LH_DFPRQX9 port map( D => n495, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_10_port);
   HI_LO_c_reg_HI_9_inst : HS65_LH_DFPRQX9 port map( D => n494, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_9_port);
   HI_LO_c_reg_HI_8_inst : HS65_LH_DFPRQX9 port map( D => n493, CP => clk, RN 
                           => n539, Q => HI_LO_c_HI_8_port);
   HI_LO_c_reg_HI_7_inst : HS65_LH_DFPRQX9 port map( D => n492, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_7_port);
   HI_LO_c_reg_HI_6_inst : HS65_LH_DFPRQX9 port map( D => n491, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_6_port);
   HI_LO_c_reg_HI_5_inst : HS65_LH_DFPRQX9 port map( D => n490, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_5_port);
   HI_LO_c_reg_HI_4_inst : HS65_LH_DFPRQX9 port map( D => n489, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_4_port);
   HI_LO_c_reg_HI_3_inst : HS65_LH_DFPRQX9 port map( D => n488, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_3_port);
   HI_LO_c_reg_HI_2_inst : HS65_LH_DFPRQX9 port map( D => n487, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_2_port);
   HI_LO_c_reg_HI_1_inst : HS65_LH_DFPRQX9 port map( D => n486, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_1_port);
   HI_LO_c_reg_HI_0_inst : HS65_LH_DFPRQX9 port map( D => n485, CP => clk, RN 
                           => n540, Q => HI_LO_c_HI_0_port);
   HI_LO_c_reg_LO_31_inst : HS65_LH_DFPRQX9 port map( D => n484, CP => clk, RN 
                           => n540, Q => HI_LO_c_LO_31_port);
   HI_LO_c_reg_LO_30_inst : HS65_LH_DFPRQX9 port map( D => n483, CP => clk, RN 
                           => n540, Q => HI_LO_c_LO_30_port);
   HI_LO_c_reg_LO_29_inst : HS65_LH_DFPRQX9 port map( D => n482, CP => clk, RN 
                           => n540, Q => HI_LO_c_LO_29_port);
   HI_LO_c_reg_LO_28_inst : HS65_LH_DFPRQX9 port map( D => n481, CP => clk, RN 
                           => n540, Q => HI_LO_c_LO_28_port);
   HI_LO_c_reg_LO_27_inst : HS65_LH_DFPRQX9 port map( D => n480, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_27_port);
   HI_LO_c_reg_LO_26_inst : HS65_LH_DFPRQX9 port map( D => n479, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_26_port);
   HI_LO_c_reg_LO_25_inst : HS65_LH_DFPRQX9 port map( D => n478, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_25_port);
   HI_LO_c_reg_LO_24_inst : HS65_LH_DFPRQX9 port map( D => n477, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_24_port);
   HI_LO_c_reg_LO_23_inst : HS65_LH_DFPRQX9 port map( D => n476, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_23_port);
   HI_LO_c_reg_LO_22_inst : HS65_LH_DFPRQX9 port map( D => n475, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_22_port);
   HI_LO_c_reg_LO_21_inst : HS65_LH_DFPRQX9 port map( D => n474, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_21_port);
   HI_LO_c_reg_LO_20_inst : HS65_LH_DFPRQX9 port map( D => n473, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_20_port);
   HI_LO_c_reg_LO_19_inst : HS65_LH_DFPRQX9 port map( D => n472, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_19_port);
   HI_LO_c_reg_LO_18_inst : HS65_LH_DFPRQX9 port map( D => n471, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_18_port);
   HI_LO_c_reg_LO_17_inst : HS65_LH_DFPRQX9 port map( D => n470, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_17_port);
   HI_LO_c_reg_LO_16_inst : HS65_LH_DFPRQX9 port map( D => n469, CP => clk, RN 
                           => n541, Q => HI_LO_c_LO_16_port);
   HI_LO_c_reg_LO_15_inst : HS65_LH_DFPRQX9 port map( D => n468, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_15_port);
   HI_LO_c_reg_LO_14_inst : HS65_LH_DFPRQX9 port map( D => n467, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_14_port);
   HI_LO_c_reg_LO_13_inst : HS65_LH_DFPRQX9 port map( D => n466, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_13_port);
   HI_LO_c_reg_LO_12_inst : HS65_LH_DFPRQX9 port map( D => n465, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_12_port);
   HI_LO_c_reg_LO_11_inst : HS65_LH_DFPRQX9 port map( D => n464, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_11_port);
   HI_LO_c_reg_LO_10_inst : HS65_LH_DFPRQX9 port map( D => n463, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_10_port);
   HI_LO_c_reg_LO_9_inst : HS65_LH_DFPRQX9 port map( D => n462, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_9_port);
   HI_LO_c_reg_LO_8_inst : HS65_LH_DFPRQX9 port map( D => n461, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_8_port);
   HI_LO_c_reg_LO_7_inst : HS65_LH_DFPRQX9 port map( D => n460, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_7_port);
   HI_LO_c_reg_LO_6_inst : HS65_LH_DFPRQX9 port map( D => n459, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_6_port);
   HI_LO_c_reg_LO_5_inst : HS65_LH_DFPRQX9 port map( D => n458, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_5_port);
   HI_LO_c_reg_LO_4_inst : HS65_LH_DFPRQX9 port map( D => n457, CP => clk, RN 
                           => n542, Q => HI_LO_c_LO_4_port);
   HI_LO_c_reg_LO_3_inst : HS65_LH_DFPRQX9 port map( D => n456, CP => clk, RN 
                           => n543, Q => HI_LO_c_LO_3_port);
   HI_LO_c_reg_LO_2_inst : HS65_LH_DFPRQX9 port map( D => n455, CP => clk, RN 
                           => n543, Q => HI_LO_c_LO_2_port);
   HI_LO_c_reg_LO_1_inst : HS65_LH_DFPRQX9 port map( D => n454, CP => clk, RN 
                           => n543, Q => HI_LO_c_LO_1_port);
   HI_LO_c_reg_LO_0_inst : HS65_LH_DFPRQX9 port map( D => n453, CP => clk, RN 
                           => n543, Q => HI_LO_c_LO_0_port);
   lt_136 : alu_DW_cmp_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           alu_i(44), A(1) => alu_i(43), A(0) => alu_i(42), 
                           B(31) => alu_i(41), B(30) => n524, B(29) => n523, 
                           B(28) => alu_i(38), B(27) => alu_i(37), B(26) => 
                           n520, B(25) => n519, B(24) => n518, B(23) => n517, 
                           B(22) => n300, B(21) => n90, B(20) => alu_i(30), 
                           B(19) => n88, B(18) => n87, B(17) => n86, B(16) => 
                           n85, B(15) => n84, B(14) => n83, B(13) => n82, B(12)
                           => n81, B(11) => alu_i(21), B(10) => n79, B(9) => 
                           n78, B(8) => n77, B(7) => n76, B(6) => n75, B(5) => 
                           n74, B(4) => alu_i(14), B(3) => alu_i(13), B(2) => 
                           alu_i(12), B(1) => n70, B(0) => n69, TC => n1, GE_LT
                           => n1, GE_GT_EQ => n2, GE_LT_GT_LE => N648, EQ_NE =>
                           n_1012);
   sub_68 : alu_DW01_sub_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           alu_i(44), A(1) => alu_i(43), A(0) => alu_i(42), 
                           B(31) => alu_i(41), B(30) => n524, B(29) => n523, 
                           B(28) => alu_i(38), B(27) => alu_i(37), B(26) => 
                           n520, B(25) => n519, B(24) => n518, B(23) => n517, 
                           B(22) => n300, B(21) => n90, B(20) => alu_i(30), 
                           B(19) => n88, B(18) => n87, B(17) => n86, B(16) => 
                           n85, B(15) => n84, B(14) => n83, B(13) => n82, B(12)
                           => n81, B(11) => alu_i(21), B(10) => n79, B(9) => 
                           n78, B(8) => n77, B(7) => n76, B(6) => n75, B(5) => 
                           n74, B(4) => alu_i(14), B(3) => alu_i(13), B(2) => 
                           alu_i(12), B(1) => n70, B(0) => n69, CI => n3, 
                           DIFF(31) => N162, DIFF(30) => N161, DIFF(29) => N160
                           , DIFF(28) => N159, DIFF(27) => N158, DIFF(26) => 
                           N157, DIFF(25) => N156, DIFF(24) => N155, DIFF(23) 
                           => N154, DIFF(22) => N153, DIFF(21) => N152, 
                           DIFF(20) => N151, DIFF(19) => N150, DIFF(18) => N149
                           , DIFF(17) => N148, DIFF(16) => N147, DIFF(15) => 
                           N146, DIFF(14) => N145, DIFF(13) => N144, DIFF(12) 
                           => N143, DIFF(11) => N142, DIFF(10) => N141, DIFF(9)
                           => N140, DIFF(8) => N139, DIFF(7) => N138, DIFF(6) 
                           => N137, DIFF(5) => N136, DIFF(4) => N135, DIFF(3) 
                           => N134, DIFF(2) => N133, DIFF(1) => N132, DIFF(0) 
                           => N131, CO => n_1013);
   r325 : alu_DW01_cmp6_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           alu_i(44), A(1) => alu_i(43), A(0) => alu_i(42), 
                           B(31) => alu_i(41), B(30) => n524, B(29) => n523, 
                           B(28) => alu_i(38), B(27) => alu_i(37), B(26) => 
                           n520, B(25) => n519, B(24) => n518, B(23) => n517, 
                           B(22) => n300, B(21) => n90, B(20) => alu_i(30), 
                           B(19) => n88, B(18) => n87, B(17) => n86, B(16) => 
                           n85, B(15) => n84, B(14) => n83, B(13) => n82, B(12)
                           => n81, B(11) => alu_i(21), B(10) => n79, B(9) => 
                           n78, B(8) => n77, B(7) => n76, B(6) => n75, B(5) => 
                           n74, B(4) => alu_i(14), B(3) => alu_i(13), B(2) => 
                           alu_i(12), B(1) => n70, B(0) => n69, TC => n4, LT =>
                           N649, GT => n_1014, EQ => N714, LE => n_1015, GE => 
                           n_1016, NE => N715);
   r321 : alu_DW01_add_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => alu_i(71), A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => alu_i(68), A(25) => alu_i(67), 
                           A(24) => alu_i(66), A(23) => alu_i(65), A(22) => 
                           alu_i(64), A(21) => alu_i(63), A(20) => alu_i(62), 
                           A(19) => alu_i(61), A(18) => alu_i(60), A(17) => 
                           alu_i(59), A(16) => alu_i(58), A(15) => alu_i(57), 
                           A(14) => alu_i(56), A(13) => alu_i(55), A(12) => 
                           alu_i(54), A(11) => alu_i(53), A(10) => alu_i(52), 
                           A(9) => alu_i(51), A(8) => alu_i(50), A(7) => 
                           alu_i(49), A(6) => alu_i(48), A(5) => alu_i(47), 
                           A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           alu_i(44), A(1) => alu_i(43), A(0) => alu_i(42), 
                           B(31) => alu_i(41), B(30) => n524, B(29) => n523, 
                           B(28) => alu_i(38), B(27) => alu_i(37), B(26) => 
                           n520, B(25) => n519, B(24) => n518, B(23) => n517, 
                           B(22) => n300, B(21) => n90, B(20) => alu_i(30), 
                           B(19) => n88, B(18) => n87, B(17) => n86, B(16) => 
                           n85, B(15) => n84, B(14) => n83, B(13) => n82, B(12)
                           => n81, B(11) => alu_i(21), B(10) => n79, B(9) => 
                           n78, B(8) => n77, B(7) => n76, B(6) => n75, B(5) => 
                           n74, B(4) => alu_i(14), B(3) => alu_i(13), B(2) => 
                           alu_i(12), B(1) => n70, B(0) => n69, CI => n5, 
                           SUM(31) => N130, SUM(30) => N129, SUM(29) => N128, 
                           SUM(28) => N127, SUM(27) => N126, SUM(26) => N125, 
                           SUM(25) => N124, SUM(24) => N123, SUM(23) => N122, 
                           SUM(22) => N121, SUM(21) => N120, SUM(20) => N119, 
                           SUM(19) => N118, SUM(18) => N117, SUM(17) => N116, 
                           SUM(16) => N115, SUM(15) => N114, SUM(14) => N113, 
                           SUM(13) => N112, SUM(12) => N111, SUM(11) => N110, 
                           SUM(10) => N109, SUM(9) => N108, SUM(8) => N107, 
                           SUM(7) => N106, SUM(6) => N105, SUM(5) => N104, 
                           SUM(4) => N103, SUM(3) => N102, SUM(2) => N101, 
                           SUM(1) => N100, SUM(0) => N99, CO => n_1017);
   mult_71 : alu_DW_mult_uns_0 port map( a(31) => alu_i(73), a(30) => alu_i(72)
                           , a(29) => alu_i(71), a(28) => alu_i(70), a(27) => 
                           alu_i(69), a(26) => alu_i(68), a(25) => alu_i(67), 
                           a(24) => alu_i(66), a(23) => alu_i(65), a(22) => 
                           alu_i(64), a(21) => alu_i(63), a(20) => alu_i(62), 
                           a(19) => alu_i(61), a(18) => alu_i(60), a(17) => 
                           alu_i(59), a(16) => alu_i(58), a(15) => alu_i(57), 
                           a(14) => alu_i(56), a(13) => alu_i(55), a(12) => 
                           alu_i(54), a(11) => alu_i(53), a(10) => alu_i(52), 
                           a(9) => alu_i(51), a(8) => alu_i(50), a(7) => 
                           alu_i(49), a(6) => alu_i(48), a(5) => alu_i(47), 
                           a(4) => alu_i(46), a(3) => alu_i(45), a(2) => 
                           alu_i(44), a(1) => alu_i(43), a(0) => alu_i(42), 
                           b(31) => alu_i(41), b(30) => n524, b(29) => n523, 
                           b(28) => alu_i(38), b(27) => alu_i(37), b(26) => 
                           n520, b(25) => n519, b(24) => n518, b(23) => n517, 
                           b(22) => n300, b(21) => n90, b(20) => alu_i(30), 
                           b(19) => n88, b(18) => n87, b(17) => n86, b(16) => 
                           n85, b(15) => n84, b(14) => n83, b(13) => n82, b(12)
                           => n81, b(11) => alu_i(21), b(10) => n79, b(9) => 
                           n78, b(8) => n77, b(7) => n76, b(6) => n75, b(5) => 
                           n74, b(4) => alu_i(14), b(3) => alu_i(13), b(2) => 
                           alu_i(12), b(1) => n70, b(0) => n69, product(63) => 
                           N226, product(62) => N225, product(61) => N224, 
                           product(60) => N223, product(59) => N222, 
                           product(58) => N221, product(57) => N220, 
                           product(56) => N219, product(55) => N218, 
                           product(54) => N217, product(53) => N216, 
                           product(52) => N215, product(51) => N214, 
                           product(50) => N213, product(49) => N212, 
                           product(48) => N211, product(47) => N210, 
                           product(46) => N209, product(45) => N208, 
                           product(44) => N207, product(43) => N206, 
                           product(42) => N205, product(41) => N204, 
                           product(40) => N203, product(39) => N202, 
                           product(38) => N201, product(37) => N200, 
                           product(36) => N199, product(35) => N198, 
                           product(34) => N197, product(33) => N196, 
                           product(32) => N195, product(31) => N194, 
                           product(30) => N193, product(29) => N192, 
                           product(28) => N191, product(27) => N190, 
                           product(26) => N189, product(25) => N188, 
                           product(24) => N187, product(23) => N186, 
                           product(22) => N185, product(21) => N184, 
                           product(20) => N183, product(19) => N182, 
                           product(18) => N181, product(17) => N180, 
                           product(16) => N179, product(15) => N178, 
                           product(14) => N177, product(13) => N176, 
                           product(12) => N175, product(11) => N174, 
                           product(10) => N173, product(9) => N172, product(8) 
                           => N171, product(7) => N170, product(6) => N169, 
                           product(5) => N168, product(4) => N167, product(3) 
                           => N166, product(2) => N165, product(1) => N164, 
                           product(0) => N163);
   U3 : HS65_LH_NOR4ABX2 port map( A => n92, B => n93, C => n94, D => n95, Z =>
                           n91);
   U4 : HS65_LH_NOR2X6 port map( A => n98, B => alu_i(4), Z => n284);
   U5 : HS65_LH_BFX9 port map( A => alu_i(19), Z => n78);
   U6 : HS65_LH_BFX9 port map( A => alu_i(16), Z => n75);
   U7 : HS65_LH_BFX9 port map( A => alu_i(24), Z => n83);
   U13 : HS65_LH_BFX9 port map( A => alu_i(20), Z => n79);
   U14 : HS65_LH_BFX9 port map( A => alu_i(18), Z => n77);
   U15 : HS65_LH_BFX9 port map( A => alu_i(17), Z => n76);
   U16 : HS65_LH_BFX9 port map( A => alu_i(25), Z => n84);
   U17 : HS65_LH_BFX9 port map( A => alu_i(15), Z => n74);
   U18 : HS65_LH_BFX9 port map( A => alu_i(23), Z => n82);
   U19 : HS65_LH_BFX9 port map( A => alu_i(22), Z => n81);
   U20 : HS65_LH_BFX9 port map( A => alu_i(35), Z => n519);
   U21 : HS65_LH_BFX9 port map( A => alu_i(26), Z => n85);
   U22 : HS65_LH_BFX9 port map( A => alu_i(36), Z => n520);
   U23 : HS65_LH_BFX9 port map( A => alu_i(27), Z => n86);
   U24 : HS65_LH_BFX9 port map( A => alu_i(11), Z => n70);
   U25 : HS65_LH_BFX9 port map( A => alu_i(28), Z => n87);
   U26 : HS65_LH_BFX9 port map( A => alu_i(31), Z => n90);
   U27 : HS65_LH_BFX9 port map( A => alu_i(39), Z => n523);
   U28 : HS65_LH_BFX9 port map( A => alu_i(32), Z => n300);
   U29 : HS65_LH_BFX9 port map( A => alu_i(34), Z => n518);
   U30 : HS65_LH_BFX9 port map( A => alu_i(40), Z => n524);
   U31 : HS65_LH_BFX9 port map( A => alu_i(29), Z => n88);
   U32 : HS65_LH_BFX9 port map( A => alu_i(33), Z => n517);
   U33 : HS65_LH_OR2X9 port map( A => alu_i(2), B => alu_i(3), Z => n6);
   U34 : HS65_LH_IVX9 port map( A => n61, Z => n60);
   U35 : HS65_LH_IVX9 port map( A => n62, Z => n59);
   U36 : HS65_LH_IVX9 port map( A => n62, Z => n58);
   U37 : HS65_LH_IVX9 port map( A => n62, Z => n57);
   U38 : HS65_LH_IVX9 port map( A => n98, Z => n581);
   U39 : HS65_LH_IVX9 port map( A => n176_port, Z => n580);
   U40 : HS65_LH_IVX9 port map( A => n281, Z => n582);
   U41 : HS65_LH_IVX9 port map( A => n56, Z => n55);
   U42 : HS65_LH_IVX9 port map( A => n42, Z => n41);
   U43 : HS65_LH_BFX9 port map( A => n68, Z => n61);
   U44 : HS65_LH_BFX9 port map( A => n68, Z => n62);
   U45 : HS65_LH_BFX9 port map( A => n586, Z => n15);
   U46 : HS65_LH_BFX9 port map( A => n586, Z => n14);
   U47 : HS65_LH_BFX9 port map( A => n585, Z => n11);
   U48 : HS65_LH_BFX9 port map( A => n585, Z => n12);
   U49 : HS65_LH_BFX9 port map( A => n67, Z => n65);
   U50 : HS65_LH_BFX9 port map( A => n67, Z => n64);
   U51 : HS65_LH_BFX9 port map( A => n68, Z => n63);
   U52 : HS65_LH_BFX9 port map( A => n586, Z => n16);
   U53 : HS65_LH_BFX9 port map( A => n585, Z => n13);
   U54 : HS65_LH_BFX9 port map( A => n67, Z => n66);
   U55 : HS65_LH_IVX9 port map( A => n101_port, Z => n585);
   U56 : HS65_LH_IVX9 port map( A => n100_port, Z => n586);
   U57 : HS65_LH_NOR2X6 port map( A => n96, B => n189_port, Z => n279);
   U58 : HS65_LH_AOI222X2 port map( A => n275, B => n276, C => n277, D => n278,
                           E => n279, F => n214_port, Z => n274);
   U59 : HS65_LH_NAND2X7 port map( A => n442, B => n435, Z => n98);
   U60 : HS65_LH_IVX9 port map( A => n96, Z => n584);
   U61 : HS65_LH_NOR2X6 port map( A => n189_port, B => n98, Z => n115_port);
   U62 : HS65_LH_IVX9 port map( A => n208_port, Z => n579);
   U63 : HS65_LH_IVX9 port map( A => n186_port, Z => n583);
   U64 : HS65_LH_NAND2X7 port map( A => n195_port, B => n581, Z => n176_port);
   U65 : HS65_LH_NAND2X7 port map( A => n584, B => n195_port, Z => n281);
   U66 : HS65_LH_OAI211X5 port map( A => n39, B => n208_port, C => n101_port, D
                           => n40, Z => n207_port);
   U67 : HS65_LH_NOR3X4 port map( A => n48, B => n45, C => n106_port, Z => n92)
                           ;
   U68 : HS65_LH_IVX9 port map( A => n189_port, Z => n591);
   U69 : HS65_LH_IVX9 port map( A => n237, Z => n576);
   U70 : HS65_LH_AND2X4 port map( A => n275, B => n17, Z => n368);
   U71 : HS65_LH_AND2X4 port map( A => n117_port, B => n17, Z => n397);
   U72 : HS65_LH_IVX9 port map( A => n54, Z => n56);
   U73 : HS65_LH_IVX9 port map( A => n40, Z => n42);
   U74 : HS65_LH_BFX9 port map( A => n43, Z => n44);
   U75 : HS65_LH_BFX9 port map( A => n91, Z => n68);
   U76 : HS65_LH_BFX9 port map( A => n91, Z => n67);
   U77 : HS65_LH_BFX9 port map( A => n50, Z => n52);
   U78 : HS65_LH_BFX9 port map( A => n50, Z => n51);
   U79 : HS65_LH_IVX9 port map( A => n39, Z => n37);
   U80 : HS65_LH_BFX9 port map( A => n577, Z => n10);
   U81 : HS65_LH_BFX9 port map( A => n30, Z => n32);
   U82 : HS65_LH_BFX9 port map( A => n577, Z => n9);
   U83 : HS65_LH_BFX9 port map( A => n43, Z => n45);
   U84 : HS65_LH_BFX9 port map( A => n30, Z => n33);
   U85 : HS65_LH_BFX9 port map( A => n31, Z => n34);
   U86 : HS65_LH_IVX9 port map( A => n39, Z => n38);
   U87 : HS65_LH_BFX9 port map( A => n19, Z => n21);
   U88 : HS65_LH_BFX9 port map( A => n19, Z => n23);
   U89 : HS65_LH_BFX9 port map( A => n19, Z => n22);
   U90 : HS65_LH_BFX9 port map( A => n20, Z => n24);
   U91 : HS65_LH_IVX9 port map( A => n317, Z => n572);
   U92 : HS65_LH_BFX9 port map( A => n50, Z => n53);
   U93 : HS65_LH_IVX9 port map( A => n144_port, Z => n569);
   U94 : HS65_LH_IVX9 port map( A => n130_port, Z => n571);
   U95 : HS65_LH_IVX9 port map( A => n212_port, Z => n570);
   U96 : HS65_LH_BFX9 port map( A => n20, Z => n25);
   U97 : HS65_LH_BFX9 port map( A => n31, Z => n35);
   U98 : HS65_LH_NAND4ABX3 port map( A => n42, B => n53, C => n578, D => n10, Z
                           => n94);
   U99 : HS65_LH_NAND3X5 port map( A => n96, B => n55, C => n98, Z => n95);
   U100 : HS65_LH_NOR4ABX2 port map( A => n100_port, B => n101_port, C => 
                           n102_port, D => n103_port, Z => n93);
   U101 : HS65_LH_IVX9 port map( A => n180_port, Z => n577);
   U102 : HS65_LH_AOI222X2 port map( A => n32, B => n70, C => n27, D => n69, E 
                           => n196_port, F => alu_i(12), Z => n237);
   U103 : HS65_LH_NOR2X6 port map( A => n592, B => n96, Z => n275);
   U104 : HS65_LH_NAND2X7 port map( A => n436, B => n442, Z => n96);
   U105 : HS65_LH_AOI222X2 port map( A => n284, B => n387, C => n277, D => n314
                           , E => n279, F => n317, Z => n386);
   U106 : HS65_LH_AOI222X2 port map( A => n284, B => n360, C => n277, D => n302
                           , E => n279, F => n306, Z => n380);
   U107 : HS65_LH_AOI222X2 port map( A => n284, B => n239, C => n277, D => n336
                           , E => n279, F => n292, Z => n373);
   U108 : HS65_LH_AOI222X2 port map( A => n284, B => n566, C => n277, D => n326
                           , E => n279, F => n278, Z => n366);
   U109 : HS65_LH_IVX9 port map( A => n190_port, Z => n566);
   U110 : HS65_LH_AOI222X2 port map( A => n284, B => n174_port, C => n277, D =>
                           n316, E => n279, F => n266, Z => n349);
   U111 : HS65_LH_AOI222X2 port map( A => n275, B => n165_port, C => n279, D =>
                           n254, E => n284, F => n166_port, Z => n343);
   U112 : HS65_LH_AOI222X2 port map( A => n275, B => n153_port, C => n279, D =>
                           n229, E => n284, F => n155_port, Z => n333);
   U113 : HS65_LH_AOI222X2 port map( A => n275, B => n141_port, C => n279, D =>
                           n212_port, E => n284, F => n143_port, Z => n323);
   U114 : HS65_LH_AOI222X2 port map( A => n275, B => n129_port, C => n279, D =>
                           n268, E => n284, F => n131_port, Z => n312);
   U115 : HS65_LH_AOI222X2 port map( A => n275, B => n112_port, C => n279, D =>
                           n256, E => n284, F => n116_port, Z => n298);
   U116 : HS65_LH_AOI222X2 port map( A => n275, B => n290, C => n279, D => n231
                           , E => n284, F => n291, Z => n289);
   U117 : HS65_LH_AOI212X4 port map( A => alu_i(53), B => n180_port, C => n56, 
                           D => n529, E => n42, Z => n421);
   U118 : HS65_LH_AOI212X4 port map( A => alu_i(62), B => n180_port, C => n56, 
                           D => n532, E => n42, Z => n350);
   U119 : HS65_LH_NAND2X7 port map( A => n301, B => n592, Z => n189_port);
   U120 : HS65_LH_OAI212X5 port map( A => n574, B => n189_port, C => n190_port,
                           D => n592, E => n191_port, Z => n183_port);
   U121 : HS65_LH_IVX9 port map( A => n140_port, Z => n574);
   U122 : HS65_LH_AOI222X2 port map( A => n192_port, B => n145_port, C => 
                           n193_port, D => n194_port, E => n195_port, F => 
                           n142_port, Z => n191_port);
   U123 : HS65_LH_MX41X7 port map( D0 => alu_i(13), S0 => n37, D1 => alu_i(14),
                           S1 => n33, D2 => n74, S2 => n28, D3 => n75, S3 => 
                           n23, Z => n194_port);
   U124 : HS65_LH_OAI212X5 port map( A => n568, B => n189_port, C => n264, D =>
                           n592, E => n265, Z => n259);
   U125 : HS65_LH_IVX9 port map( A => n269, Z => n568);
   U126 : HS65_LH_AOI222X2 port map( A => n192_port, B => n266, C => n193_port,
                           D => n267, E => n195_port, F => n268, Z => n265);
   U127 : HS65_LH_MX41X7 port map( D0 => alu_i(38), S0 => n36, D1 => alu_i(37),
                           S1 => n32, D2 => n520, S2 => n27, D3 => n519, S3 => 
                           n21, Z => n267);
   U128 : HS65_LH_OAI212X5 port map( A => n236, B => n71, C => n237, D => 
                           n186_port, E => n238, Z => n235);
   U129 : HS65_LH_CBI4I1X5 port map( A => n56, B => n71, C => n42, D => 
                           alu_i(44), Z => n238);
   U130 : HS65_LH_AOI212X4 port map( A => alu_i(44), B => n180_port, C => n56, 
                           D => n526, E => n42, Z => n236);
   U131 : HS65_LH_NOR2X6 port map( A => n594, B => n593, Z => n374);
   U132 : HS65_LH_OAI212X5 port map( A => alu_i(71), B => n55, C => n9, D => 
                           n535, E => n41, Z => n248);
   U133 : HS65_LH_NOR2X6 port map( A => n592, B => n98, Z => n117_port);
   U134 : HS65_LH_OAI212X5 port map( A => alu_i(56), B => n54, C => n10, D => 
                           n530, E => n123_port, Z => n403);
   U135 : HS65_LH_OAI212X5 port map( A => alu_i(59), B => n54, C => n10, D => 
                           n531, E => n40, Z => n381);
   U136 : HS65_LH_OAI212X5 port map( A => alu_i(47), B => n55, C => n9, D => 
                           n527, E => n41, Z => n167_port);
   U137 : HS65_LH_OAI212X5 port map( A => alu_i(50), B => n55, C => n9, D => 
                           n528, E => n41, Z => n134_port);
   U138 : HS65_LH_OAI212X5 port map( A => alu_i(65), B => n55, C => n9, D => 
                           n533, E => n41, Z => n328);
   U139 : HS65_LH_OAI212X5 port map( A => alu_i(68), B => n55, C => n9, D => 
                           n534, E => n41, Z => n293);
   U140 : HS65_LH_AOI32X5 port map( A => n178_port, B => n593, C => n275, D => 
                           alu_i(62), E => n352, Z => n351);
   U141 : HS65_LH_OAI21X3 port map( A => alu_i(30), B => n54, C => n40, Z => 
                           n352);
   U142 : HS65_LH_AND2X4 port map( A => n192_port, B => n584, Z => n277);
   U143 : HS65_LH_NOR2X6 port map( A => n588, B => n590, Z => n435);
   U144 : HS65_LH_AOI32X5 port map( A => n283, B => n593, C => n117_port, D => 
                           alu_i(53), E => n423, Z => n422);
   U145 : HS65_LH_OAI21X3 port map( A => alu_i(21), B => n54, C => n123_port, Z
                           => n423);
   U146 : HS65_LH_NAND2X7 port map( A => n193_port, B => n581, Z => n208_port);
   U147 : HS65_LH_MX41X7 port map( D0 => n81, S0 => n38, D1 => alu_i(21), S1 =>
                           n34, D2 => n79, S2 => n29, D3 => n21, S3 => n78, Z 
                           => n317);
   U148 : HS65_LH_AND2X4 port map( A => n390, B => n391, Z => n106_port);
   U149 : HS65_LH_MX41X7 port map( D0 => n77, S0 => n38, D1 => n76, S1 => n34, 
                           D2 => n75, S2 => n28, D3 => n74, S3 => n23, Z => 
                           n316);
   U150 : HS65_LH_MX41X7 port map( D0 => n84, S0 => n38, D1 => n85, S1 => n34, 
                           D2 => n86, S2 => n29, D3 => n87, S3 => n24, Z => 
                           n145_port);
   U151 : HS65_LH_MX41X7 port map( D0 => n85, S0 => n37, D1 => n84, S1 => n33, 
                           D2 => n83, S2 => n28, D3 => n82, S3 => n22, Z => 
                           n266);
   U152 : HS65_LH_MX41X7 port map( D0 => n84, S0 => n37, D1 => n83, S1 => n33, 
                           D2 => n82, S2 => n28, D3 => n81, S3 => n22, Z => 
                           n278);
   U153 : HS65_LH_NOR2AX3 port map( A => n69, B => n39, Z => n315);
   U154 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n88, D1 => n32, S1 =>
                           alu_i(30), D2 => n90, S2 => n29, D3 => n300, S3 => 
                           n24, Z => n144_port);
   U155 : HS65_LH_MX41X7 port map( D0 => alu_i(38), S0 => n38, D1 => n523, S1 
                           => n34, D2 => n524, S2 => n29, D3 => alu_i(41), S3 
                           => n25, Z => n263);
   U156 : HS65_LH_MX41X7 port map( D0 => alu_i(13), S0 => n38, D1 => alu_i(12),
                           S1 => n34, D2 => n70, S2 => n29, D3 => n69, S3 => 
                           n24, Z => n188_port);
   U157 : HS65_LH_NAND2X7 port map( A => n193_port, B => n584, Z => n186_port);
   U158 : HS65_LH_MX41X7 port map( D0 => n81, S0 => n38, D1 => n82, S1 => n34, 
                           D2 => n83, S2 => n29, D3 => n84, S3 => n25, Z => 
                           n130_port);
   U159 : HS65_LH_MX41X7 port map( D0 => n36, S0 => n88, D1 => n87, S1 => n33, 
                           D2 => n86, S2 => n28, D3 => n85, S3 => n22, Z => 
                           n212_port);
   U160 : HS65_LH_MX41X7 port map( D0 => n517, S0 => n38, D1 => n518, S1 => n34
                           , D2 => n519, S2 => n29, D3 => n520, S3 => n24, Z =>
                           n325);
   U161 : HS65_LH_MX41X7 port map( D0 => n83, S0 => n38, D1 => n84, S1 => n34, 
                           D2 => n85, S2 => n29, D3 => n86, S3 => n24, Z => 
                           n157_port);
   U162 : HS65_LH_MX41X7 port map( D0 => n82, S0 => n37, D1 => n83, S1 => n33, 
                           D2 => n84, S2 => n28, D3 => n85, S3 => n23, Z => 
                           n114_port);
   U163 : HS65_LH_MX41X7 port map( D0 => alu_i(21), S0 => n38, D1 => n81, S1 =>
                           n34, D2 => n82, S2 => n29, D3 => n83, S3 => n23, Z 
                           => n142_port);
   U164 : HS65_LH_MX41X7 port map( D0 => n74, S0 => n37, D1 => alu_i(14), S1 =>
                           n33, D2 => alu_i(13), S2 => n28, D3 => alu_i(12), S3
                           => n23, Z => n302);
   U165 : HS65_LH_MX41X7 port map( D0 => n75, S0 => n38, D1 => n74, S1 => n34, 
                           D2 => alu_i(14), S2 => n29, D3 => alu_i(13), S3 => 
                           n24, Z => n336);
   U166 : HS65_LH_MX41X7 port map( D0 => n76, S0 => n38, D1 => n75, S1 => n34, 
                           D2 => n74, S2 => n29, D3 => alu_i(14), S3 => n24, Z 
                           => n326);
   U167 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n87, D1 => n86, S1 =>
                           n33, D2 => n85, S2 => n28, D3 => n84, S3 => n22, Z 
                           => n229);
   U168 : HS65_LH_MX41X7 port map( D0 => n36, S0 => alu_i(30), D1 => n32, S1 =>
                           n88, D2 => n87, S2 => n28, D3 => n86, S3 => n22, Z 
                           => n268);
   U169 : HS65_LH_AND2X4 port map( A => n445, B => n587, Z => n442);
   U170 : HS65_LH_MX41X7 port map( D0 => n86, S0 => n37, D1 => n85, S1 => n33, 
                           D2 => n84, S2 => n28, D3 => n83, S3 => n22, Z => 
                           n254);
   U171 : HS65_LH_MX41X7 port map( D0 => n83, S0 => n37, D1 => n82, S1 => n33, 
                           D2 => n81, S2 => n28, D3 => alu_i(21), S3 => n23, Z 
                           => n292);
   U172 : HS65_LH_MX41X7 port map( D0 => n82, S0 => n37, D1 => n81, S1 => n33, 
                           D2 => alu_i(21), S2 => n28, D3 => n79, S3 => n23, Z 
                           => n306);
   U173 : HS65_LH_CBI4I6X5 port map( A => n69, B => n55, C => n123_port, D => 
                           n565, Z => n440);
   U174 : HS65_LH_CBI4I6X5 port map( A => n70, B => n55, C => n40, D => n564, Z
                           => n358);
   U175 : HS65_LH_CBI4I6X5 port map( A => n523, B => n55, C => n123_port, D => 
                           n535, Z => n249);
   U176 : HS65_LH_CBI4I6X5 port map( A => n524, B => n55, C => n40, D => n545, 
                           Z => n224_port);
   U177 : HS65_LH_AO222X4 port map( A => n34, B => n524, C => n27, D => 
                           alu_i(41), E => n36, F => n523, Z => n247);
   U178 : HS65_LH_AND2X4 port map( A => n448, B => n594, Z => n195_port);
   U179 : HS65_LH_MX41X7 port map( D0 => n518, S0 => n38, D1 => n519, S1 => n34
                           , D2 => n520, S2 => n29, D3 => alu_i(37), S3 => n25,
                           Z => n313);
   U180 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n78, D1 => n79, S1 =>
                           n33, D2 => alu_i(21), S2 => n28, D3 => n81, S3 => 
                           n22, Z => n111_port);
   U181 : HS65_LH_MX41X7 port map( D0 => n79, S0 => n38, D1 => alu_i(21), S1 =>
                           n34, D2 => n81, S2 => n29, D3 => n82, S3 => n24, Z 
                           => n154_port);
   U182 : HS65_LH_MX41X7 port map( D0 => n519, S0 => n37, D1 => n520, S1 => n33
                           , D2 => alu_i(37), S2 => n28, D3 => alu_i(38), S3 =>
                           n23, Z => n299);
   U183 : HS65_LH_MX41X7 port map( D0 => n520, S0 => n38, D1 => alu_i(37), S1 
                           => n34, D2 => alu_i(38), S2 => n29, D3 => n523, S3 
                           => n24, Z => n334);
   U184 : HS65_LH_MX41X7 port map( D0 => n85, S0 => n196_port, D1 => n86, S1 =>
                           n34, D2 => n87, S2 => n29, D3 => n88, S3 => n25, Z 
                           => n133_port);
   U185 : HS65_LH_MX41X7 port map( D0 => n36, S0 => alu_i(30), D1 => n90, S1 =>
                           n34, D2 => n300, S2 => n29, D3 => n517, S3 => n25, Z
                           => n132_port);
   U186 : HS65_LH_MX41X7 port map( D0 => n300, S0 => n37, D1 => n90, S1 => n33,
                           D2 => n27, S2 => alu_i(30), D3 => n88, S3 => n22, Z 
                           => n231);
   U187 : HS65_LH_MX41X7 port map( D0 => n300, S0 => n38, D1 => n517, S1 => n34
                           , D2 => n518, S2 => n29, D3 => n519, S3 => n24, Z =>
                           n335);
   U188 : HS65_LH_MX41X7 port map( D0 => n79, S0 => n38, D1 => n32, S1 => n78, 
                           D2 => n77, S2 => n29, D3 => n76, S3 => n24, Z => 
                           n337);
   U189 : HS65_LH_MX41X7 port map( D0 => n90, S0 => n37, D1 => n300, S1 => n33,
                           D2 => n517, S2 => n28, D3 => n518, S3 => n23, Z => 
                           n119_port);
   U190 : HS65_LH_MX41X7 port map( D0 => n90, S0 => n37, D1 => n32, S1 => 
                           alu_i(30), D2 => n88, S2 => n27, D3 => n87, S3 => 
                           n22, Z => n256);
   U191 : HS65_LH_NOR2X6 port map( A => n525, B => n39, Z => n216_port);
   U192 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n78, D1 => n77, S1 =>
                           n33, D2 => n76, S2 => n28, D3 => n75, S3 => n23, Z 
                           => n305);
   U193 : HS65_LH_MX41X7 port map( D0 => alu_i(21), S0 => n38, D1 => n79, S1 =>
                           n34, D2 => n27, S2 => n78, D3 => n77, S3 => n23, Z 
                           => n327);
   U194 : HS65_LH_MX41X7 port map( D0 => alu_i(14), S0 => n38, D1 => alu_i(13),
                           S1 => n33, D2 => alu_i(12), S2 => n28, D3 => n70, S3
                           => n23, Z => n314);
   U195 : HS65_LH_MX41X7 port map( D0 => n86, S0 => n37, D1 => n87, S1 => n33, 
                           D2 => n88, S2 => n28, D3 => alu_i(30), S3 => n23, Z 
                           => n120_port);
   U196 : HS65_LH_MX41X7 port map( D0 => n36, S0 => n87, D1 => n32, S1 => n88, 
                           D2 => n27, S2 => alu_i(30), D3 => n90, S3 => n24, Z 
                           => n156_port);
   U197 : HS65_LH_MX41X7 port map( D0 => n77, S0 => n38, D1 => n32, S1 => n78, 
                           D2 => n79, S2 => n29, D3 => alu_i(21), S3 => n25, Z 
                           => n128_port);
   U198 : HS65_LH_MX41X7 port map( D0 => n517, S0 => n37, D1 => n300, S1 => n32
                           , D2 => n90, S2 => n27, D3 => alu_i(30), S3 => n22, 
                           Z => n214_port);
   U199 : HS65_LH_NAND2X7 port map( A => n434, B => n438, Z => n101_port);
   U200 : HS65_LH_MX41X7 port map( D0 => n76, S0 => n37, D1 => n77, S1 => n32, 
                           D2 => n27, S2 => n78, D3 => n79, S3 => n21, Z => 
                           n140_port);
   U201 : HS65_LH_AND2X4 port map( A => n192_port, B => n581, Z => n118_port);
   U202 : HS65_LH_AO22X9 port map( A => n196_port, B => n70, C => n32, D => n69
                           , Z => n303);
   U203 : HS65_LH_AO22X9 port map( A => n36, B => n524, C => n32, D => 
                           alu_i(41), Z => n222_port);
   U204 : HS65_LH_MX41X7 port map( D0 => alu_i(37), S0 => n38, D1 => alu_i(38),
                           S1 => n34, D2 => n523, S2 => n29, D3 => n524, S3 => 
                           n24, Z => n324);
   U205 : HS65_LH_MX41X7 port map( D0 => alu_i(14), S0 => n196_port, D1 => n74,
                           S1 => n32, D2 => n75, S2 => n27, D3 => n76, S3 => 
                           n21, Z => n173_port);
   U206 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n133_port, D1 => n301, S1 
                           => n132_port, D2 => n304, S2 => n313, D3 => n374, S3
                           => n263, Z => n387);
   U207 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n120_port, D1 => n7, S1 => 
                           n119_port, D2 => n304, S2 => n299, D3 => n374, S3 =>
                           n247, Z => n360);
   U208 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n156_port, D1 => n8, S1 => 
                           n335, D2 => n304, S2 => n334, D3 => n374, S3 => 
                           n222_port, Z => n239);
   U209 : HS65_LH_MX41X7 port map( D0 => n74, S0 => n37, D1 => n75, S1 => n33, 
                           D2 => n76, S2 => n28, D3 => n77, S3 => n22, Z => 
                           n164_port);
   U210 : HS65_LH_MX41X7 port map( D0 => n75, S0 => n37, D1 => n76, S1 => n32, 
                           D2 => n77, S2 => n27, D3 => n21, S3 => n78, Z => 
                           n152_port);
   U211 : HS65_LH_AO222X4 port map( A => n313, B => n301, C => n263, D => n304,
                           E => n132_port, F => n17, Z => n174_port);
   U212 : HS65_LH_AO222X4 port map( A => n326, B => n8, C => n188_port, D => 
                           n304, E => n327, F => n17, Z => n276);
   U213 : HS65_LH_AO222X4 port map( A => n314, B => n7, C => n304, D => n315, E
                           => n316, F => n18, Z => n129_port);
   U214 : HS65_LH_AO222X4 port map( A => n302, B => n8, C => n303, D => n304, E
                           => n305, F => n18, Z => n112_port);
   U215 : HS65_LH_AO222X4 port map( A => n336, B => n7, C => n576, D => n304, E
                           => n337, F => n17, Z => n290);
   U216 : HS65_LH_MX41X7 port map( D0 => n518, S0 => n36, D1 => n517, S1 => n33
                           , D2 => n300, S2 => n27, D3 => n90, S3 => n21, Z => 
                           n269);
   U217 : HS65_LH_AO222X4 port map( A => n324, B => n301, C => n304, D => 
                           n216_port, E => n325, F => n18, Z => n143_port);
   U218 : HS65_LH_AO222X4 port map( A => n299, B => n7, C => n247, D => n304, E
                           => n119_port, F => n17, Z => n166_port);
   U219 : HS65_LH_AO222X4 port map( A => n334, B => n8, C => n222_port, D => 
                           n304, E => n335, F => n18, Z => n155_port);
   U220 : HS65_LH_MX41X7 port map( D0 => n520, S0 => n196_port, D1 => n519, S1 
                           => n32, D2 => n518, S2 => n27, D3 => n517, S3 => n21
                           , Z => n226_port);
   U221 : HS65_LH_MX41X7 port map( D0 => n519, S0 => n37, D1 => n518, S1 => n32
                           , D2 => n517, S2 => n27, D3 => n300, S3 => n22, Z =>
                           n251);
   U222 : HS65_LH_MX41X7 port map( D0 => alu_i(37), S0 => n36, D1 => n520, S1 
                           => n32, D2 => n519, S2 => n27, D3 => n518, S3 => n21
                           , Z => n209_port);
   U223 : HS65_LH_OAI21X3 port map( A => n74, B => n97, C => n40, Z => 
                           n168_port);
   U224 : HS65_LH_OAI21X3 port map( A => n75, B => n54, C => n40, Z => 
                           n159_port);
   U225 : HS65_LH_OAI21X3 port map( A => n76, B => n97, C => n123_port, Z => 
                           n147_port);
   U226 : HS65_LH_OAI21X3 port map( A => n77, B => n54, C => n40, Z => 
                           n135_port);
   U227 : HS65_LH_OAI21X3 port map( A => n79, B => n97, C => n123_port, Z => 
                           n429);
   U228 : HS65_LH_OAI21X3 port map( A => n81, B => n54, C => n40, Z => n416);
   U229 : HS65_LH_OAI21X3 port map( A => n82, B => n97, C => n123_port, Z => 
                           n410);
   U230 : HS65_LH_OAI21X3 port map( A => n83, B => n54, C => n40, Z => n404);
   U231 : HS65_LH_OAI21X3 port map( A => n84, B => n97, C => n123_port, Z => 
                           n398);
   U232 : HS65_LH_OAI21X3 port map( A => n85, B => n54, C => n123_port, Z => 
                           n389);
   U233 : HS65_LH_OAI21X3 port map( A => n86, B => n97, C => n40, Z => n382);
   U234 : HS65_LH_OAI21X3 port map( A => n88, B => n54, C => n123_port, Z => 
                           n369);
   U235 : HS65_LH_OAI21X3 port map( A => n518, B => n97, C => n40, Z => n319);
   U236 : HS65_LH_OAI21X3 port map( A => n519, B => n54, C => n123_port, Z => 
                           n308);
   U237 : HS65_LH_OAI21X3 port map( A => n520, B => n97, C => n40, Z => n294);
   U238 : HS65_LH_OAI21X3 port map( A => n90, B => n97, C => n123_port, Z => 
                           n345);
   U239 : HS65_LH_OAI21X3 port map( A => n300, B => n54, C => n40, Z => n339);
   U240 : HS65_LH_OAI21X3 port map( A => n517, B => n97, C => n123_port, Z => 
                           n329);
   U241 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n306, D1 => n7, S1 => n305,
                           D2 => n304, S2 => n302, D3 => n374, S3 => n303, Z =>
                           n252);
   U242 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n292, D1 => n8, S1 => n337,
                           D2 => n304, S2 => n336, D3 => n374, S3 => n576, Z =>
                           n227);
   U243 : HS65_LH_MX41X7 port map( D0 => n17, S0 => n278, D1 => n301, S1 => 
                           n327, D2 => n304, S2 => n326, D3 => n374, S3 => 
                           n188_port, Z => n210_port);
   U244 : HS65_LH_NAND2X7 port map( A => n434, B => n435, Z => n100_port);
   U245 : HS65_LH_OAI21X3 port map( A => n78, B => n97, C => n40, Z => 
                           n122_port);
   U246 : HS65_LH_OAI21X3 port map( A => n87, B => n97, C => n40, Z => n376);
   U247 : HS65_LH_IVX9 port map( A => n36, Z => n39);
   U248 : HS65_LH_IVX9 port map( A => n6, Z => n17);
   U249 : HS65_LH_NAND3X5 port map( A => n243, B => n244, C => n245, Z => 
                           alu_o(29));
   U250 : HS65_LH_AOI22X6 port map( A => N128, B => n48, C => n584, D => n250, 
                           Z => n243);
   U251 : HS65_LH_AOI212X4 port map( A => n13, B => n524, C => N160, D => n53, 
                           E => n246, Z => n245);
   U252 : HS65_LH_AOI212X4 port map( A => n579, B => n247, C => n523, D => n248
                           , E => n249, Z => n244);
   U253 : HS65_LH_NAND3X5 port map( A => n218_port, B => n219_port, C => 
                           n220_port, Z => alu_o(30));
   U254 : HS65_LH_AOI22X6 port map( A => N129, B => n48, C => n584, D => 
                           n225_port, Z => n218_port);
   U255 : HS65_LH_AOI212X4 port map( A => n13, B => alu_i(41), C => N161, D => 
                           n53, E => n221_port, Z => n220_port);
   U256 : HS65_LH_AOI212X4 port map( A => n579, B => n222_port, C => n524, D =>
                           n223_port, E => n224_port, Z => n219_port);
   U257 : HS65_LH_NAND3X5 port map( A => n353, B => n354, C => n355, Z => 
                           alu_o(1));
   U258 : HS65_LH_AOI22X6 port map( A => N100, B => n48, C => n581, D => n359, 
                           Z => n353);
   U259 : HS65_LH_AOI212X4 port map( A => n12, B => alu_i(12), C => N132, D => 
                           n53, E => n356, Z => n355);
   U260 : HS65_LH_AOI212X4 port map( A => n583, B => n303, C => n70, D => n357,
                           E => n358, Z => n354);
   U261 : HS65_LH_BFX9 port map( A => n97, Z => n54);
   U262 : HS65_LH_NAND2X7 port map( A => n391, B => n442, Z => n97);
   U263 : HS65_LH_BFX9 port map( A => n123_port, Z => n40);
   U264 : HS65_LH_NAND2X7 port map( A => n438, B => n442, Z => n123_port);
   U265 : HS65_LH_AO22X9 port map( A => n302, B => n17, C => n303, D => n7, Z 
                           => n165_port);
   U266 : HS65_LH_AO22X9 port map( A => n336, B => n17, C => n576, D => n8, Z 
                           => n153_port);
   U267 : HS65_LH_AO22X9 port map( A => n326, B => n17, C => n188_port, D => 
                           n301, Z => n141_port);
   U268 : HS65_LH_AO22X9 port map( A => n313, B => n17, C => n263, D => n7, Z 
                           => n131_port);
   U269 : HS65_LH_AO22X9 port map( A => n299, B => n17, C => n247, D => n8, Z 
                           => n116_port);
   U270 : HS65_LH_AO22X9 port map( A => n334, B => n17, C => n222_port, D => 
                           n301, Z => n291);
   U271 : HS65_LH_BFX9 port map( A => n199_port, Z => n19);
   U272 : HS65_LH_BFX9 port map( A => n105_port, Z => n43);
   U273 : HS65_LH_NOR2AX3 port map( A => n390, B => n589, Z => n105_port);
   U274 : HS65_LH_BFX9 port map( A => n99_port, Z => n50);
   U275 : HS65_LH_NOR2X6 port map( A => n590, B => n437, Z => n99_port);
   U276 : HS65_LH_BFX9 port map( A => n46, Z => n48);
   U277 : HS65_LH_IVX9 port map( A => n438, Z => n589);
   U278 : HS65_LH_BFX9 port map( A => n46, Z => n47);
   U279 : HS65_LH_AND2X4 port map( A => n434, B => n391, Z => n102_port);
   U280 : HS65_LH_BFX9 port map( A => n197_port, Z => n30);
   U281 : HS65_LH_BFX9 port map( A => n197_port, Z => n31);
   U282 : HS65_LH_BFX9 port map( A => n26, Z => n27);
   U283 : HS65_LH_IVX9 port map( A => n264, Z => n573);
   U284 : HS65_LH_AND2X4 port map( A => n434, B => n436, Z => n103_port);
   U285 : HS65_LH_BFX9 port map( A => n26, Z => n29);
   U286 : HS65_LH_BFX9 port map( A => n26, Z => n28);
   U287 : HS65_LH_BFX9 port map( A => n199_port, Z => n20);
   U288 : HS65_LH_IVX9 port map( A => n6, Z => n18);
   U289 : HS65_LH_BFX9 port map( A => n537, Z => n542);
   U290 : HS65_LH_BFX9 port map( A => n537, Z => n541);
   U291 : HS65_LH_BFX9 port map( A => n536, Z => n540);
   U292 : HS65_LH_BFX9 port map( A => n536, Z => n539);
   U293 : HS65_LH_BFX9 port map( A => n536, Z => n538);
   U294 : HS65_LH_BFX9 port map( A => n46, Z => n49);
   U295 : HS65_LH_BFX9 port map( A => n537, Z => n543);
   U296 : HS65_LH_AO22X9 port map( A => N167, B => n63, C => HI_LO_c_LO_4_port,
                           D => n57, Z => n457);
   U297 : HS65_LH_AO22X9 port map( A => N168, B => n63, C => HI_LO_c_LO_5_port,
                           D => n57, Z => n458);
   U298 : HS65_LH_AO22X9 port map( A => N169, B => n62, C => HI_LO_c_LO_6_port,
                           D => n57, Z => n459);
   U299 : HS65_LH_AO22X9 port map( A => N170, B => n61, C => HI_LO_c_LO_7_port,
                           D => n57, Z => n460);
   U300 : HS65_LH_AO22X9 port map( A => N171, B => n66, C => HI_LO_c_LO_8_port,
                           D => n59, Z => n461);
   U301 : HS65_LH_AO22X9 port map( A => N172, B => n66, C => HI_LO_c_LO_9_port,
                           D => n58, Z => n462);
   U302 : HS65_LH_AO22X9 port map( A => N173, B => n65, C => HI_LO_c_LO_10_port
                           , D => n57, Z => n463);
   U303 : HS65_LH_AO22X9 port map( A => N174, B => n65, C => HI_LO_c_LO_11_port
                           , D => n60, Z => n464);
   U304 : HS65_LH_AO22X9 port map( A => N175, B => n65, C => HI_LO_c_LO_12_port
                           , D => n60, Z => n465);
   U305 : HS65_LH_AO22X9 port map( A => N176, B => n65, C => HI_LO_c_LO_13_port
                           , D => n60, Z => n466);
   U306 : HS65_LH_AO22X9 port map( A => N177, B => n65, C => HI_LO_c_LO_14_port
                           , D => n60, Z => n467);
   U307 : HS65_LH_AO22X9 port map( A => N178, B => n65, C => HI_LO_c_LO_15_port
                           , D => n60, Z => n468);
   U308 : HS65_LH_AO22X9 port map( A => N199, B => n64, C => HI_LO_c_HI_4_port,
                           D => n59, Z => n489);
   U309 : HS65_LH_AO22X9 port map( A => N200, B => n64, C => HI_LO_c_HI_5_port,
                           D => n59, Z => n490);
   U310 : HS65_LH_AO22X9 port map( A => N201, B => n64, C => HI_LO_c_HI_6_port,
                           D => n59, Z => n491);
   U311 : HS65_LH_AO22X9 port map( A => N202, B => n64, C => HI_LO_c_HI_7_port,
                           D => n59, Z => n492);
   U312 : HS65_LH_AO22X9 port map( A => N203, B => n64, C => HI_LO_c_HI_8_port,
                           D => n59, Z => n493);
   U313 : HS65_LH_AO22X9 port map( A => N204, B => n64, C => HI_LO_c_HI_9_port,
                           D => n59, Z => n494);
   U314 : HS65_LH_AO22X9 port map( A => N205, B => n64, C => HI_LO_c_HI_10_port
                           , D => n59, Z => n495);
   U315 : HS65_LH_AO22X9 port map( A => N206, B => n64, C => HI_LO_c_HI_11_port
                           , D => n59, Z => n496);
   U316 : HS65_LH_AO22X9 port map( A => N207, B => n64, C => HI_LO_c_HI_12_port
                           , D => n59, Z => n497);
   U317 : HS65_LH_AO22X9 port map( A => N208, B => n64, C => HI_LO_c_HI_13_port
                           , D => n59, Z => n498);
   U318 : HS65_LH_AO22X9 port map( A => N209, B => n64, C => HI_LO_c_HI_14_port
                           , D => n59, Z => n499);
   U319 : HS65_LH_AO22X9 port map( A => N210, B => n64, C => HI_LO_c_HI_15_port
                           , D => n59, Z => n500);
   U320 : HS65_LH_AO22X9 port map( A => N211, B => n64, C => HI_LO_c_HI_16_port
                           , D => n58, Z => n501);
   U321 : HS65_LH_AO22X9 port map( A => N212, B => n64, C => HI_LO_c_HI_17_port
                           , D => n58, Z => n502);
   U322 : HS65_LH_AO22X9 port map( A => N213, B => n63, C => HI_LO_c_HI_18_port
                           , D => n58, Z => n503);
   U323 : HS65_LH_AO22X9 port map( A => N214, B => n63, C => HI_LO_c_HI_19_port
                           , D => n58, Z => n504);
   U324 : HS65_LH_AO22X9 port map( A => N215, B => n63, C => HI_LO_c_HI_20_port
                           , D => n58, Z => n505);
   U325 : HS65_LH_AO22X9 port map( A => N216, B => n63, C => HI_LO_c_HI_21_port
                           , D => n58, Z => n506);
   U326 : HS65_LH_AO22X9 port map( A => N217, B => n63, C => HI_LO_c_HI_22_port
                           , D => n58, Z => n507);
   U327 : HS65_LH_AO22X9 port map( A => N218, B => n63, C => HI_LO_c_HI_23_port
                           , D => n58, Z => n508);
   U328 : HS65_LH_AO22X9 port map( A => N219, B => n63, C => HI_LO_c_HI_24_port
                           , D => n58, Z => n509);
   U329 : HS65_LH_AO22X9 port map( A => N220, B => n63, C => HI_LO_c_HI_25_port
                           , D => n58, Z => n510);
   U330 : HS65_LH_AO22X9 port map( A => N221, B => n63, C => HI_LO_c_HI_26_port
                           , D => n58, Z => n511);
   U331 : HS65_LH_AO22X9 port map( A => N222, B => n63, C => HI_LO_c_HI_27_port
                           , D => n58, Z => n512);
   U332 : HS65_LH_AO22X9 port map( A => N226, B => n63, C => HI_LO_c_HI_31_port
                           , D => n57, Z => n516);
   U333 : HS65_LH_AO22X9 port map( A => N163, B => n63, C => HI_LO_c_LO_0_port,
                           D => n57, Z => n453);
   U334 : HS65_LH_AO22X9 port map( A => N164, B => n63, C => HI_LO_c_LO_1_port,
                           D => n57, Z => n454);
   U335 : HS65_LH_AO22X9 port map( A => N165, B => n63, C => HI_LO_c_LO_2_port,
                           D => n57, Z => n455);
   U336 : HS65_LH_AO22X9 port map( A => N166, B => n63, C => HI_LO_c_LO_3_port,
                           D => n57, Z => n456);
   U337 : HS65_LH_AO22X9 port map( A => N194, B => n64, C => HI_LO_c_LO_31_port
                           , D => n59, Z => n484);
   U338 : HS65_LH_AO22X9 port map( A => N196, B => n64, C => HI_LO_c_HI_1_port,
                           D => n58, Z => n486);
   U339 : HS65_LH_AO22X9 port map( A => N197, B => n64, C => HI_LO_c_HI_2_port,
                           D => n57, Z => n487);
   U340 : HS65_LH_AO22X9 port map( A => N198, B => n64, C => HI_LO_c_HI_3_port,
                           D => n60, Z => n488);
   U341 : HS65_LH_AO22X9 port map( A => N223, B => n63, C => HI_LO_c_HI_28_port
                           , D => n57, Z => n513);
   U342 : HS65_LH_AO22X9 port map( A => N224, B => n63, C => HI_LO_c_HI_29_port
                           , D => n57, Z => n514);
   U343 : HS65_LH_AO22X9 port map( A => N225, B => n63, C => HI_LO_c_HI_30_port
                           , D => n57, Z => n515);
   U344 : HS65_LH_AO22X9 port map( A => N179, B => n65, C => HI_LO_c_LO_16_port
                           , D => n60, Z => n469);
   U345 : HS65_LH_AO22X9 port map( A => N180, B => n65, C => HI_LO_c_LO_17_port
                           , D => n60, Z => n470);
   U346 : HS65_LH_AO22X9 port map( A => N181, B => n65, C => HI_LO_c_LO_18_port
                           , D => n60, Z => n471);
   U347 : HS65_LH_AO22X9 port map( A => N182, B => n65, C => HI_LO_c_LO_19_port
                           , D => n60, Z => n472);
   U348 : HS65_LH_AO22X9 port map( A => N183, B => n65, C => HI_LO_c_LO_20_port
                           , D => n60, Z => n473);
   U349 : HS65_LH_AO22X9 port map( A => N184, B => n65, C => HI_LO_c_LO_21_port
                           , D => n60, Z => n474);
   U350 : HS65_LH_AO22X9 port map( A => N185, B => n65, C => HI_LO_c_LO_22_port
                           , D => n60, Z => n475);
   U351 : HS65_LH_AO22X9 port map( A => N186, B => n65, C => HI_LO_c_LO_23_port
                           , D => n60, Z => n476);
   U352 : HS65_LH_AO22X9 port map( A => N187, B => n65, C => HI_LO_c_LO_24_port
                           , D => n59, Z => n477);
   U353 : HS65_LH_AO22X9 port map( A => N188, B => n65, C => HI_LO_c_LO_25_port
                           , D => n58, Z => n478);
   U354 : HS65_LH_AO22X9 port map( A => N189, B => n65, C => HI_LO_c_LO_26_port
                           , D => n57, Z => n479);
   U355 : HS65_LH_AO22X9 port map( A => N190, B => n65, C => HI_LO_c_LO_27_port
                           , D => n60, Z => n480);
   U356 : HS65_LH_AO22X9 port map( A => N191, B => n65, C => HI_LO_c_LO_28_port
                           , D => n59, Z => n481);
   U357 : HS65_LH_AO22X9 port map( A => N192, B => n65, C => HI_LO_c_LO_29_port
                           , D => n58, Z => n482);
   U358 : HS65_LH_AO22X9 port map( A => N193, B => n64, C => HI_LO_c_LO_30_port
                           , D => n57, Z => n483);
   U359 : HS65_LH_AO22X9 port map( A => N195, B => n64, C => HI_LO_c_HI_0_port,
                           D => n60, Z => n485);
   U360 : HS65_LH_NOR4ABX4 port map( A => n578, B => n435, C => alu_i(8), D => 
                           alu_i(7), Z => n180_port);
   U361 : HS65_LH_NOR3X4 port map( A => alu_i(7), B => alu_i(9), C => n587, Z 
                           => n434);
   U362 : HS65_LH_AND2X4 port map( A => alu_i(1), B => alu_i(0), Z => n199_port
                           );
   U363 : HS65_LH_AOI222X2 port map( A => n317, B => n17, C => n316, D => n7, E
                           => n178_port, F => alu_i(3), Z => n264);
   U364 : HS65_LH_AOI222X2 port map( A => n144_port, B => n17, C => n325, D => 
                           n8, E => n283, F => alu_i(3), Z => n190_port);
   U365 : HS65_LH_NOR2X6 port map( A => n594, B => alu_i(3), Z => n7);
   U366 : HS65_LH_NOR2X6 port map( A => n594, B => alu_i(3), Z => n8);
   U367 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_4_port, C => 
                           n579, D => n173_port, E => N103, F => n47, Z => 
                           n172_port);
   U368 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_5_port, C => 
                           n579, D => n164_port, E => N104, F => n47, Z => 
                           n163_port);
   U369 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_6_port, C => 
                           n579, D => n152_port, E => N105, F => n47, Z => 
                           n151_port);
   U370 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_7_port, C => 
                           n579, D => n140_port, E => N106, F => n47, Z => 
                           n139_port);
   U371 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_8_port, C => 
                           n579, D => n128_port, E => N107, F => n47, Z => 
                           n127_port);
   U372 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_9_port, C => 
                           n579, D => n111_port, E => N108, F => n47, Z => 
                           n110_port);
   U373 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_10_port, C => 
                           n579, D => n154_port, E => N109, F => n47, Z => n427
                           );
   U374 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_11_port, C => 
                           n579, D => n142_port, E => N110, F => n47, Z => n420
                           );
   U375 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_12_port, C => 
                           n579, D => n130_port, E => N111, F => n47, Z => n414
                           );
   U376 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_13_port, C => 
                           n579, D => n114_port, E => N112, F => n47, Z => n408
                           );
   U377 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_14_port, C => 
                           n579, D => n157_port, E => N113, F => n47, Z => n402
                           );
   U378 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_15_port, C => 
                           n579, D => n145_port, E => N114, F => n47, Z => n395
                           );
   U379 : HS65_LH_NOR2AX3 port map( A => alu_i(0), B => alu_i(1), Z => 
                           n197_port);
   U380 : HS65_LH_AOI212X4 port map( A => alu_i(46), B => n180_port, C => n56, 
                           D => n562, E => n42, Z => n175_port);
   U381 : HS65_LH_IVX9 port map( A => alu_i(46), Z => n562);
   U382 : HS65_LH_AOI212X4 port map( A => alu_i(69), B => n180_port, C => n56, 
                           D => n547, E => n42, Z => n280);
   U383 : HS65_LH_IVX9 port map( A => alu_i(69), Z => n547);
   U384 : HS65_LH_NOR2X6 port map( A => n96, B => alu_i(4), Z => n113_port);
   U385 : HS65_LH_NOR2X6 port map( A => n594, B => alu_i(3), Z => n301);
   U386 : HS65_LH_IVX9 port map( A => alu_i(3), Z => n593);
   U387 : HS65_LH_NOR2X6 port map( A => n593, B => alu_i(2), Z => n304);
   U388 : HS65_LH_OAI212X5 port map( A => n185_port, B => n72, C => n575, D => 
                           n186_port, E => n187_port, Z => n184_port);
   U389 : HS65_LH_IVX9 port map( A => n188_port, Z => n575);
   U390 : HS65_LH_CBI4I1X5 port map( A => n56, B => n72, C => n42, D => 
                           alu_i(45), Z => n187_port);
   U391 : HS65_LH_AOI212X4 port map( A => alu_i(45), B => n180_port, C => n56, 
                           D => n563, E => n42, Z => n185_port);
   U392 : HS65_LH_OAI212X5 port map( A => n261, B => n522, C => n567, D => 
                           n208_port, E => n262, Z => n260);
   U393 : HS65_LH_IVX9 port map( A => n263, Z => n567);
   U394 : HS65_LH_CBI4I1X5 port map( A => n56, B => n522, C => n42, D => 
                           alu_i(70), Z => n262);
   U395 : HS65_LH_AOI212X4 port map( A => alu_i(70), B => n180_port, C => n56, 
                           D => n546, E => n42, Z => n261);
   U396 : HS65_LH_OAI212X5 port map( A => alu_i(42), B => n55, C => n9, D => 
                           n565, E => n441, Z => n439);
   U397 : HS65_LH_AOI12X2 port map( A => n583, B => n196_port, C => n42, Z => 
                           n441);
   U398 : HS65_LH_OAI212X5 port map( A => alu_i(72), B => n55, C => n9, D => 
                           n545, E => n41, Z => n223_port);
   U399 : HS65_LH_OAI212X5 port map( A => alu_i(43), B => n97, C => n10, D => 
                           n564, E => n41, Z => n357);
   U400 : HS65_LH_NOR2X6 port map( A => n6, B => alu_i(4), Z => n193_port);
   U401 : HS65_LH_OAI212X5 port map( A => alu_i(54), B => n54, C => n10, D => 
                           n557, E => n123_port, Z => n415);
   U402 : HS65_LH_IVX9 port map( A => alu_i(54), Z => n557);
   U403 : HS65_LH_OAI212X5 port map( A => alu_i(55), B => n97, C => n10, D => 
                           n556, E => n40, Z => n409);
   U404 : HS65_LH_IVX9 port map( A => alu_i(55), Z => n556);
   U405 : HS65_LH_OAI212X5 port map( A => alu_i(57), B => n54, C => n10, D => 
                           n555, E => n123_port, Z => n396);
   U406 : HS65_LH_IVX9 port map( A => alu_i(57), Z => n555);
   U407 : HS65_LH_OAI212X5 port map( A => alu_i(58), B => n97, C => n10, D => 
                           n554, E => n41, Z => n388);
   U408 : HS65_LH_IVX9 port map( A => alu_i(58), Z => n554);
   U409 : HS65_LH_OAI212X5 port map( A => alu_i(60), B => n54, C => n10, D => 
                           n553, E => n40, Z => n375);
   U410 : HS65_LH_IVX9 port map( A => alu_i(60), Z => n553);
   U411 : HS65_LH_OAI212X5 port map( A => alu_i(61), B => n97, C => n10, D => 
                           n552, E => n123_port, Z => n367);
   U412 : HS65_LH_IVX9 port map( A => alu_i(61), Z => n552);
   U413 : HS65_LH_OAI212X5 port map( A => alu_i(48), B => n55, C => n9, D => 
                           n561, E => n41, Z => n158_port);
   U414 : HS65_LH_IVX9 port map( A => alu_i(48), Z => n561);
   U415 : HS65_LH_OAI212X5 port map( A => alu_i(49), B => n55, C => n9, D => 
                           n560, E => n41, Z => n146_port);
   U416 : HS65_LH_IVX9 port map( A => alu_i(49), Z => n560);
   U417 : HS65_LH_OAI212X5 port map( A => alu_i(51), B => n55, C => n559, D => 
                           n10, E => n123_port, Z => n121_port);
   U418 : HS65_LH_IVX9 port map( A => alu_i(51), Z => n559);
   U419 : HS65_LH_OAI212X5 port map( A => alu_i(66), B => n55, C => n9, D => 
                           n549, E => n41, Z => n318);
   U420 : HS65_LH_IVX9 port map( A => alu_i(66), Z => n549);
   U421 : HS65_LH_AOI32X5 port map( A => n283, B => n593, C => n284, D => 
                           alu_i(69), E => n285, Z => n282);
   U422 : HS65_LH_OAI21X3 port map( A => alu_i(37), B => n54, C => n123_port, Z
                           => n285);
   U423 : HS65_LH_OAI212X5 port map( A => alu_i(52), B => n54, C => n10, D => 
                           n558, E => n41, Z => n428);
   U424 : HS65_LH_IVX9 port map( A => alu_i(52), Z => n558);
   U425 : HS65_LH_OAI212X5 port map( A => alu_i(63), B => n97, C => n10, D => 
                           n551, E => n41, Z => n344);
   U426 : HS65_LH_IVX9 port map( A => alu_i(63), Z => n551);
   U427 : HS65_LH_OAI212X5 port map( A => alu_i(64), B => n54, C => n9, D => 
                           n550, E => n41, Z => n338);
   U428 : HS65_LH_IVX9 port map( A => alu_i(64), Z => n550);
   U429 : HS65_LH_OAI212X5 port map( A => alu_i(67), B => n97, C => n9, D => 
                           n548, E => n41, Z => n307);
   U430 : HS65_LH_IVX9 port map( A => alu_i(67), Z => n548);
   U431 : HS65_LH_AOI32X5 port map( A => n178_port, B => n593, C => n113_port, 
                           D => alu_i(46), E => n179_port, Z => n177_port);
   U432 : HS65_LH_OAI21X3 port map( A => alu_i(14), B => n97, C => n40, Z => 
                           n179_port);
   U433 : HS65_LH_NOR2X6 port map( A => n590, B => alu_i(6), Z => n391);
   U434 : HS65_LH_IVX9 port map( A => alu_i(4), Z => n592);
   U435 : HS65_LH_IVX9 port map( A => alu_i(2), Z => n594);
   U436 : HS65_LH_NOR2X6 port map( A => alu_i(6), B => alu_i(5), Z => n438);
   U437 : HS65_LH_NOR2X6 port map( A => n588, B => alu_i(5), Z => n436);
   U438 : HS65_LH_NOR2X6 port map( A => n593, B => alu_i(4), Z => n448);
   U439 : HS65_LH_NAND4ABX3 port map( A => alu_i(9), B => alu_i(7), C => n588, 
                           D => n587, Z => n437);
   U440 : HS65_LH_AND2X4 port map( A => n448, B => alu_i(2), Z => n192_port);
   U441 : HS65_LH_AO22X9 port map( A => n594, B => n314, C => alu_i(2), D => 
                           n315, Z => n178_port);
   U442 : HS65_LH_AO22X9 port map( A => n594, B => n324, C => alu_i(2), D => 
                           n216_port, Z => n283);
   U443 : HS65_LH_OAI21X3 port map( A => n205_port, B => n525, C => n206_port, 
                           Z => n204_port);
   U444 : HS65_LH_CBI4I1X5 port map( A => n56, B => n525, C => n42, D => 
                           alu_i(73), Z => n206_port);
   U445 : HS65_LH_AOI212X4 port map( A => n56, B => n544, C => alu_i(73), D => 
                           n180_port, E => n207_port, Z => n205_port);
   U446 : HS65_LH_IVX9 port map( A => alu_i(73), Z => n544);
   U447 : HS65_LH_AND2X4 port map( A => n445, B => alu_i(8), Z => n390);
   U448 : HS65_LH_NOR2AX3 port map( A => alu_i(7), B => alu_i(9), Z => n445);
   U449 : HS65_LH_NAND4ABX3 port map( A => n383, B => n384, C => n385, D => 
                           n386, Z => alu_o(16));
   U450 : HS65_LH_MX41X7 port map( D0 => n582, S0 => n316, D1 => n85, S1 => 
                           n388, D2 => n368, S2 => n315, D3 => alu_i(58), S3 =>
                           n389, Z => n384);
   U451 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_16_port, D1 => 
                           n106_port, S1 => n69, D2 => N115, S2 => n49, D3 => 
                           n583, S3 => n266, Z => n383);
   U452 : HS65_LH_AOI222X2 port map( A => N147, B => n52, C => n15, D => 
                           HI_LO_c_HI_16_port, E => n12, F => n86, Z => n385);
   U453 : HS65_LH_NAND4ABX3 port map( A => n377, B => n378, C => n379, D => 
                           n380, Z => alu_o(17));
   U454 : HS65_LH_MX41X7 port map( D0 => n582, S0 => n305, D1 => n86, S1 => 
                           n381, D2 => n368, S2 => n303, D3 => alu_i(59), S3 =>
                           n382, Z => n378);
   U455 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_17_port, D1 => 
                           n106_port, S1 => n70, D2 => N116, S2 => n49, D3 => 
                           n583, S3 => n254, Z => n377);
   U456 : HS65_LH_AOI222X2 port map( A => N148, B => n52, C => n15, D => 
                           HI_LO_c_HI_17_port, E => n12, F => n87, Z => n379);
   U457 : HS65_LH_NAND4ABX3 port map( A => n370, B => n371, C => n372, D => 
                           n373, Z => alu_o(18));
   U458 : HS65_LH_MX41X7 port map( D0 => n582, S0 => n337, D1 => n87, S1 => 
                           n375, D2 => n368, S2 => n576, D3 => alu_i(60), S3 =>
                           n376, Z => n371);
   U459 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_18_port, D1 => 
                           n106_port, S1 => alu_i(12), D2 => N117, S2 => n49, 
                           D3 => n583, S3 => n229, Z => n370);
   U460 : HS65_LH_AOI222X2 port map( A => N149, B => n52, C => n15, D => 
                           HI_LO_c_HI_18_port, E => n12, F => n88, Z => n372);
   U461 : HS65_LH_NAND4ABX3 port map( A => n363, B => n364, C => n365, D => 
                           n366, Z => alu_o(19));
   U462 : HS65_LH_MX41X7 port map( D0 => n582, S0 => n327, D1 => n88, S1 => 
                           n367, D2 => n368, S2 => n188_port, D3 => alu_i(61), 
                           S3 => n369, Z => n364);
   U463 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_19_port, D1 => 
                           n106_port, S1 => alu_i(13), D2 => N118, S2 => n48, 
                           D3 => n583, S3 => n212_port, Z => n363);
   U464 : HS65_LH_AOI222X2 port map( A => N150, B => n52, C => n15, D => 
                           HI_LO_c_HI_19_port, E => n12, F => alu_i(30), Z => 
                           n365);
   U465 : HS65_LH_NAND4ABX3 port map( A => n346, B => n347, C => n348, D => 
                           n349, Z => alu_o(20));
   U466 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_20_port, D1 => 
                           n106_port, S1 => alu_i(14), D2 => N119, S2 => n48, 
                           D3 => n583, S3 => n268, Z => n346);
   U467 : HS65_LH_OAI212X5 port map( A => n350, B => n89, C => n572, D => n281,
                           E => n351, Z => n347);
   U468 : HS65_LH_AOI222X2 port map( A => N151, B => n52, C => n15, D => 
                           HI_LO_c_HI_20_port, E => n12, F => n90, Z => n348);
   U469 : HS65_LH_NAND4ABX3 port map( A => n271, B => n272, C => n273, D => 
                           n274, Z => alu_o(27));
   U470 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_27_port, D1 => 
                           n106_port, S1 => alu_i(21), D2 => N126, S2 => n48, 
                           D3 => n583, S3 => n209_port, Z => n271);
   U471 : HS65_LH_OAI212X5 port map( A => n280, B => n521, C => n570, D => n281
                           , E => n282, Z => n272);
   U472 : HS65_LH_AOI222X2 port map( A => N158, B => n51, C => n14, D => 
                           HI_LO_c_HI_27_port, E => n11, F => alu_i(38), Z => 
                           n273);
   U473 : HS65_LH_NAND4ABX3 port map( A => n340, B => n341, C => n342, D => 
                           n343, Z => alu_o(21));
   U474 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n305, D1 => n582, S1 => 
                           n306, D2 => n90, S2 => n344, D3 => alu_i(63), S3 => 
                           n345, Z => n341);
   U475 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_21_port, D1 => 
                           n106_port, S1 => n74, D2 => N120, S2 => n48, D3 => 
                           n583, S3 => n256, Z => n340);
   U476 : HS65_LH_AOI222X2 port map( A => N152, B => n52, C => n14, D => 
                           HI_LO_c_HI_21_port, E => n11, F => n300, Z => n342);
   U477 : HS65_LH_NAND4ABX3 port map( A => n330, B => n331, C => n332, D => 
                           n333, Z => alu_o(22));
   U478 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n337, D1 => n582, S1 => 
                           n292, D2 => n300, S2 => n338, D3 => alu_i(64), S3 =>
                           n339, Z => n331);
   U479 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_22_port, D1 => 
                           n106_port, S1 => n75, D2 => N121, S2 => n48, D3 => 
                           n583, S3 => n231, Z => n330);
   U480 : HS65_LH_AOI222X2 port map( A => N153, B => n51, C => n14, D => 
                           HI_LO_c_HI_22_port, E => n11, F => n517, Z => n332);
   U481 : HS65_LH_NAND4ABX3 port map( A => n320, B => n321, C => n322, D => 
                           n323, Z => alu_o(23));
   U482 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n327, D1 => n582, S1 => 
                           n278, D2 => n517, S2 => n328, D3 => alu_i(65), S3 =>
                           n329, Z => n321);
   U483 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_23_port, D1 => 
                           n106_port, S1 => n76, D2 => N122, S2 => n48, D3 => 
                           n583, S3 => n214_port, Z => n320);
   U484 : HS65_LH_AOI222X2 port map( A => N154, B => n51, C => n14, D => 
                           HI_LO_c_HI_23_port, E => n11, F => n518, Z => n322);
   U485 : HS65_LH_NAND4ABX3 port map( A => n309, B => n310, C => n311, D => 
                           n312, Z => alu_o(24));
   U486 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n317, D1 => n582, S1 => 
                           n266, D2 => n518, S2 => n318, D3 => alu_i(66), S3 =>
                           n319, Z => n310);
   U487 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_24_port, D1 => 
                           n106_port, S1 => n77, D2 => N123, S2 => n48, D3 => 
                           n583, S3 => n269, Z => n309);
   U488 : HS65_LH_AOI222X2 port map( A => N155, B => n51, C => n14, D => 
                           HI_LO_c_HI_24_port, E => n11, F => n519, Z => n311);
   U489 : HS65_LH_NAND4ABX3 port map( A => n295, B => n296, C => n297, D => 
                           n298, Z => alu_o(25));
   U490 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n306, D1 => n582, S1 => 
                           n254, D2 => n519, S2 => n307, D3 => alu_i(67), S3 =>
                           n308, Z => n296);
   U491 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_25_port, D1 => 
                           n106_port, S1 => n78, D2 => N124, S2 => n48, D3 => 
                           n583, S3 => n251, Z => n295);
   U492 : HS65_LH_AOI222X2 port map( A => N156, B => n51, C => n14, D => 
                           HI_LO_c_HI_25_port, E => n11, F => n520, Z => n297);
   U493 : HS65_LH_NAND4ABX3 port map( A => n286, B => n287, C => n288, D => 
                           n289, Z => alu_o(26));
   U494 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n292, D1 => n582, S1 => 
                           n229, D2 => n520, S2 => n293, D3 => alu_i(68), S3 =>
                           n294, Z => n287);
   U495 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_26_port, D1 => 
                           n106_port, S1 => n79, D2 => N125, S2 => n48, D3 => 
                           n583, S3 => n226_port, Z => n286);
   U496 : HS65_LH_AOI222X2 port map( A => N157, B => n51, C => n14, D => 
                           HI_LO_c_HI_26_port, E => n11, F => alu_i(37), Z => 
                           n288);
   U497 : HS65_LH_NAND4ABX3 port map( A => n169_port, B => n170_port, C => 
                           n171_port, D => n172_port, Z => alu_o(4));
   U498 : HS65_LH_AO222X4 port map( A => n128_port, B => n115_port, C => 
                           n133_port, D => n118_port, E => n174_port, F => 
                           n117_port, Z => n170_port);
   U499 : HS65_LH_OAI212X5 port map( A => n175_port, B => n73, C => n571, D => 
                           n176_port, E => n177_port, Z => n169_port);
   U500 : HS65_LH_AOI222X2 port map( A => N135, B => n51, C => n14, D => 
                           HI_LO_c_HI_4_port, E => n11, F => n74, Z => 
                           n171_port);
   U501 : HS65_LH_NAND4ABX3 port map( A => n160_port, B => n161_port, C => 
                           n162_port, D => n163_port, Z => alu_o(5));
   U502 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n120_port, D1 => n580
                           , S1 => n114_port, D2 => n74, S2 => n167_port, D3 =>
                           alu_i(47), S3 => n168_port, Z => n160_port);
   U503 : HS65_LH_AO222X4 port map( A => n165_port, B => n113_port, C => 
                           n111_port, D => n115_port, E => n166_port, F => 
                           n117_port, Z => n161_port);
   U504 : HS65_LH_AOI222X2 port map( A => N136, B => n51, C => n15, D => 
                           HI_LO_c_HI_5_port, E => n11, F => n75, Z => 
                           n162_port);
   U505 : HS65_LH_NAND4ABX3 port map( A => n148_port, B => n149_port, C => 
                           n150_port, D => n151_port, Z => alu_o(6));
   U506 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n156_port, D1 => n580
                           , S1 => n157_port, D2 => n75, S2 => n158_port, D3 =>
                           alu_i(48), S3 => n159_port, Z => n148_port);
   U507 : HS65_LH_AO222X4 port map( A => n153_port, B => n113_port, C => 
                           n154_port, D => n115_port, E => n155_port, F => 
                           n117_port, Z => n149_port);
   U508 : HS65_LH_AOI222X2 port map( A => N137, B => n51, C => n14, D => 
                           HI_LO_c_HI_6_port, E => n11, F => n76, Z => 
                           n150_port);
   U509 : HS65_LH_NAND4ABX3 port map( A => n136_port, B => n137_port, C => 
                           n138_port, D => n139_port, Z => alu_o(7));
   U510 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n144_port, D1 => n580
                           , S1 => n145_port, D2 => n76, S2 => n146_port, D3 =>
                           alu_i(49), S3 => n147_port, Z => n136_port);
   U511 : HS65_LH_AO222X4 port map( A => n141_port, B => n113_port, C => 
                           n142_port, D => n115_port, E => n143_port, F => 
                           n117_port, Z => n137_port);
   U512 : HS65_LH_AOI222X2 port map( A => N138, B => n51, C => n14, D => 
                           HI_LO_c_HI_7_port, E => n11, F => n77, Z => 
                           n138_port);
   U513 : HS65_LH_NAND4ABX3 port map( A => n124_port, B => n125_port, C => 
                           n126_port, D => n127_port, Z => alu_o(8));
   U514 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n132_port, D1 => n580
                           , S1 => n133_port, D2 => n77, S2 => n134_port, D3 =>
                           alu_i(50), S3 => n135_port, Z => n124_port);
   U515 : HS65_LH_AO222X4 port map( A => n129_port, B => n113_port, C => 
                           n130_port, D => n115_port, E => n131_port, F => 
                           n117_port, Z => n125_port);
   U516 : HS65_LH_AOI222X2 port map( A => N139, B => n51, C => n14, D => 
                           HI_LO_c_HI_8_port, E => n11, F => n78, Z => 
                           n126_port);
   U517 : HS65_LH_NAND4ABX3 port map( A => n107_port, B => n108_port, C => 
                           n109_port, D => n110_port, Z => alu_o(9));
   U518 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n119_port, D1 => n580
                           , S1 => n120_port, D2 => n78, S2 => n121_port, D3 =>
                           alu_i(51), S3 => n122_port, Z => n107_port);
   U519 : HS65_LH_AO222X4 port map( A => n112_port, B => n113_port, C => 
                           n114_port, D => n115_port, E => n116_port, F => 
                           n117_port, Z => n108_port);
   U520 : HS65_LH_AOI222X2 port map( A => N140, B => n51, C => n14, D => 
                           HI_LO_c_HI_9_port, E => n11, F => n79, Z => 
                           n109_port);
   U521 : HS65_LH_NAND4ABX3 port map( A => n424, B => n425, C => n426, D => 
                           n427, Z => alu_o(10));
   U522 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n335, D1 => n580, S1 
                           => n156_port, D2 => n79, S2 => n428, D3 => alu_i(52)
                           , S3 => n429, Z => n424);
   U523 : HS65_LH_AO222X4 port map( A => n290, B => n113_port, C => n157_port, 
                           D => n115_port, E => n291, F => n117_port, Z => n425
                           );
   U524 : HS65_LH_AOI222X2 port map( A => N141, B => n52, C => n15, D => 
                           HI_LO_c_HI_10_port, E => n12, F => alu_i(21), Z => 
                           n426);
   U525 : HS65_LH_NAND4ABX3 port map( A => n417, B => n418, C => n419, D => 
                           n420, Z => alu_o(11));
   U526 : HS65_LH_AO222X4 port map( A => n145_port, B => n115_port, C => n325, 
                           D => n118_port, E => n276, F => n113_port, Z => n418
                           );
   U527 : HS65_LH_OAI212X5 port map( A => n421, B => n80, C => n569, D => 
                           n176_port, E => n422, Z => n417);
   U528 : HS65_LH_AOI222X2 port map( A => N142, B => n52, C => n15, D => 
                           HI_LO_c_HI_11_port, E => n12, F => n81, Z => n419);
   U529 : HS65_LH_NAND4ABX3 port map( A => n411, B => n412, C => n413, D => 
                           n414, Z => alu_o(12));
   U530 : HS65_LH_MX41X7 port map( D0 => n580, S0 => n132_port, D1 => n81, S1 
                           => n415, D2 => n397, S2 => n263, D3 => alu_i(54), S3
                           => n416, Z => n411);
   U531 : HS65_LH_AO222X4 port map( A => n133_port, B => n115_port, C => n313, 
                           D => n118_port, E => n573, F => n113_port, Z => n412
                           );
   U532 : HS65_LH_AOI222X2 port map( A => N143, B => n52, C => n15, D => 
                           HI_LO_c_HI_12_port, E => n12, F => n82, Z => n413);
   U533 : HS65_LH_NAND4ABX3 port map( A => n405, B => n406, C => n407, D => 
                           n408, Z => alu_o(13));
   U534 : HS65_LH_MX41X7 port map( D0 => n580, S0 => n119_port, D1 => n82, S1 
                           => n409, D2 => n397, S2 => n247, D3 => alu_i(55), S3
                           => n410, Z => n405);
   U535 : HS65_LH_AO222X4 port map( A => n120_port, B => n115_port, C => n299, 
                           D => n118_port, E => n252, F => n113_port, Z => n406
                           );
   U536 : HS65_LH_AOI222X2 port map( A => N144, B => n52, C => n15, D => 
                           HI_LO_c_HI_13_port, E => n12, F => n83, Z => n407);
   U537 : HS65_LH_NAND4ABX3 port map( A => n399, B => n400, C => n401, D => 
                           n402, Z => alu_o(14));
   U538 : HS65_LH_MX41X7 port map( D0 => n580, S0 => n335, D1 => n83, S1 => 
                           n403, D2 => n397, S2 => n222_port, D3 => alu_i(56), 
                           S3 => n404, Z => n399);
   U539 : HS65_LH_AO222X4 port map( A => n156_port, B => n115_port, C => n334, 
                           D => n118_port, E => n227, F => n113_port, Z => n400
                           );
   U540 : HS65_LH_AOI222X2 port map( A => N145, B => n52, C => n15, D => 
                           HI_LO_c_HI_14_port, E => n12, F => n84, Z => n401);
   U541 : HS65_LH_NAND4ABX3 port map( A => n392, B => n393, C => n394, D => 
                           n395, Z => alu_o(15));
   U542 : HS65_LH_MX41X7 port map( D0 => n580, S0 => n325, D1 => n84, S1 => 
                           n396, D2 => n397, S2 => n216_port, D3 => alu_i(57), 
                           S3 => n398, Z => n392);
   U543 : HS65_LH_AO222X4 port map( A => n144_port, B => n115_port, C => n324, 
                           D => n118_port, E => n210_port, F => n113_port, Z =>
                           n393);
   U544 : HS65_LH_AOI222X2 port map( A => N146, B => n52, C => n15, D => 
                           HI_LO_c_HI_15_port, E => n12, F => n85, Z => n394);
   U545 : HS65_LH_AO222X4 port map( A => N649, B => n103_port, C => n16, D => 
                           HI_LO_c_HI_0_port, E => N648, F => n102_port, Z => 
                           n433);
   U546 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_29_port, B => n45, C => n82
                           , D => n106_port, E => HI_LO_c_HI_29_port, F => n16,
                           Z => n246);
   U547 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_30_port, B => n105_port, C 
                           => n83, D => n106_port, E => HI_LO_c_HI_30_port, F 
                           => n16, Z => n221_port);
   U548 : HS65_LH_IVX9 port map( A => alu_i(9), Z => n578);
   U549 : HS65_LH_AO212X4 port map( A => n173_port, B => n591, C => n387, D => 
                           alu_i(4), E => n446, Z => n444);
   U550 : HS65_LH_AO222X4 port map( A => n192_port, B => n130_port, C => 
                           n193_port, D => n447, E => n195_port, F => n128_port
                           , Z => n446);
   U551 : HS65_LH_AO212X4 port map( A => n27, B => alu_i(12), C => n35, D => 
                           n70, E => n449, Z => n447);
   U552 : HS65_LH_AO12X9 port map( A => alu_i(13), B => n21, C => n315, Z => 
                           n449);
   U553 : HS65_LH_AO212X4 port map( A => n164_port, B => n591, C => n360, D => 
                           alu_i(4), E => n361, Z => n359);
   U554 : HS65_LH_AO222X4 port map( A => n192_port, B => n114_port, C => 
                           n193_port, D => n362, E => n195_port, F => n111_port
                           , Z => n361);
   U555 : HS65_LH_MX41X7 port map( D0 => n70, S0 => n37, D1 => alu_i(12), S1 =>
                           n33, D2 => alu_i(13), S2 => n28, D3 => alu_i(14), S3
                           => n22, Z => n362);
   U556 : HS65_LH_AO212X4 port map( A => n251, B => n591, C => n252, D => 
                           alu_i(4), E => n253, Z => n250);
   U557 : HS65_LH_AO222X4 port map( A => n192_port, B => n254, C => n193_port, 
                           D => n255, E => n195_port, F => n256, Z => n253);
   U558 : HS65_LH_MX41X7 port map( D0 => n523, S0 => n196_port, D1 => alu_i(38)
                           , S1 => n32, D2 => alu_i(37), S2 => n27, D3 => n520,
                           S3 => n21, Z => n255);
   U559 : HS65_LH_AO212X4 port map( A => n226_port, B => n591, C => n227, D => 
                           alu_i(4), E => n228, Z => n225_port);
   U560 : HS65_LH_AO222X4 port map( A => n192_port, B => n229, C => n193_port, 
                           D => n230, E => n195_port, F => n231, Z => n228);
   U561 : HS65_LH_MX41X7 port map( D0 => n524, S0 => n37, D1 => n523, S1 => n32
                           , D2 => alu_i(38), S2 => n27, D3 => alu_i(37), S3 =>
                           n21, Z => n230);
   U562 : HS65_LH_NAND3X5 port map( A => n430, B => n431, C => n432, Z => 
                           alu_o(0));
   U563 : HS65_LH_AOI22X6 port map( A => n581, B => n444, C => n45, D => 
                           HI_LO_c_LO_0_port, Z => n430);
   U564 : HS65_LH_AOI212X4 port map( A => n13, B => n70, C => N131, D => n53, E
                           => n433, Z => n432);
   U565 : HS65_LH_AOI212X4 port map( A => N99, B => n48, C => n69, D => n439, E
                           => n440, Z => n431);
   U566 : HS65_LH_BFX9 port map( A => n196_port, Z => n36);
   U567 : HS65_LH_NOR2X6 port map( A => alu_i(0), B => alu_i(1), Z => n196_port
                           );
   U568 : HS65_LH_AO212X4 port map( A => n152_port, B => n591, C => n239, D => 
                           alu_i(4), E => n240, Z => n234);
   U569 : HS65_LH_AO222X4 port map( A => n192_port, B => n157_port, C => 
                           n193_port, D => n241, E => n195_port, F => n154_port
                           , Z => n240);
   U570 : HS65_LH_MX41X7 port map( D0 => alu_i(12), S0 => n36, D1 => alu_i(13),
                           S1 => n32, D2 => alu_i(14), S2 => n27, D3 => n74, S3
                           => n21, Z => n241);
   U571 : HS65_LH_AO212X4 port map( A => n209_port, B => n591, C => n210_port, 
                           D => alu_i(4), E => n211_port, Z => n203_port);
   U572 : HS65_LH_AO222X4 port map( A => n192_port, B => n212_port, C => 
                           n193_port, D => n213_port, E => n195_port, F => 
                           n214_port, Z => n211_port);
   U573 : HS65_LH_AO212X4 port map( A => n27, B => n523, C => n35, D => n524, E
                           => n215_port, Z => n213_port);
   U574 : HS65_LH_AO12X9 port map( A => alu_i(38), B => n21, C => n216_port, Z 
                           => n215_port);
   U575 : HS65_LH_BFX9 port map( A => alu_i(10), Z => n69);
   U576 : HS65_LH_IVX9 port map( A => alu_i(6), Z => n588);
   U577 : HS65_LH_IVX9 port map( A => alu_i(5), Z => n590);
   U578 : HS65_LH_IVX9 port map( A => alu_i(8), Z => n587);
   U579 : HS65_LH_IVX9 port map( A => alu_i(41), Z => n525);
   U580 : HS65_LH_IVX9 port map( A => alu_i(12), Z => n71);
   U581 : HS65_LH_IVX9 port map( A => alu_i(13), Z => n72);
   U582 : HS65_LH_IVX9 port map( A => alu_i(38), Z => n522);
   U583 : HS65_LH_IVX9 port map( A => alu_i(71), Z => n535);
   U584 : HS65_LH_BFX9 port map( A => n104_port, Z => n46);
   U585 : HS65_LH_OAI21X3 port map( A => alu_i(5), B => n437, C => n443, Z => 
                           n104_port);
   U586 : HS65_LH_OAI21X3 port map( A => n436, B => n435, C => n390, Z => n443)
                           ;
   U587 : HS65_LH_BFX9 port map( A => n198_port, Z => n26);
   U588 : HS65_LH_NOR2AX3 port map( A => alu_i(1), B => alu_i(0), Z => 
                           n198_port);
   U589 : HS65_LH_IVX9 port map( A => alu_i(14), Z => n73);
   U590 : HS65_LH_IVX9 port map( A => alu_i(21), Z => n80);
   U591 : HS65_LH_IVX9 port map( A => alu_i(30), Z => n89);
   U592 : HS65_LH_IVX9 port map( A => alu_i(37), Z => n521);
   U593 : HS65_LH_IVX9 port map( A => alu_i(47), Z => n527);
   U594 : HS65_LH_IVX9 port map( A => alu_i(50), Z => n528);
   U595 : HS65_LH_IVX9 port map( A => alu_i(56), Z => n530);
   U596 : HS65_LH_IVX9 port map( A => alu_i(59), Z => n531);
   U597 : HS65_LH_IVX9 port map( A => alu_i(65), Z => n533);
   U598 : HS65_LH_IVX9 port map( A => alu_i(68), Z => n534);
   U599 : HS65_LH_IVX9 port map( A => alu_i(44), Z => n526);
   U600 : HS65_LH_IVX9 port map( A => alu_i(53), Z => n529);
   U601 : HS65_LH_IVX9 port map( A => alu_i(62), Z => n532);
   U602 : HS65_LH_BFX9 port map( A => rst_n, Z => n537);
   U603 : HS65_LH_BFX9 port map( A => rst_n, Z => n536);
   U604 : HS65_LH_AO112X9 port map( A => N714, B => n450, C => n451, D => n452,
                           Z => alu_o(32));
   U605 : HS65_LH_AO222X4 port map( A => n391, B => n450, C => n438, D => n450,
                           E => n436, F => n450, Z => n452);
   U606 : HS65_LH_NOR4ABX2 port map( A => N715, B => n587, C => n578, D => n589
                           , Z => n451);
   U607 : HS65_LH_NOR3X4 port map( A => alu_i(7), B => alu_i(8), C => n578, Z 
                           => n450);
   U608 : HS65_LH_NAND2X7 port map( A => n257, B => n258, Z => alu_o(28));
   U609 : HS65_LH_AOI212X4 port map( A => n12, B => n523, C => N159, D => n53, 
                           E => n270, Z => n257);
   U610 : HS65_LH_AOI212X4 port map( A => N127, B => n48, C => n584, D => n259,
                           E => n260, Z => n258);
   U611 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_28_port, B => n45, C => n81
                           , D => n106_port, E => HI_LO_c_HI_28_port, F => n16,
                           Z => n270);
   U612 : HS65_LH_NAND2X7 port map( A => n201_port, B => n202_port, Z => 
                           alu_o(31));
   U613 : HS65_LH_AOI212X4 port map( A => n16, B => HI_LO_c_HI_31_port, C => 
                           N162, D => n53, E => n217_port, Z => n201_port);
   U614 : HS65_LH_AOI212X4 port map( A => N130, B => n48, C => n584, D => 
                           n203_port, E => n204_port, Z => n202_port);
   U615 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_31_port, B => n45, C => n84,
                           D => n106_port, Z => n217_port);
   U616 : HS65_LH_NAND2X7 port map( A => n232, B => n233, Z => alu_o(2));
   U617 : HS65_LH_AOI212X4 port map( A => n13, B => alu_i(13), C => N133, D => 
                           n53, E => n242, Z => n232);
   U618 : HS65_LH_AOI212X4 port map( A => N101, B => n48, C => n581, D => n234,
                           E => n235, Z => n233);
   U619 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_2_port, B => n16, C => 
                           HI_LO_c_LO_2_port, D => n45, Z => n242);
   U620 : HS65_LH_NAND2X7 port map( A => n181_port, B => n182_port, Z => 
                           alu_o(3));
   U621 : HS65_LH_AOI212X4 port map( A => n13, B => alu_i(14), C => N134, D => 
                           n53, E => n200_port, Z => n181_port);
   U622 : HS65_LH_AOI212X4 port map( A => N102, B => n48, C => n581, D => 
                           n183_port, E => n184_port, Z => n182_port);
   U623 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_3_port, B => n16, C => 
                           HI_LO_c_LO_3_port, D => n45, Z => n200_port);
   U624 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_1_port, B => n16, C => 
                           HI_LO_c_LO_1_port, D => n45, Z => n356);
   U625 : HS65_LH_IVX9 port map( A => alu_i(42), Z => n565);
   U626 : HS65_LH_IVX9 port map( A => alu_i(43), Z => n564);
   U627 : HS65_LH_IVX9 port map( A => alu_i(72), Z => n545);
   U628 : HS65_LH_IVX9 port map( A => alu_i(45), Z => n563);
   U629 : HS65_LH_IVX9 port map( A => alu_i(70), Z => n546);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_top is

   port( clk, rst_n : in std_logic;  src_a, src_b : in std_logic_vector (31 
         downto 0);  op, shamt : in std_logic_vector (4 downto 0);  result : 
         out std_logic_vector (31 downto 0);  branch : out std_logic);

end alu_top;

architecture SYN_Behavioral of alu_top is

   component alu
      port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 
            0);  alu_o : out std_logic_vector (32 downto 0));
   end component;

begin
   
   alu_inst : alu port map( clk => clk, rst_n => rst_n, alu_i(73) => src_a(31),
                           alu_i(72) => src_a(30), alu_i(71) => src_a(29), 
                           alu_i(70) => src_a(28), alu_i(69) => src_a(27), 
                           alu_i(68) => src_a(26), alu_i(67) => src_a(25), 
                           alu_i(66) => src_a(24), alu_i(65) => src_a(23), 
                           alu_i(64) => src_a(22), alu_i(63) => src_a(21), 
                           alu_i(62) => src_a(20), alu_i(61) => src_a(19), 
                           alu_i(60) => src_a(18), alu_i(59) => src_a(17), 
                           alu_i(58) => src_a(16), alu_i(57) => src_a(15), 
                           alu_i(56) => src_a(14), alu_i(55) => src_a(13), 
                           alu_i(54) => src_a(12), alu_i(53) => src_a(11), 
                           alu_i(52) => src_a(10), alu_i(51) => src_a(9), 
                           alu_i(50) => src_a(8), alu_i(49) => src_a(7), 
                           alu_i(48) => src_a(6), alu_i(47) => src_a(5), 
                           alu_i(46) => src_a(4), alu_i(45) => src_a(3), 
                           alu_i(44) => src_a(2), alu_i(43) => src_a(1), 
                           alu_i(42) => src_a(0), alu_i(41) => src_b(31), 
                           alu_i(40) => src_b(30), alu_i(39) => src_b(29), 
                           alu_i(38) => src_b(28), alu_i(37) => src_b(27), 
                           alu_i(36) => src_b(26), alu_i(35) => src_b(25), 
                           alu_i(34) => src_b(24), alu_i(33) => src_b(23), 
                           alu_i(32) => src_b(22), alu_i(31) => src_b(21), 
                           alu_i(30) => src_b(20), alu_i(29) => src_b(19), 
                           alu_i(28) => src_b(18), alu_i(27) => src_b(17), 
                           alu_i(26) => src_b(16), alu_i(25) => src_b(15), 
                           alu_i(24) => src_b(14), alu_i(23) => src_b(13), 
                           alu_i(22) => src_b(12), alu_i(21) => src_b(11), 
                           alu_i(20) => src_b(10), alu_i(19) => src_b(9), 
                           alu_i(18) => src_b(8), alu_i(17) => src_b(7), 
                           alu_i(16) => src_b(6), alu_i(15) => src_b(5), 
                           alu_i(14) => src_b(4), alu_i(13) => src_b(3), 
                           alu_i(12) => src_b(2), alu_i(11) => src_b(1), 
                           alu_i(10) => src_b(0), alu_i(9) => op(4), alu_i(8) 
                           => op(3), alu_i(7) => op(2), alu_i(6) => op(1), 
                           alu_i(5) => op(0), alu_i(4) => shamt(4), alu_i(3) =>
                           shamt(3), alu_i(2) => shamt(2), alu_i(1) => shamt(1)
                           , alu_i(0) => shamt(0), alu_o(32) => branch, 
                           alu_o(31) => result(31), alu_o(30) => result(30), 
                           alu_o(29) => result(29), alu_o(28) => result(28), 
                           alu_o(27) => result(27), alu_o(26) => result(26), 
                           alu_o(25) => result(25), alu_o(24) => result(24), 
                           alu_o(23) => result(23), alu_o(22) => result(22), 
                           alu_o(21) => result(21), alu_o(20) => result(20), 
                           alu_o(19) => result(19), alu_o(18) => result(18), 
                           alu_o(17) => result(17), alu_o(16) => result(16), 
                           alu_o(15) => result(15), alu_o(14) => result(14), 
                           alu_o(13) => result(13), alu_o(12) => result(12), 
                           alu_o(11) => result(11), alu_o(10) => result(10), 
                           alu_o(9) => result(9), alu_o(8) => result(8), 
                           alu_o(7) => result(7), alu_o(6) => result(6), 
                           alu_o(5) => result(5), alu_o(4) => result(4), 
                           alu_o(3) => result(3), alu_o(2) => result(2), 
                           alu_o(1) => result(1), alu_o(0) => result(0));

end SYN_Behavioral;
