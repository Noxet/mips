
module alu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328;

  HS65_LH_IVX9 U157 ( .A(n305), .Z(n256) );
  HS65_LH_OR2X9 U158 ( .A(B[11]), .B(n241), .Z(n327) );
  HS65_LH_IVX9 U159 ( .A(n316), .Z(n266) );
  HS65_LH_IVX9 U160 ( .A(B[3]), .Z(n228) );
  HS65_LH_IVX9 U161 ( .A(B[4]), .Z(n229) );
  HS65_LH_IVX9 U162 ( .A(A[17]), .Z(n243) );
  HS65_LH_IVX9 U163 ( .A(A[11]), .Z(n241) );
  HS65_LH_IVX9 U164 ( .A(B[27]), .Z(n237) );
  HS65_LH_IVX9 U165 ( .A(B[2]), .Z(n227) );
  HS65_LH_IVX9 U166 ( .A(A[14]), .Z(n242) );
  HS65_LH_IVX9 U167 ( .A(A[8]), .Z(n240) );
  HS65_LH_IVX9 U168 ( .A(A[20]), .Z(n244) );
  HS65_LH_IVX9 U169 ( .A(A[5]), .Z(n239) );
  HS65_LH_IVX9 U170 ( .A(A[29]), .Z(n245) );
  HS65_LH_IVX9 U171 ( .A(n321), .Z(n257) );
  HS65_LH_IVX9 U172 ( .A(n306), .Z(n260) );
  HS65_LH_IVX9 U173 ( .A(n296), .Z(n247) );
  HS65_LH_OR2X9 U174 ( .A(B[17]), .B(n243), .Z(n281) );
  HS65_LH_IVX9 U175 ( .A(n279), .Z(n252) );
  HS65_LH_IVX9 U176 ( .A(n297), .Z(n246) );
  HS65_LH_IVX9 U177 ( .A(n284), .Z(n250) );
  HS65_LH_IVX9 U178 ( .A(n320), .Z(n254) );
  HS65_LH_IVX9 U179 ( .A(n308), .Z(n263) );
  HS65_LH_IVX9 U180 ( .A(B[1]), .Z(n226) );
  HS65_LH_IVX9 U181 ( .A(B[23]), .Z(n233) );
  HS65_LH_IVX9 U182 ( .A(B[19]), .Z(n231) );
  HS65_LH_IVX9 U183 ( .A(B[26]), .Z(n236) );
  HS65_LH_IVX9 U184 ( .A(B[22]), .Z(n232) );
  HS65_LH_IVX9 U185 ( .A(B[18]), .Z(n230) );
  HS65_LH_IVX9 U186 ( .A(B[24]), .Z(n234) );
  HS65_LH_IVX9 U187 ( .A(B[30]), .Z(n238) );
  HS65_LH_IVX9 U188 ( .A(A[15]), .Z(n255) );
  HS65_LH_IVX9 U189 ( .A(A[7]), .Z(n264) );
  HS65_LH_IVX9 U190 ( .A(A[1]), .Z(n268) );
  HS65_LH_IVX9 U191 ( .A(B[25]), .Z(n235) );
  HS65_LH_AND2X4 U192 ( .A(A[3]), .B(n228), .Z(n318) );
  HS65_LH_IVX9 U193 ( .A(A[9]), .Z(n262) );
  HS65_LH_IVX9 U194 ( .A(A[31]), .Z(n248) );
  HS65_LH_IVX9 U195 ( .A(A[21]), .Z(n251) );
  HS65_LH_IVX9 U196 ( .A(A[16]), .Z(n253) );
  HS65_LH_IVX9 U197 ( .A(A[13]), .Z(n258) );
  HS65_LH_IVX9 U198 ( .A(A[12]), .Z(n259) );
  HS65_LH_IVX9 U199 ( .A(A[28]), .Z(n249) );
  HS65_LH_IVX9 U200 ( .A(A[6]), .Z(n265) );
  HS65_LH_IVX9 U201 ( .A(A[10]), .Z(n261) );
  HS65_LH_IVX9 U202 ( .A(A[4]), .Z(n267) );
  HS65_LH_OAI12X2 U203 ( .A(n269), .B(n270), .C(n271), .Z(GE_LT_GT_LE) );
  HS65_LH_OAI32X2 U204 ( .A(n272), .B(n273), .C(n274), .D(n275), .E(n272), .Z(
        n271) );
  HS65_LH_AOI212X2 U205 ( .A(n276), .B(n277), .C(n277), .D(n252), .E(n278), 
        .Z(n274) );
  HS65_LH_OA32X4 U206 ( .A(n230), .B(A[18]), .C(n280), .D(A[19]), .E(n231), 
        .Z(n277) );
  HS65_LH_AOI32X3 U207 ( .A(n281), .B(n253), .C(B[16]), .D(B[17]), .E(n243), 
        .Z(n276) );
  HS65_LH_AOI22X1 U208 ( .A(n282), .B(n283), .C(n283), .D(n250), .Z(n273) );
  HS65_LH_OA32X4 U209 ( .A(n232), .B(A[22]), .C(n285), .D(A[23]), .E(n233), 
        .Z(n283) );
  HS65_LH_AOI32X3 U210 ( .A(n286), .B(n244), .C(B[20]), .D(B[21]), .E(n251), 
        .Z(n282) );
  HS65_LH_CBI4I1X3 U211 ( .A(n247), .B(n246), .C(n287), .D(n288), .Z(n272) );
  HS65_LH_OAI212X3 U212 ( .A(n289), .B(n290), .C(n291), .D(n289), .E(n292), 
        .Z(n288) );
  HS65_LH_OAI32X2 U213 ( .A(n234), .B(A[24]), .C(n293), .D(A[25]), .E(n235), 
        .Z(n290) );
  HS65_LH_OAI32X2 U214 ( .A(n236), .B(A[26]), .C(n294), .D(A[27]), .E(n237), 
        .Z(n289) );
  HS65_LH_AOI312X2 U215 ( .A(n295), .B(n249), .C(B[28]), .D(B[29]), .E(n245), 
        .F(n296), .Z(n287) );
  HS65_LH_OAI32X2 U216 ( .A(n238), .B(A[30]), .C(n298), .D(B[31]), .E(n248), 
        .Z(n296) );
  HS65_LH_NAND3AX3 U217 ( .A(n278), .B(n279), .C(n275), .Z(n270) );
  HS65_LH_AND3X4 U218 ( .A(n291), .B(n292), .C(n299), .Z(n275) );
  HS65_LH_AOI12X2 U219 ( .A(A[24]), .B(n234), .C(n293), .Z(n299) );
  HS65_LH_NOR2AX3 U220 ( .A(A[25]), .B(B[25]), .Z(n293) );
  HS65_LH_OA112X4 U221 ( .A(B[28]), .B(n249), .C(n295), .D(n297), .Z(n292) );
  HS65_LH_AOI12X2 U222 ( .A(n238), .B(A[30]), .C(n298), .Z(n297) );
  HS65_LH_AND2X4 U223 ( .A(B[31]), .B(n248), .Z(n298) );
  HS65_LH_OR2X4 U224 ( .A(B[29]), .B(n245), .Z(n295) );
  HS65_LH_AOI12X2 U225 ( .A(n236), .B(A[26]), .C(n294), .Z(n291) );
  HS65_LH_AND2X4 U226 ( .A(A[27]), .B(n237), .Z(n294) );
  HS65_LH_AOI12X2 U227 ( .A(n230), .B(A[18]), .C(n280), .Z(n279) );
  HS65_LH_AND2X4 U228 ( .A(A[19]), .B(n231), .Z(n280) );
  HS65_LH_OAI112X1 U229 ( .A(B[20]), .B(n244), .C(n286), .D(n284), .Z(n278) );
  HS65_LH_AOI12X2 U230 ( .A(n232), .B(A[22]), .C(n285), .Z(n284) );
  HS65_LH_AND2X4 U231 ( .A(A[23]), .B(n233), .Z(n285) );
  HS65_LH_OR2X4 U232 ( .A(B[21]), .B(n251), .Z(n286) );
  HS65_LH_OAI212X3 U233 ( .A(n300), .B(n301), .C(n302), .D(n300), .E(n303), 
        .Z(n269) );
  HS65_LH_OA12X4 U234 ( .A(n253), .B(B[16]), .C(n281), .Z(n303) );
  HS65_LH_NOR3X1 U235 ( .A(n304), .B(n305), .C(n306), .Z(n302) );
  HS65_LH_OAI12X2 U236 ( .A(B[8]), .B(n240), .C(n307), .Z(n304) );
  HS65_LH_CBI4I1X3 U237 ( .A(n308), .B(n309), .C(n310), .D(n311), .Z(n301) );
  HS65_LH_NAND3AX3 U238 ( .A(n309), .B(n312), .C(n313), .Z(n311) );
  HS65_LH_AOI212X2 U239 ( .A(n314), .B(n315), .C(A[4]), .D(n229), .E(n316), 
        .Z(n313) );
  HS65_LH_AOI22X1 U240 ( .A(B[1]), .B(n268), .C(n317), .D(B[0]), .Z(n314) );
  HS65_LH_AOI12X2 U241 ( .A(A[1]), .B(n226), .C(A[0]), .Z(n317) );
  HS65_LH_CBI4I1X3 U242 ( .A(A[2]), .B(n227), .C(n318), .D(n315), .Z(n312) );
  HS65_LH_OA32X4 U243 ( .A(n227), .B(A[2]), .C(n318), .D(A[3]), .E(n228), .Z(
        n315) );
  HS65_LH_AOI312X2 U244 ( .A(n266), .B(n267), .C(B[4]), .D(B[5]), .E(n239), 
        .F(n263), .Z(n310) );
  HS65_LH_NOR2X2 U245 ( .A(n239), .B(B[5]), .Z(n316) );
  HS65_LH_OAI12X2 U246 ( .A(B[6]), .B(n265), .C(n319), .Z(n309) );
  HS65_LH_AOI32X3 U247 ( .A(B[6]), .B(n265), .C(n319), .D(n264), .E(B[7]), .Z(
        n308) );
  HS65_LH_NAND2AX4 U248 ( .A(B[7]), .B(A[7]), .Z(n319) );
  HS65_LH_CBI4I1X3 U249 ( .A(n320), .B(n321), .C(n322), .D(n323), .Z(n300) );
  HS65_LH_OAI212X3 U250 ( .A(n324), .B(n325), .C(n260), .D(n324), .E(n256), 
        .Z(n323) );
  HS65_LH_OAI112X1 U251 ( .A(B[12]), .B(n259), .C(n326), .D(n257), .Z(n305) );
  HS65_LH_OAI12X2 U252 ( .A(B[10]), .B(n261), .C(n327), .Z(n306) );
  HS65_LH_AO32X4 U253 ( .A(B[8]), .B(n240), .C(n307), .D(n262), .E(B[9]), .Z(
        n325) );
  HS65_LH_NAND2AX4 U254 ( .A(B[9]), .B(A[9]), .Z(n307) );
  HS65_LH_AO32X4 U255 ( .A(B[10]), .B(n261), .C(n327), .D(n241), .E(B[11]), 
        .Z(n324) );
  HS65_LH_AOI312X2 U256 ( .A(n326), .B(n259), .C(B[12]), .D(B[13]), .E(n258), 
        .F(n254), .Z(n322) );
  HS65_LH_OR2X4 U257 ( .A(B[13]), .B(n258), .Z(n326) );
  HS65_LH_OAI12X2 U258 ( .A(B[14]), .B(n242), .C(n328), .Z(n321) );
  HS65_LH_AOI32X3 U259 ( .A(B[14]), .B(n242), .C(n328), .D(n255), .E(B[15]), 
        .Z(n320) );
  HS65_LH_NAND2AX4 U260 ( .A(B[15]), .B(A[15]), .Z(n328) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  HS65_LHS_XOR3X2 U2_31 ( .A(A[31]), .B(n33), .C(carry[31]), .Z(DIFF[31]) );
  HS65_LH_FA1X4 U2_30 ( .A0(A[30]), .B0(n32), .CI(carry[30]), .CO(carry[31]), 
        .S0(DIFF[30]) );
  HS65_LH_FA1X4 U2_28 ( .A0(A[28]), .B0(n30), .CI(carry[28]), .CO(carry[29]), 
        .S0(DIFF[28]) );
  HS65_LH_FA1X4 U2_27 ( .A0(A[27]), .B0(n29), .CI(carry[27]), .CO(carry[28]), 
        .S0(DIFF[27]) );
  HS65_LH_FA1X4 U2_25 ( .A0(A[25]), .B0(n27), .CI(carry[25]), .CO(carry[26]), 
        .S0(DIFF[25]) );
  HS65_LH_FA1X4 U2_24 ( .A0(A[24]), .B0(n26), .CI(carry[24]), .CO(carry[25]), 
        .S0(DIFF[24]) );
  HS65_LH_FA1X4 U2_22 ( .A0(A[22]), .B0(n24), .CI(carry[22]), .CO(carry[23]), 
        .S0(DIFF[22]) );
  HS65_LH_FA1X4 U2_21 ( .A0(A[21]), .B0(n23), .CI(carry[21]), .CO(carry[22]), 
        .S0(DIFF[21]) );
  HS65_LH_FA1X4 U2_19 ( .A0(A[19]), .B0(n21), .CI(carry[19]), .CO(carry[20]), 
        .S0(DIFF[19]) );
  HS65_LH_FA1X4 U2_18 ( .A0(A[18]), .B0(n20), .CI(carry[18]), .CO(carry[19]), 
        .S0(DIFF[18]) );
  HS65_LH_FA1X4 U2_16 ( .A0(A[16]), .B0(n18), .CI(carry[16]), .CO(carry[17]), 
        .S0(DIFF[16]) );
  HS65_LH_FA1X4 U2_15 ( .A0(A[15]), .B0(n17), .CI(carry[15]), .CO(carry[16]), 
        .S0(DIFF[15]) );
  HS65_LH_FA1X4 U2_13 ( .A0(A[13]), .B0(n15), .CI(carry[13]), .CO(carry[14]), 
        .S0(DIFF[13]) );
  HS65_LH_FA1X4 U2_12 ( .A0(A[12]), .B0(n14), .CI(carry[12]), .CO(carry[13]), 
        .S0(DIFF[12]) );
  HS65_LH_FA1X4 U2_10 ( .A0(A[10]), .B0(n12), .CI(carry[10]), .CO(carry[11]), 
        .S0(DIFF[10]) );
  HS65_LH_FA1X4 U2_9 ( .A0(A[9]), .B0(n11), .CI(carry[9]), .CO(carry[10]), 
        .S0(DIFF[9]) );
  HS65_LH_FA1X4 U2_7 ( .A0(A[7]), .B0(n9), .CI(carry[7]), .CO(carry[8]), .S0(
        DIFF[7]) );
  HS65_LH_FA1X4 U2_6 ( .A0(A[6]), .B0(n8), .CI(carry[6]), .CO(carry[7]), .S0(
        DIFF[6]) );
  HS65_LH_FA1X4 U2_4 ( .A0(A[4]), .B0(n6), .CI(carry[4]), .CO(carry[5]), .S0(
        DIFF[4]) );
  HS65_LH_FA1X4 U2_3 ( .A0(A[3]), .B0(n5), .CI(carry[3]), .CO(carry[4]), .S0(
        DIFF[3]) );
  HS65_LH_FA1X4 U2_1 ( .A0(A[1]), .B0(n3), .CI(carry[1]), .CO(carry[2]), .S0(
        DIFF[1]) );
  HS65_LH_FA1X4 U2_23 ( .A0(A[23]), .B0(n25), .CI(carry[23]), .CO(carry[24]), 
        .S0(DIFF[23]) );
  HS65_LH_FA1X4 U2_2 ( .A0(A[2]), .B0(n4), .CI(carry[2]), .CO(carry[3]), .S0(
        DIFF[2]) );
  HS65_LH_FA1X4 U2_29 ( .A0(A[29]), .B0(n31), .CI(carry[29]), .CO(carry[30]), 
        .S0(DIFF[29]) );
  HS65_LH_FA1X4 U2_26 ( .A0(A[26]), .B0(n28), .CI(carry[26]), .CO(carry[27]), 
        .S0(DIFF[26]) );
  HS65_LH_FA1X4 U2_20 ( .A0(A[20]), .B0(n22), .CI(carry[20]), .CO(carry[21]), 
        .S0(DIFF[20]) );
  HS65_LH_FA1X4 U2_17 ( .A0(A[17]), .B0(n19), .CI(carry[17]), .CO(carry[18]), 
        .S0(DIFF[17]) );
  HS65_LH_FA1X4 U2_11 ( .A0(A[11]), .B0(n13), .CI(carry[11]), .CO(carry[12]), 
        .S0(DIFF[11]) );
  HS65_LH_FA1X4 U2_5 ( .A0(A[5]), .B0(n7), .CI(carry[5]), .CO(carry[6]), .S0(
        DIFF[5]) );
  HS65_LH_FA1X4 U2_14 ( .A0(A[14]), .B0(n16), .CI(carry[14]), .CO(carry[15]), 
        .S0(DIFF[14]) );
  HS65_LH_FA1X4 U2_8 ( .A0(A[8]), .B0(n10), .CI(carry[8]), .CO(carry[9]), .S0(
        DIFF[8]) );
  HS65_LH_IVX9 U1 ( .A(B[8]), .Z(n10) );
  HS65_LH_IVX9 U2 ( .A(B[14]), .Z(n16) );
  HS65_LH_IVX9 U3 ( .A(B[5]), .Z(n7) );
  HS65_LH_IVX9 U4 ( .A(B[11]), .Z(n13) );
  HS65_LH_IVX9 U5 ( .A(B[17]), .Z(n19) );
  HS65_LH_IVX9 U6 ( .A(B[20]), .Z(n22) );
  HS65_LH_IVX9 U7 ( .A(B[26]), .Z(n28) );
  HS65_LH_IVX9 U8 ( .A(B[29]), .Z(n31) );
  HS65_LH_IVX9 U9 ( .A(B[2]), .Z(n4) );
  HS65_LH_IVX9 U10 ( .A(B[23]), .Z(n25) );
  HS65_LH_IVX9 U11 ( .A(B[0]), .Z(n2) );
  HS65_LHS_XNOR2X6 U12 ( .A(A[0]), .B(n2), .Z(DIFF[0]) );
  HS65_LH_IVX9 U13 ( .A(B[1]), .Z(n3) );
  HS65_LH_NAND2X7 U14 ( .A(n1), .B(B[0]), .Z(carry[1]) );
  HS65_LH_IVX9 U15 ( .A(A[0]), .Z(n1) );
  HS65_LH_IVX9 U16 ( .A(B[3]), .Z(n5) );
  HS65_LH_IVX9 U17 ( .A(B[4]), .Z(n6) );
  HS65_LH_IVX9 U18 ( .A(B[6]), .Z(n8) );
  HS65_LH_IVX9 U19 ( .A(B[7]), .Z(n9) );
  HS65_LH_IVX9 U20 ( .A(B[9]), .Z(n11) );
  HS65_LH_IVX9 U21 ( .A(B[10]), .Z(n12) );
  HS65_LH_IVX9 U22 ( .A(B[12]), .Z(n14) );
  HS65_LH_IVX9 U23 ( .A(B[13]), .Z(n15) );
  HS65_LH_IVX9 U24 ( .A(B[15]), .Z(n17) );
  HS65_LH_IVX9 U25 ( .A(B[16]), .Z(n18) );
  HS65_LH_IVX9 U26 ( .A(B[18]), .Z(n20) );
  HS65_LH_IVX9 U27 ( .A(B[19]), .Z(n21) );
  HS65_LH_IVX9 U28 ( .A(B[21]), .Z(n23) );
  HS65_LH_IVX9 U29 ( .A(B[22]), .Z(n24) );
  HS65_LH_IVX9 U30 ( .A(B[24]), .Z(n26) );
  HS65_LH_IVX9 U31 ( .A(B[25]), .Z(n27) );
  HS65_LH_IVX9 U32 ( .A(B[27]), .Z(n29) );
  HS65_LH_IVX9 U33 ( .A(B[28]), .Z(n30) );
  HS65_LH_IVX9 U34 ( .A(B[30]), .Z(n32) );
  HS65_LH_IVX9 U35 ( .A(B[31]), .Z(n33) );
endmodule


module alu_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115;

  HS65_LH_IVX9 U1 ( .A(n54), .Z(n35) );
  HS65_LH_IVX9 U2 ( .A(EQ), .Z(NE) );
  HS65_LH_IVX9 U3 ( .A(n115), .Z(n40) );
  HS65_LH_IVX9 U4 ( .A(A[14]), .Z(n21) );
  HS65_LH_IVX9 U5 ( .A(A[26]), .Z(n22) );
  HS65_LH_IVX9 U6 ( .A(B[2]), .Z(n1) );
  HS65_LH_IVX9 U7 ( .A(B[3]), .Z(n2) );
  HS65_LH_IVX9 U8 ( .A(B[27]), .Z(n16) );
  HS65_LH_IVX9 U9 ( .A(B[20]), .Z(n12) );
  HS65_LH_IVX9 U10 ( .A(B[11]), .Z(n6) );
  HS65_LH_IVX9 U11 ( .A(A[8]), .Z(n20) );
  HS65_LH_IVX9 U12 ( .A(B[28]), .Z(n17) );
  HS65_LH_IVX9 U13 ( .A(B[31]), .Z(n19) );
  HS65_LH_IVX9 U14 ( .A(n102), .Z(n38) );
  HS65_LH_IVX9 U15 ( .A(n67), .Z(n27) );
  HS65_LH_OR2X9 U16 ( .A(B[26]), .B(n22), .Z(n66) );
  HS65_LH_OR2X9 U17 ( .A(B[14]), .B(n21), .Z(n50) );
  HS65_LH_IVX9 U18 ( .A(B[23]), .Z(n14) );
  HS65_LH_IVX9 U19 ( .A(B[19]), .Z(n11) );
  HS65_LH_IVX9 U20 ( .A(B[25]), .Z(n15) );
  HS65_LH_IVX9 U21 ( .A(B[12]), .Z(n7) );
  HS65_LH_IVX9 U22 ( .A(B[13]), .Z(n8) );
  HS65_LH_IVX9 U23 ( .A(B[21]), .Z(n13) );
  HS65_LH_IVX9 U24 ( .A(B[15]), .Z(n9) );
  HS65_LH_IVX9 U25 ( .A(B[7]), .Z(n4) );
  HS65_LH_IVX9 U26 ( .A(B[5]), .Z(n3) );
  HS65_LH_IVX9 U27 ( .A(B[29]), .Z(n18) );
  HS65_LH_IVX9 U28 ( .A(B[9]), .Z(n5) );
  HS65_LH_IVX9 U29 ( .A(B[17]), .Z(n10) );
  HS65_LH_IVX9 U30 ( .A(n76), .Z(n24) );
  HS65_LH_IVX9 U31 ( .A(n60), .Z(n25) );
  HS65_LH_IVX9 U32 ( .A(n64), .Z(n28) );
  HS65_LH_IVX9 U33 ( .A(n51), .Z(n37) );
  HS65_LH_IVX9 U34 ( .A(A[22]), .Z(n30) );
  HS65_LH_IVX9 U35 ( .A(A[6]), .Z(n39) );
  HS65_LH_IVX9 U36 ( .A(n71), .Z(n33) );
  HS65_LH_IVX9 U37 ( .A(n70), .Z(n31) );
  HS65_LH_IVX9 U38 ( .A(A[1]), .Z(n42) );
  HS65_LH_IVX9 U39 ( .A(A[18]), .Z(n32) );
  HS65_LH_IVX9 U40 ( .A(A[4]), .Z(n41) );
  HS65_LH_IVX9 U41 ( .A(A[16]), .Z(n34) );
  HS65_LH_IVX9 U42 ( .A(A[24]), .Z(n29) );
  HS65_LH_IVX9 U43 ( .A(A[30]), .Z(n26) );
  HS65_LH_IVX9 U44 ( .A(A[10]), .Z(n36) );
  HS65_LH_NOR4ABX2 U45 ( .A(n43), .B(n44), .C(n45), .D(n46), .Z(EQ) );
  HS65_LH_NAND4X4 U46 ( .A(n47), .B(n48), .C(n49), .D(n50), .Z(n46) );
  HS65_LH_NAND4ABX3 U47 ( .A(n51), .B(n35), .C(n52), .D(n53), .Z(n45) );
  HS65_LH_NOR4ABX2 U48 ( .A(n55), .B(n56), .C(n57), .D(n58), .Z(n44) );
  HS65_LH_NAND4ABX3 U49 ( .A(n59), .B(n60), .C(n61), .D(n62), .Z(n58) );
  HS65_LH_AOI22X1 U50 ( .A(n42), .B(n63), .C(n63), .D(B[1]), .Z(n59) );
  HS65_LH_NAND2AX4 U51 ( .A(B[0]), .B(A[0]), .Z(n63) );
  HS65_LH_NAND4ABX3 U52 ( .A(n64), .B(n27), .C(n65), .D(n66), .Z(n57) );
  HS65_LH_NOR4ABX2 U53 ( .A(n68), .B(n69), .C(n70), .D(n71), .Z(n56) );
  HS65_LH_AND4X3 U54 ( .A(n72), .B(n73), .C(n74), .D(n75), .Z(n55) );
  HS65_LH_NOR4ABX2 U55 ( .A(n76), .B(n77), .C(n78), .D(LT), .Z(n43) );
  HS65_LH_OAI22X1 U56 ( .A(A[31]), .B(n19), .C(n24), .D(n79), .Z(LT) );
  HS65_LH_AOI32X3 U57 ( .A(n62), .B(n25), .C(n80), .D(B[30]), .E(n26), .Z(n79)
         );
  HS65_LH_OAI212X3 U58 ( .A(A[28]), .B(n17), .C(A[29]), .D(n18), .E(n81), .Z(
        n80) );
  HS65_LH_NAND3X2 U59 ( .A(n61), .B(n67), .C(n82), .Z(n81) );
  HS65_LH_OAI12X2 U60 ( .A(A[27]), .B(n16), .C(n83), .Z(n82) );
  HS65_LH_AOI32X3 U61 ( .A(n66), .B(n65), .C(n84), .D(B[26]), .E(n22), .Z(n83)
         );
  HS65_LH_OAI12X2 U62 ( .A(A[25]), .B(n15), .C(n85), .Z(n84) );
  HS65_LH_AOI32X3 U63 ( .A(n28), .B(n72), .C(n86), .D(B[24]), .E(n29), .Z(n85)
         );
  HS65_LH_OAI12X2 U64 ( .A(A[23]), .B(n14), .C(n87), .Z(n86) );
  HS65_LH_AOI32X3 U65 ( .A(n73), .B(n75), .C(n88), .D(B[22]), .E(n30), .Z(n87)
         );
  HS65_LH_OAI212X3 U66 ( .A(A[20]), .B(n12), .C(A[21]), .D(n13), .E(n89), .Z(
        n88) );
  HS65_LH_NAND3X2 U67 ( .A(n74), .B(n68), .C(n90), .Z(n89) );
  HS65_LH_OAI12X2 U68 ( .A(A[19]), .B(n11), .C(n91), .Z(n90) );
  HS65_LH_AOI32X3 U69 ( .A(n31), .B(n69), .C(n92), .D(B[18]), .E(n32), .Z(n91)
         );
  HS65_LH_OAI12X2 U70 ( .A(A[17]), .B(n10), .C(n93), .Z(n92) );
  HS65_LH_AOI32X3 U71 ( .A(n33), .B(n49), .C(n94), .D(B[16]), .E(n34), .Z(n93)
         );
  HS65_LH_OAI12X2 U72 ( .A(A[15]), .B(n9), .C(n95), .Z(n94) );
  HS65_LH_AOI32X3 U73 ( .A(n50), .B(n48), .C(n96), .D(B[14]), .E(n21), .Z(n95)
         );
  HS65_LH_OAI212X3 U74 ( .A(A[12]), .B(n7), .C(A[13]), .D(n8), .E(n97), .Z(n96) );
  HS65_LH_NAND3X2 U75 ( .A(n47), .B(n54), .C(n98), .Z(n97) );
  HS65_LH_OAI12X2 U76 ( .A(A[11]), .B(n6), .C(n99), .Z(n98) );
  HS65_LH_AOI32X3 U77 ( .A(n53), .B(n52), .C(n100), .D(B[10]), .E(n36), .Z(n99) );
  HS65_LH_OAI12X2 U78 ( .A(A[9]), .B(n5), .C(n101), .Z(n100) );
  HS65_LH_AOI32X3 U79 ( .A(n37), .B(n102), .C(n103), .D(B[8]), .E(n20), .Z(
        n101) );
  HS65_LH_OAI12X2 U80 ( .A(A[7]), .B(n4), .C(n104), .Z(n103) );
  HS65_LH_AOI32X3 U81 ( .A(n105), .B(n106), .C(n107), .D(B[6]), .E(n39), .Z(
        n104) );
  HS65_LH_OAI12X2 U82 ( .A(A[5]), .B(n3), .C(n108), .Z(n107) );
  HS65_LH_AOI32X3 U83 ( .A(n40), .B(n109), .C(n110), .D(B[4]), .E(n41), .Z(
        n108) );
  HS65_LH_OAI212X3 U84 ( .A(A[2]), .B(n1), .C(A[3]), .D(n2), .E(n111), .Z(n110) );
  HS65_LH_OAI212X3 U85 ( .A(B[1]), .B(n112), .C(n113), .D(n42), .E(n114), .Z(
        n111) );
  HS65_LH_AND2X4 U86 ( .A(n113), .B(n42), .Z(n112) );
  HS65_LH_NOR2AX3 U87 ( .A(B[0]), .B(A[0]), .Z(n113) );
  HS65_LH_NOR2X2 U88 ( .A(n20), .B(B[8]), .Z(n51) );
  HS65_LH_NAND2X2 U89 ( .A(A[9]), .B(n5), .Z(n52) );
  HS65_LH_NAND2AX4 U90 ( .A(B[10]), .B(A[10]), .Z(n53) );
  HS65_LH_NAND2X2 U91 ( .A(A[11]), .B(n6), .Z(n54) );
  HS65_LH_NAND2X2 U92 ( .A(A[12]), .B(n7), .Z(n47) );
  HS65_LH_NAND2X2 U93 ( .A(A[13]), .B(n8), .Z(n48) );
  HS65_LH_NAND2X2 U94 ( .A(A[15]), .B(n9), .Z(n49) );
  HS65_LH_NOR2X2 U95 ( .A(n34), .B(B[16]), .Z(n71) );
  HS65_LH_NAND2X2 U96 ( .A(A[17]), .B(n10), .Z(n69) );
  HS65_LH_NOR2X2 U97 ( .A(B[18]), .B(n32), .Z(n70) );
  HS65_LH_NAND2X2 U98 ( .A(A[19]), .B(n11), .Z(n68) );
  HS65_LH_NAND2X2 U99 ( .A(A[20]), .B(n12), .Z(n74) );
  HS65_LH_NAND2X2 U100 ( .A(A[21]), .B(n13), .Z(n75) );
  HS65_LH_NAND2AX4 U101 ( .A(B[22]), .B(A[22]), .Z(n73) );
  HS65_LH_NAND2X2 U102 ( .A(A[23]), .B(n14), .Z(n72) );
  HS65_LH_NOR2X2 U103 ( .A(n29), .B(B[24]), .Z(n64) );
  HS65_LH_NAND2X2 U104 ( .A(A[25]), .B(n15), .Z(n65) );
  HS65_LH_NAND2X2 U105 ( .A(A[27]), .B(n16), .Z(n67) );
  HS65_LH_NAND2X2 U106 ( .A(A[28]), .B(n17), .Z(n61) );
  HS65_LH_NOR2X2 U107 ( .A(n26), .B(B[30]), .Z(n60) );
  HS65_LH_NAND2X2 U108 ( .A(A[29]), .B(n18), .Z(n62) );
  HS65_LH_NAND4ABX3 U109 ( .A(n115), .B(n38), .C(n106), .D(n105), .Z(n78) );
  HS65_LH_NAND2AX4 U110 ( .A(B[6]), .B(A[6]), .Z(n105) );
  HS65_LH_NAND2X2 U111 ( .A(A[5]), .B(n3), .Z(n106) );
  HS65_LH_NAND2X2 U112 ( .A(A[7]), .B(n4), .Z(n102) );
  HS65_LH_NOR2X2 U113 ( .A(n41), .B(B[4]), .Z(n115) );
  HS65_LH_AND2X4 U114 ( .A(n114), .B(n109), .Z(n77) );
  HS65_LH_NAND2X2 U115 ( .A(A[3]), .B(n2), .Z(n109) );
  HS65_LH_NAND2X2 U116 ( .A(A[2]), .B(n1), .Z(n114) );
  HS65_LH_NAND2X2 U117 ( .A(A[31]), .B(n19), .Z(n76) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  HS65_LHS_XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Z(SUM[31]) );
  HS65_LH_FA1X4 U1_30 ( .A0(A[30]), .B0(B[30]), .CI(carry[30]), .CO(carry[31]), 
        .S0(SUM[30]) );
  HS65_LH_FA1X4 U1_28 ( .A0(A[28]), .B0(B[28]), .CI(carry[28]), .CO(carry[29]), 
        .S0(SUM[28]) );
  HS65_LH_FA1X4 U1_27 ( .A0(A[27]), .B0(B[27]), .CI(carry[27]), .CO(carry[28]), 
        .S0(SUM[27]) );
  HS65_LH_FA1X4 U1_25 ( .A0(A[25]), .B0(B[25]), .CI(carry[25]), .CO(carry[26]), 
        .S0(SUM[25]) );
  HS65_LH_FA1X4 U1_24 ( .A0(A[24]), .B0(B[24]), .CI(carry[24]), .CO(carry[25]), 
        .S0(SUM[24]) );
  HS65_LH_FA1X4 U1_22 ( .A0(A[22]), .B0(B[22]), .CI(carry[22]), .CO(carry[23]), 
        .S0(SUM[22]) );
  HS65_LH_FA1X4 U1_21 ( .A0(A[21]), .B0(B[21]), .CI(carry[21]), .CO(carry[22]), 
        .S0(SUM[21]) );
  HS65_LH_FA1X4 U1_19 ( .A0(A[19]), .B0(B[19]), .CI(carry[19]), .CO(carry[20]), 
        .S0(SUM[19]) );
  HS65_LH_FA1X4 U1_18 ( .A0(A[18]), .B0(B[18]), .CI(carry[18]), .CO(carry[19]), 
        .S0(SUM[18]) );
  HS65_LH_FA1X4 U1_16 ( .A0(A[16]), .B0(B[16]), .CI(carry[16]), .CO(carry[17]), 
        .S0(SUM[16]) );
  HS65_LH_FA1X4 U1_3 ( .A0(A[3]), .B0(B[3]), .CI(carry[3]), .CO(carry[4]), 
        .S0(SUM[3]) );
  HS65_LH_FA1X4 U1_1 ( .A0(A[1]), .B0(B[1]), .CI(n1), .CO(carry[2]), .S0(
        SUM[1]) );
  HS65_LH_FA1X4 U1_15 ( .A0(A[15]), .B0(B[15]), .CI(carry[15]), .CO(carry[16]), 
        .S0(SUM[15]) );
  HS65_LH_FA1X4 U1_13 ( .A0(A[13]), .B0(B[13]), .CI(carry[13]), .CO(carry[14]), 
        .S0(SUM[13]) );
  HS65_LH_FA1X4 U1_12 ( .A0(A[12]), .B0(B[12]), .CI(carry[12]), .CO(carry[13]), 
        .S0(SUM[12]) );
  HS65_LH_FA1X4 U1_10 ( .A0(A[10]), .B0(B[10]), .CI(carry[10]), .CO(carry[11]), 
        .S0(SUM[10]) );
  HS65_LH_FA1X4 U1_9 ( .A0(A[9]), .B0(B[9]), .CI(carry[9]), .CO(carry[10]), 
        .S0(SUM[9]) );
  HS65_LH_FA1X4 U1_7 ( .A0(A[7]), .B0(B[7]), .CI(carry[7]), .CO(carry[8]), 
        .S0(SUM[7]) );
  HS65_LH_FA1X4 U1_6 ( .A0(A[6]), .B0(B[6]), .CI(carry[6]), .CO(carry[7]), 
        .S0(SUM[6]) );
  HS65_LH_FA1X4 U1_4 ( .A0(A[4]), .B0(B[4]), .CI(carry[4]), .CO(carry[5]), 
        .S0(SUM[4]) );
  HS65_LH_FA1X4 U1_23 ( .A0(A[23]), .B0(B[23]), .CI(carry[23]), .CO(carry[24]), 
        .S0(SUM[23]) );
  HS65_LH_FA1X4 U1_2 ( .A0(A[2]), .B0(B[2]), .CI(carry[2]), .CO(carry[3]), 
        .S0(SUM[2]) );
  HS65_LH_FA1X4 U1_29 ( .A0(A[29]), .B0(B[29]), .CI(carry[29]), .CO(carry[30]), 
        .S0(SUM[29]) );
  HS65_LH_FA1X4 U1_26 ( .A0(A[26]), .B0(B[26]), .CI(carry[26]), .CO(carry[27]), 
        .S0(SUM[26]) );
  HS65_LH_FA1X4 U1_20 ( .A0(A[20]), .B0(B[20]), .CI(carry[20]), .CO(carry[21]), 
        .S0(SUM[20]) );
  HS65_LH_FA1X4 U1_17 ( .A0(A[17]), .B0(B[17]), .CI(carry[17]), .CO(carry[18]), 
        .S0(SUM[17]) );
  HS65_LH_FA1X4 U1_11 ( .A0(A[11]), .B0(B[11]), .CI(carry[11]), .CO(carry[12]), 
        .S0(SUM[11]) );
  HS65_LH_FA1X4 U1_5 ( .A0(A[5]), .B0(B[5]), .CI(carry[5]), .CO(carry[6]), 
        .S0(SUM[5]) );
  HS65_LH_FA1X4 U1_14 ( .A0(A[14]), .B0(B[14]), .CI(carry[14]), .CO(carry[15]), 
        .S0(SUM[14]) );
  HS65_LH_FA1X4 U1_8 ( .A0(A[8]), .B0(B[8]), .CI(carry[8]), .CO(carry[9]), 
        .S0(SUM[8]) );
  HS65_LH_AND2X4 U1 ( .A(A[0]), .B(B[0]), .Z(n1) );
  HS65_LHS_XOR2X6 U2 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
endmodule


module alu_DW_mult_uns_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n7, n19, n31, n43, n55, n67, n79, n91, n103, n115, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n292, n293, n294, n295, n296, n297,
         n299, n300, n302, n303, n304, n305, n306, n307, n308, n309, n311,
         n312, n313, n314, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
         n360, n361, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
  assign n7 = a[2];
  assign n19 = a[5];
  assign n31 = a[8];
  assign n43 = a[11];
  assign n55 = a[14];
  assign n67 = a[17];
  assign n79 = a[20];
  assign n91 = a[23];
  assign n103 = a[26];
  assign n115 = a[29];

  HS65_LH_FA1X4 U228 ( .A0(n293), .B0(n292), .CI(n228), .CO(n227), .S0(
        product[62]) );
  HS65_LH_FA1X4 U229 ( .A0(n295), .B0(n294), .CI(n229), .CO(n228), .S0(
        product[61]) );
  HS65_LH_FA1X4 U230 ( .A0(n296), .B0(n299), .CI(n230), .CO(n229), .S0(
        product[60]) );
  HS65_LH_FA1X4 U231 ( .A0(n300), .B0(n302), .CI(n231), .CO(n230), .S0(
        product[59]) );
  HS65_LH_FA1X4 U232 ( .A0(n303), .B0(n305), .CI(n232), .CO(n231), .S0(
        product[58]) );
  HS65_LH_FA1X4 U233 ( .A0(n306), .B0(n311), .CI(n233), .CO(n232), .S0(
        product[57]) );
  HS65_LH_FA1X4 U234 ( .A0(n312), .B0(n316), .CI(n234), .CO(n233), .S0(
        product[56]) );
  HS65_LH_FA1X4 U235 ( .A0(n317), .B0(n322), .CI(n235), .CO(n234), .S0(
        product[55]) );
  HS65_LH_FA1X4 U236 ( .A0(n323), .B0(n330), .CI(n236), .CO(n235), .S0(
        product[54]) );
  HS65_LH_FA1X4 U237 ( .A0(n331), .B0(n337), .CI(n237), .CO(n236), .S0(
        product[53]) );
  HS65_LH_FA1X4 U238 ( .A0(n338), .B0(n344), .CI(n238), .CO(n237), .S0(
        product[52]) );
  HS65_LH_FA1X4 U239 ( .A0(n345), .B0(n354), .CI(n239), .CO(n238), .S0(
        product[51]) );
  HS65_LH_FA1X4 U240 ( .A0(n355), .B0(n363), .CI(n240), .CO(n239), .S0(
        product[50]) );
  HS65_LH_FA1X4 U241 ( .A0(n364), .B0(n373), .CI(n241), .CO(n240), .S0(
        product[49]) );
  HS65_LH_FA1X4 U242 ( .A0(n374), .B0(n385), .CI(n242), .CO(n241), .S0(
        product[48]) );
  HS65_LH_FA1X4 U243 ( .A0(n386), .B0(n396), .CI(n243), .CO(n242), .S0(
        product[47]) );
  HS65_LH_FA1X4 U244 ( .A0(n397), .B0(n407), .CI(n244), .CO(n243), .S0(
        product[46]) );
  HS65_LH_FA1X4 U245 ( .A0(n408), .B0(n421), .CI(n245), .CO(n244), .S0(
        product[45]) );
  HS65_LH_FA1X4 U246 ( .A0(n422), .B0(n434), .CI(n246), .CO(n245), .S0(
        product[44]) );
  HS65_LH_FA1X4 U247 ( .A0(n435), .B0(n448), .CI(n247), .CO(n246), .S0(
        product[43]) );
  HS65_LH_FA1X4 U248 ( .A0(n449), .B0(n464), .CI(n248), .CO(n247), .S0(
        product[42]) );
  HS65_LH_FA1X4 U249 ( .A0(n465), .B0(n479), .CI(n249), .CO(n248), .S0(
        product[41]) );
  HS65_LH_FA1X4 U250 ( .A0(n480), .B0(n494), .CI(n250), .CO(n249), .S0(
        product[40]) );
  HS65_LH_FA1X4 U251 ( .A0(n495), .B0(n512), .CI(n251), .CO(n250), .S0(
        product[39]) );
  HS65_LH_FA1X4 U252 ( .A0(n513), .B0(n529), .CI(n252), .CO(n251), .S0(
        product[38]) );
  HS65_LH_FA1X4 U253 ( .A0(n530), .B0(n546), .CI(n253), .CO(n252), .S0(
        product[37]) );
  HS65_LH_FA1X4 U254 ( .A0(n547), .B0(n564), .CI(n254), .CO(n253), .S0(
        product[36]) );
  HS65_LH_FA1X4 U255 ( .A0(n565), .B0(n582), .CI(n255), .CO(n254), .S0(
        product[35]) );
  HS65_LH_FA1X4 U256 ( .A0(n583), .B0(n600), .CI(n256), .CO(n255), .S0(
        product[34]) );
  HS65_LH_FA1X4 U257 ( .A0(n601), .B0(n1386), .CI(n257), .CO(n256), .S0(
        product[33]) );
  HS65_LH_FA1X4 U258 ( .A0(n1387), .B0(n619), .CI(n258), .CO(n257), .S0(
        product[32]) );
  HS65_LH_FA1X4 U259 ( .A0(n1388), .B0(n637), .CI(n259), .CO(n258), .S0(
        product[31]) );
  HS65_LH_FA1X4 U260 ( .A0(n1389), .B0(n655), .CI(n260), .CO(n259), .S0(
        product[30]) );
  HS65_LH_FA1X4 U261 ( .A0(n1390), .B0(n673), .CI(n261), .CO(n260), .S0(
        product[29]) );
  HS65_LH_FA1X4 U262 ( .A0(n1391), .B0(n691), .CI(n262), .CO(n261), .S0(
        product[28]) );
  HS65_LH_FA1X4 U263 ( .A0(n1392), .B0(n709), .CI(n263), .CO(n262), .S0(
        product[27]) );
  HS65_LH_FA1X4 U264 ( .A0(n1393), .B0(n727), .CI(n264), .CO(n263), .S0(
        product[26]) );
  HS65_LH_FA1X4 U265 ( .A0(n1394), .B0(n743), .CI(n265), .CO(n264), .S0(
        product[25]) );
  HS65_LH_FA1X4 U266 ( .A0(n1395), .B0(n759), .CI(n266), .CO(n265), .S0(
        product[24]) );
  HS65_LH_FA1X4 U267 ( .A0(n1396), .B0(n775), .CI(n267), .CO(n266), .S0(
        product[23]) );
  HS65_LH_FA1X4 U268 ( .A0(n1397), .B0(n789), .CI(n268), .CO(n267), .S0(
        product[22]) );
  HS65_LH_FA1X4 U269 ( .A0(n1398), .B0(n803), .CI(n269), .CO(n268), .S0(
        product[21]) );
  HS65_LH_FA1X4 U270 ( .A0(n1399), .B0(n817), .CI(n270), .CO(n269), .S0(
        product[20]) );
  HS65_LH_FA1X4 U271 ( .A0(n1400), .B0(n829), .CI(n271), .CO(n270), .S0(
        product[19]) );
  HS65_LH_FA1X4 U272 ( .A0(n1401), .B0(n841), .CI(n272), .CO(n271), .S0(
        product[18]) );
  HS65_LH_FA1X4 U273 ( .A0(n1402), .B0(n853), .CI(n273), .CO(n272), .S0(
        product[17]) );
  HS65_LH_FA1X4 U274 ( .A0(n1403), .B0(n863), .CI(n274), .CO(n273), .S0(
        product[16]) );
  HS65_LH_FA1X4 U275 ( .A0(n1404), .B0(n873), .CI(n275), .CO(n274), .S0(
        product[15]) );
  HS65_LH_FA1X4 U276 ( .A0(n1405), .B0(n883), .CI(n276), .CO(n275), .S0(
        product[14]) );
  HS65_LH_FA1X4 U277 ( .A0(n1406), .B0(n891), .CI(n277), .CO(n276), .S0(
        product[13]) );
  HS65_LH_FA1X4 U278 ( .A0(n1407), .B0(n899), .CI(n278), .CO(n277), .S0(
        product[12]) );
  HS65_LH_FA1X4 U279 ( .A0(n1408), .B0(n907), .CI(n279), .CO(n278), .S0(
        product[11]) );
  HS65_LH_FA1X4 U280 ( .A0(n1409), .B0(n913), .CI(n280), .CO(n279), .S0(
        product[10]) );
  HS65_LH_FA1X4 U281 ( .A0(n1410), .B0(n919), .CI(n281), .CO(n280), .S0(
        product[9]) );
  HS65_LH_FA1X4 U282 ( .A0(n1411), .B0(n925), .CI(n282), .CO(n281), .S0(
        product[8]) );
  HS65_LH_FA1X4 U283 ( .A0(n1412), .B0(n929), .CI(n283), .CO(n282), .S0(
        product[7]) );
  HS65_LH_FA1X4 U284 ( .A0(n1413), .B0(n933), .CI(n284), .CO(n283), .S0(
        product[6]) );
  HS65_LH_FA1X4 U285 ( .A0(n1414), .B0(n937), .CI(n285), .CO(n284), .S0(
        product[5]) );
  HS65_LH_FA1X4 U286 ( .A0(n1415), .B0(n939), .CI(n286), .CO(n285), .S0(
        product[4]) );
  HS65_LH_FA1X4 U287 ( .A0(n1416), .B0(n941), .CI(n287), .CO(n286), .S0(
        product[3]) );
  HS65_LH_HA1X4 U288 ( .A0(n1417), .B0(n288), .CO(n287), .S0(product[2]) );
  HS65_LH_HA1X4 U289 ( .A0(n1418), .B0(n289), .CO(n288), .S0(product[1]) );
  HS65_LH_HA1X4 U290 ( .A0(n7), .B0(n1419), .CO(n289), .S0(product[0]) );
  HS65_LH_FA1X4 U293 ( .A0(n297), .B0(n2646), .CI(n1041), .CO(n293), .S0(n294)
         );
  HS65_LH_FA1X4 U294 ( .A0(n1042), .B0(n2647), .CI(n1071), .CO(n295), .S0(n296) );
  HS65_LH_FA1X4 U296 ( .A0(n2647), .B0(n1043), .CI(n1072), .CO(n299), .S0(n300) );
  HS65_LH_FA1X4 U298 ( .A0(n1073), .B0(n304), .CI(n307), .CO(n302), .S0(n303)
         );
  HS65_LH_FA1X4 U299 ( .A0(n309), .B0(n2644), .CI(n1044), .CO(n297), .S0(n304)
         );
  HS65_LH_FA1X4 U300 ( .A0(n1106), .B0(n1074), .CI(n308), .CO(n305), .S0(n306)
         );
  HS65_LH_FA1X4 U301 ( .A0(n1045), .B0(n2652), .CI(n313), .CO(n307), .S0(n308)
         );
  HS65_LH_FA1X4 U303 ( .A0(n314), .B0(n318), .CI(n1107), .CO(n311), .S0(n312)
         );
  HS65_LH_FA1X4 U304 ( .A0(n2652), .B0(n320), .CI(n1075), .CO(n313), .S0(n314)
         );
  HS65_LH_FA1X4 U306 ( .A0(n1108), .B0(n319), .CI(n324), .CO(n316), .S0(n317)
         );
  HS65_LH_FA1X4 U307 ( .A0(n326), .B0(n321), .CI(n1076), .CO(n318), .S0(n319)
         );
  HS65_LH_FA1X4 U308 ( .A0(n328), .B0(n2642), .CI(n1046), .CO(n320), .S0(n321)
         );
  HS65_LH_FA1X4 U309 ( .A0(n1141), .B0(n1109), .CI(n325), .CO(n322), .S0(n323)
         );
  HS65_LH_FA1X4 U310 ( .A0(n327), .B0(n334), .CI(n332), .CO(n324), .S0(n325)
         );
  HS65_LH_FA1X4 U311 ( .A0(n1047), .B0(n2648), .CI(n1077), .CO(n326), .S0(n327) );
  HS65_LH_FA1X4 U313 ( .A0(n333), .B0(n339), .CI(n1142), .CO(n330), .S0(n331)
         );
  HS65_LH_FA1X4 U314 ( .A0(n335), .B0(n341), .CI(n1110), .CO(n332), .S0(n333)
         );
  HS65_LH_FA1X4 U315 ( .A0(n2648), .B0(n1048), .CI(n1078), .CO(n334), .S0(n335) );
  HS65_LH_FA1X4 U317 ( .A0(n1143), .B0(n340), .CI(n346), .CO(n337), .S0(n338)
         );
  HS65_LH_FA1X4 U318 ( .A0(n348), .B0(n342), .CI(n1111), .CO(n339), .S0(n340)
         );
  HS65_LH_FA1X4 U319 ( .A0(n1079), .B0(n343), .CI(n350), .CO(n341), .S0(n342)
         );
  HS65_LH_FA1X4 U320 ( .A0(n352), .B0(n2640), .CI(n1049), .CO(n328), .S0(n343)
         );
  HS65_LH_FA1X4 U321 ( .A0(n1176), .B0(n1144), .CI(n347), .CO(n344), .S0(n345)
         );
  HS65_LH_FA1X4 U322 ( .A0(n349), .B0(n358), .CI(n356), .CO(n346), .S0(n347)
         );
  HS65_LH_FA1X4 U323 ( .A0(n351), .B0(n1080), .CI(n1112), .CO(n348), .S0(n349)
         );
  HS65_LH_FA1X4 U324 ( .A0(n1050), .B0(n2653), .CI(n360), .CO(n350), .S0(n351)
         );
  HS65_LH_FA1X4 U326 ( .A0(n357), .B0(n365), .CI(n1177), .CO(n354), .S0(n355)
         );
  HS65_LH_FA1X4 U327 ( .A0(n359), .B0(n367), .CI(n1145), .CO(n356), .S0(n357)
         );
  HS65_LH_FA1X4 U328 ( .A0(n361), .B0(n369), .CI(n1113), .CO(n358), .S0(n359)
         );
  HS65_LH_FA1X4 U329 ( .A0(n2653), .B0(n371), .CI(n1081), .CO(n360), .S0(n361)
         );
  HS65_LH_FA1X4 U331 ( .A0(n1178), .B0(n366), .CI(n375), .CO(n363), .S0(n364)
         );
  HS65_LH_FA1X4 U332 ( .A0(n377), .B0(n368), .CI(n1146), .CO(n365), .S0(n366)
         );
  HS65_LH_FA1X4 U333 ( .A0(n1114), .B0(n370), .CI(n379), .CO(n367), .S0(n368)
         );
  HS65_LH_FA1X4 U334 ( .A0(n381), .B0(n372), .CI(n1082), .CO(n369), .S0(n370)
         );
  HS65_LH_FA1X4 U335 ( .A0(n383), .B0(n2638), .CI(n1051), .CO(n371), .S0(n372)
         );
  HS65_LH_FA1X4 U336 ( .A0(n1211), .B0(n1179), .CI(n376), .CO(n373), .S0(n374)
         );
  HS65_LH_FA1X4 U337 ( .A0(n378), .B0(n389), .CI(n387), .CO(n375), .S0(n376)
         );
  HS65_LH_FA1X4 U338 ( .A0(n380), .B0(n1115), .CI(n1147), .CO(n377), .S0(n378)
         );
  HS65_LH_FA1X4 U339 ( .A0(n382), .B0(n393), .CI(n391), .CO(n379), .S0(n380)
         );
  HS65_LH_FA1X4 U340 ( .A0(n1052), .B0(n2649), .CI(n1083), .CO(n381), .S0(n382) );
  HS65_LH_FA1X4 U342 ( .A0(n388), .B0(n398), .CI(n1212), .CO(n385), .S0(n386)
         );
  HS65_LH_FA1X4 U343 ( .A0(n390), .B0(n400), .CI(n1180), .CO(n387), .S0(n388)
         );
  HS65_LH_FA1X4 U344 ( .A0(n392), .B0(n402), .CI(n1148), .CO(n389), .S0(n390)
         );
  HS65_LH_FA1X4 U345 ( .A0(n394), .B0(n404), .CI(n1116), .CO(n391), .S0(n392)
         );
  HS65_LH_FA1X4 U346 ( .A0(n2649), .B0(n1053), .CI(n1084), .CO(n393), .S0(n394) );
  HS65_LH_FA1X4 U348 ( .A0(n1213), .B0(n399), .CI(n409), .CO(n396), .S0(n397)
         );
  HS65_LH_FA1X4 U349 ( .A0(n411), .B0(n401), .CI(n1181), .CO(n398), .S0(n399)
         );
  HS65_LH_FA1X4 U350 ( .A0(n1149), .B0(n403), .CI(n413), .CO(n400), .S0(n401)
         );
  HS65_LH_FA1X4 U351 ( .A0(n415), .B0(n405), .CI(n1117), .CO(n402), .S0(n403)
         );
  HS65_LH_FA1X4 U352 ( .A0(n1085), .B0(n406), .CI(n417), .CO(n404), .S0(n405)
         );
  HS65_LH_FA1X4 U353 ( .A0(n419), .B0(n2636), .CI(n1054), .CO(n383), .S0(n406)
         );
  HS65_LH_FA1X4 U354 ( .A0(n1246), .B0(n1214), .CI(n410), .CO(n407), .S0(n408)
         );
  HS65_LH_FA1X4 U355 ( .A0(n412), .B0(n425), .CI(n423), .CO(n409), .S0(n410)
         );
  HS65_LH_FA1X4 U356 ( .A0(n414), .B0(n1150), .CI(n1182), .CO(n411), .S0(n412)
         );
  HS65_LH_FA1X4 U357 ( .A0(n416), .B0(n429), .CI(n427), .CO(n413), .S0(n414)
         );
  HS65_LH_FA1X4 U358 ( .A0(n418), .B0(n1086), .CI(n1118), .CO(n415), .S0(n416)
         );
  HS65_LH_FA1X4 U359 ( .A0(n1055), .B0(n2654), .CI(n431), .CO(n417), .S0(n418)
         );
  HS65_LH_FA1X4 U361 ( .A0(n424), .B0(n436), .CI(n1247), .CO(n421), .S0(n422)
         );
  HS65_LH_FA1X4 U362 ( .A0(n426), .B0(n438), .CI(n1215), .CO(n423), .S0(n424)
         );
  HS65_LH_FA1X4 U363 ( .A0(n428), .B0(n440), .CI(n1183), .CO(n425), .S0(n426)
         );
  HS65_LH_FA1X4 U364 ( .A0(n430), .B0(n442), .CI(n1151), .CO(n427), .S0(n428)
         );
  HS65_LH_FA1X4 U365 ( .A0(n432), .B0(n444), .CI(n1119), .CO(n429), .S0(n430)
         );
  HS65_LH_FA1X4 U366 ( .A0(n2654), .B0(n446), .CI(n1087), .CO(n431), .S0(n432)
         );
  HS65_LH_FA1X4 U368 ( .A0(n1248), .B0(n437), .CI(n450), .CO(n434), .S0(n435)
         );
  HS65_LH_FA1X4 U369 ( .A0(n452), .B0(n439), .CI(n1216), .CO(n436), .S0(n437)
         );
  HS65_LH_FA1X4 U370 ( .A0(n1184), .B0(n441), .CI(n454), .CO(n438), .S0(n439)
         );
  HS65_LH_FA1X4 U371 ( .A0(n456), .B0(n443), .CI(n1152), .CO(n440), .S0(n441)
         );
  HS65_LH_FA1X4 U372 ( .A0(n1120), .B0(n445), .CI(n458), .CO(n442), .S0(n443)
         );
  HS65_LH_FA1X4 U373 ( .A0(n460), .B0(n447), .CI(n1088), .CO(n444), .S0(n445)
         );
  HS65_LH_FA1X4 U374 ( .A0(n462), .B0(n2634), .CI(n1056), .CO(n446), .S0(n447)
         );
  HS65_LH_FA1X4 U375 ( .A0(n1281), .B0(n1249), .CI(n451), .CO(n448), .S0(n449)
         );
  HS65_LH_FA1X4 U376 ( .A0(n453), .B0(n468), .CI(n466), .CO(n450), .S0(n451)
         );
  HS65_LH_FA1X4 U377 ( .A0(n455), .B0(n1185), .CI(n1217), .CO(n452), .S0(n453)
         );
  HS65_LH_FA1X4 U378 ( .A0(n457), .B0(n472), .CI(n470), .CO(n454), .S0(n455)
         );
  HS65_LH_FA1X4 U379 ( .A0(n459), .B0(n1121), .CI(n1153), .CO(n456), .S0(n457)
         );
  HS65_LH_FA1X4 U380 ( .A0(n461), .B0(n476), .CI(n474), .CO(n458), .S0(n459)
         );
  HS65_LH_FA1X4 U381 ( .A0(n1057), .B0(n2650), .CI(n1089), .CO(n460), .S0(n461) );
  HS65_LH_FA1X4 U383 ( .A0(n467), .B0(n481), .CI(n1282), .CO(n464), .S0(n465)
         );
  HS65_LH_FA1X4 U384 ( .A0(n469), .B0(n483), .CI(n1250), .CO(n466), .S0(n467)
         );
  HS65_LH_FA1X4 U385 ( .A0(n471), .B0(n485), .CI(n1218), .CO(n468), .S0(n469)
         );
  HS65_LH_FA1X4 U386 ( .A0(n473), .B0(n487), .CI(n1186), .CO(n470), .S0(n471)
         );
  HS65_LH_FA1X4 U387 ( .A0(n475), .B0(n489), .CI(n1154), .CO(n472), .S0(n473)
         );
  HS65_LH_FA1X4 U388 ( .A0(n477), .B0(n491), .CI(n1122), .CO(n474), .S0(n475)
         );
  HS65_LH_FA1X4 U389 ( .A0(n2650), .B0(n1058), .CI(n1090), .CO(n476), .S0(n477) );
  HS65_LH_FA1X4 U391 ( .A0(n1283), .B0(n482), .CI(n496), .CO(n479), .S0(n480)
         );
  HS65_LH_FA1X4 U392 ( .A0(n498), .B0(n484), .CI(n1251), .CO(n481), .S0(n482)
         );
  HS65_LH_FA1X4 U393 ( .A0(n1219), .B0(n486), .CI(n500), .CO(n483), .S0(n484)
         );
  HS65_LH_FA1X4 U394 ( .A0(n502), .B0(n488), .CI(n1187), .CO(n485), .S0(n486)
         );
  HS65_LH_FA1X4 U395 ( .A0(n1155), .B0(n490), .CI(n504), .CO(n487), .S0(n488)
         );
  HS65_LH_FA1X4 U396 ( .A0(n506), .B0(n492), .CI(n1123), .CO(n489), .S0(n490)
         );
  HS65_LH_FA1X4 U397 ( .A0(n1091), .B0(n493), .CI(n508), .CO(n491), .S0(n492)
         );
  HS65_LH_FA1X4 U398 ( .A0(n510), .B0(n2632), .CI(n1059), .CO(n462), .S0(n493)
         );
  HS65_LH_FA1X4 U399 ( .A0(n1316), .B0(n1284), .CI(n497), .CO(n494), .S0(n495)
         );
  HS65_LH_FA1X4 U400 ( .A0(n499), .B0(n516), .CI(n514), .CO(n496), .S0(n497)
         );
  HS65_LH_FA1X4 U401 ( .A0(n501), .B0(n1220), .CI(n1252), .CO(n498), .S0(n499)
         );
  HS65_LH_FA1X4 U402 ( .A0(n503), .B0(n520), .CI(n518), .CO(n500), .S0(n501)
         );
  HS65_LH_FA1X4 U403 ( .A0(n505), .B0(n1156), .CI(n1188), .CO(n502), .S0(n503)
         );
  HS65_LH_FA1X4 U404 ( .A0(n507), .B0(n524), .CI(n522), .CO(n504), .S0(n505)
         );
  HS65_LH_FA1X4 U405 ( .A0(n509), .B0(n1092), .CI(n1124), .CO(n506), .S0(n507)
         );
  HS65_LH_FA1X4 U406 ( .A0(n1060), .B0(n2651), .CI(n526), .CO(n508), .S0(n509)
         );
  HS65_LH_FA1X4 U408 ( .A0(n515), .B0(n531), .CI(n1317), .CO(n512), .S0(n513)
         );
  HS65_LH_FA1X4 U409 ( .A0(n517), .B0(n533), .CI(n1285), .CO(n514), .S0(n515)
         );
  HS65_LH_FA1X4 U410 ( .A0(n519), .B0(n535), .CI(n1253), .CO(n516), .S0(n517)
         );
  HS65_LH_FA1X4 U411 ( .A0(n521), .B0(n537), .CI(n1221), .CO(n518), .S0(n519)
         );
  HS65_LH_FA1X4 U412 ( .A0(n523), .B0(n539), .CI(n1189), .CO(n520), .S0(n521)
         );
  HS65_LH_FA1X4 U413 ( .A0(n525), .B0(n541), .CI(n1157), .CO(n522), .S0(n523)
         );
  HS65_LH_FA1X4 U414 ( .A0(n527), .B0(n543), .CI(n1125), .CO(n524), .S0(n525)
         );
  HS65_LH_FA1X4 U415 ( .A0(n2651), .B0(n1061), .CI(n1093), .CO(n526), .S0(n527) );
  HS65_LH_FA1X4 U417 ( .A0(n1318), .B0(n532), .CI(n548), .CO(n529), .S0(n530)
         );
  HS65_LH_FA1X4 U418 ( .A0(n550), .B0(n534), .CI(n1286), .CO(n531), .S0(n532)
         );
  HS65_LH_FA1X4 U419 ( .A0(n1254), .B0(n536), .CI(n552), .CO(n533), .S0(n534)
         );
  HS65_LH_FA1X4 U420 ( .A0(n554), .B0(n538), .CI(n1222), .CO(n535), .S0(n536)
         );
  HS65_LH_FA1X4 U421 ( .A0(n1190), .B0(n540), .CI(n556), .CO(n537), .S0(n538)
         );
  HS65_LH_FA1X4 U422 ( .A0(n1158), .B0(n542), .CI(n558), .CO(n539), .S0(n540)
         );
  HS65_LH_FA1X4 U423 ( .A0(n1126), .B0(n544), .CI(n560), .CO(n541), .S0(n542)
         );
  HS65_LH_FA1X4 U424 ( .A0(n562), .B0(n545), .CI(n1094), .CO(n543), .S0(n544)
         );
  HS65_LH_FA1X4 U425 ( .A0(n2630), .B0(n2628), .CI(n1062), .CO(n510), .S0(n545) );
  HS65_LH_FA1X4 U426 ( .A0(n1351), .B0(n1319), .CI(n549), .CO(n546), .S0(n547)
         );
  HS65_LH_FA1X4 U427 ( .A0(n551), .B0(n1287), .CI(n566), .CO(n548), .S0(n549)
         );
  HS65_LH_FA1X4 U428 ( .A0(n553), .B0(n1255), .CI(n568), .CO(n550), .S0(n551)
         );
  HS65_LH_FA1X4 U429 ( .A0(n555), .B0(n572), .CI(n570), .CO(n552), .S0(n553)
         );
  HS65_LH_FA1X4 U430 ( .A0(n557), .B0(n1191), .CI(n1223), .CO(n554), .S0(n555)
         );
  HS65_LH_FA1X4 U431 ( .A0(n559), .B0(n576), .CI(n574), .CO(n556), .S0(n557)
         );
  HS65_LH_FA1X4 U432 ( .A0(n561), .B0(n1127), .CI(n1159), .CO(n558), .S0(n559)
         );
  HS65_LH_FA1X4 U433 ( .A0(n563), .B0(n1095), .CI(n578), .CO(n560), .S0(n561)
         );
  HS65_LH_FA1X4 U434 ( .A0(n1063), .B0(n7), .CI(n580), .CO(n562), .S0(n563) );
  HS65_LH_FA1X4 U435 ( .A0(n567), .B0(n1320), .CI(n1352), .CO(n564), .S0(n565)
         );
  HS65_LH_FA1X4 U436 ( .A0(n569), .B0(n1288), .CI(n584), .CO(n566), .S0(n567)
         );
  HS65_LH_FA1X4 U437 ( .A0(n571), .B0(n1256), .CI(n586), .CO(n568), .S0(n569)
         );
  HS65_LH_FA1X4 U438 ( .A0(n573), .B0(n590), .CI(n588), .CO(n570), .S0(n571)
         );
  HS65_LH_FA1X4 U439 ( .A0(n575), .B0(n1192), .CI(n1224), .CO(n572), .S0(n573)
         );
  HS65_LH_FA1X4 U440 ( .A0(n577), .B0(n594), .CI(n592), .CO(n574), .S0(n575)
         );
  HS65_LH_FA1X4 U441 ( .A0(n579), .B0(n1128), .CI(n1160), .CO(n576), .S0(n577)
         );
  HS65_LH_FA1X4 U442 ( .A0(n581), .B0(n1096), .CI(n596), .CO(n578), .S0(n579)
         );
  HS65_LH_FA1X4 U443 ( .A0(n1064), .B0(n7), .CI(n598), .CO(n580), .S0(n581) );
  HS65_LH_FA1X4 U444 ( .A0(n585), .B0(n602), .CI(n1353), .CO(n582), .S0(n583)
         );
  HS65_LH_FA1X4 U445 ( .A0(n587), .B0(n604), .CI(n1321), .CO(n584), .S0(n585)
         );
  HS65_LH_FA1X4 U446 ( .A0(n589), .B0(n606), .CI(n1289), .CO(n586), .S0(n587)
         );
  HS65_LH_FA1X4 U447 ( .A0(n591), .B0(n608), .CI(n1257), .CO(n588), .S0(n589)
         );
  HS65_LH_FA1X4 U448 ( .A0(n593), .B0(n610), .CI(n1225), .CO(n590), .S0(n591)
         );
  HS65_LH_FA1X4 U449 ( .A0(n595), .B0(n612), .CI(n1193), .CO(n592), .S0(n593)
         );
  HS65_LH_FA1X4 U450 ( .A0(n597), .B0(n614), .CI(n1161), .CO(n594), .S0(n595)
         );
  HS65_LH_FA1X4 U451 ( .A0(n599), .B0(n616), .CI(n1129), .CO(n596), .S0(n597)
         );
  HS65_LH_FA1X4 U452 ( .A0(n1065), .B0(n7), .CI(n1097), .CO(n598), .S0(n599)
         );
  HS65_LH_FA1X4 U453 ( .A0(n1354), .B0(n603), .CI(n618), .CO(n600), .S0(n601)
         );
  HS65_LH_FA1X4 U454 ( .A0(n1322), .B0(n605), .CI(n620), .CO(n602), .S0(n603)
         );
  HS65_LH_FA1X4 U455 ( .A0(n1290), .B0(n607), .CI(n622), .CO(n604), .S0(n605)
         );
  HS65_LH_FA1X4 U456 ( .A0(n1258), .B0(n609), .CI(n624), .CO(n606), .S0(n607)
         );
  HS65_LH_FA1X4 U457 ( .A0(n1226), .B0(n611), .CI(n626), .CO(n608), .S0(n609)
         );
  HS65_LH_FA1X4 U458 ( .A0(n1194), .B0(n613), .CI(n628), .CO(n610), .S0(n611)
         );
  HS65_LH_FA1X4 U459 ( .A0(n1162), .B0(n615), .CI(n630), .CO(n612), .S0(n613)
         );
  HS65_LH_FA1X4 U460 ( .A0(n1130), .B0(n617), .CI(n632), .CO(n614), .S0(n615)
         );
  HS65_LH_FA1X4 U461 ( .A0(n1098), .B0(n1066), .CI(n634), .CO(n616), .S0(n617)
         );
  HS65_LH_FA1X4 U462 ( .A0(n1355), .B0(n621), .CI(n636), .CO(n618), .S0(n619)
         );
  HS65_LH_FA1X4 U463 ( .A0(n1323), .B0(n623), .CI(n638), .CO(n620), .S0(n621)
         );
  HS65_LH_FA1X4 U464 ( .A0(n1291), .B0(n625), .CI(n640), .CO(n622), .S0(n623)
         );
  HS65_LH_FA1X4 U465 ( .A0(n1259), .B0(n627), .CI(n642), .CO(n624), .S0(n625)
         );
  HS65_LH_FA1X4 U466 ( .A0(n1227), .B0(n629), .CI(n644), .CO(n626), .S0(n627)
         );
  HS65_LH_FA1X4 U467 ( .A0(n1195), .B0(n631), .CI(n646), .CO(n628), .S0(n629)
         );
  HS65_LH_FA1X4 U468 ( .A0(n1163), .B0(n633), .CI(n648), .CO(n630), .S0(n631)
         );
  HS65_LH_FA1X4 U469 ( .A0(n1131), .B0(n635), .CI(n650), .CO(n632), .S0(n633)
         );
  HS65_LH_FA1X4 U470 ( .A0(n1099), .B0(n1067), .CI(n652), .CO(n634), .S0(n635)
         );
  HS65_LH_FA1X4 U471 ( .A0(n1356), .B0(n639), .CI(n654), .CO(n636), .S0(n637)
         );
  HS65_LH_FA1X4 U472 ( .A0(n1324), .B0(n641), .CI(n656), .CO(n638), .S0(n639)
         );
  HS65_LH_FA1X4 U473 ( .A0(n1292), .B0(n643), .CI(n658), .CO(n640), .S0(n641)
         );
  HS65_LH_FA1X4 U474 ( .A0(n1260), .B0(n645), .CI(n660), .CO(n642), .S0(n643)
         );
  HS65_LH_FA1X4 U475 ( .A0(n1228), .B0(n647), .CI(n662), .CO(n644), .S0(n645)
         );
  HS65_LH_FA1X4 U476 ( .A0(n1196), .B0(n649), .CI(n664), .CO(n646), .S0(n647)
         );
  HS65_LH_FA1X4 U477 ( .A0(n1164), .B0(n651), .CI(n666), .CO(n648), .S0(n649)
         );
  HS65_LH_FA1X4 U478 ( .A0(n1132), .B0(n653), .CI(n668), .CO(n650), .S0(n651)
         );
  HS65_LH_FA1X4 U479 ( .A0(n1100), .B0(n1068), .CI(n670), .CO(n652), .S0(n653)
         );
  HS65_LH_FA1X4 U480 ( .A0(n1357), .B0(n657), .CI(n672), .CO(n654), .S0(n655)
         );
  HS65_LH_FA1X4 U481 ( .A0(n1325), .B0(n659), .CI(n674), .CO(n656), .S0(n657)
         );
  HS65_LH_FA1X4 U482 ( .A0(n1293), .B0(n661), .CI(n676), .CO(n658), .S0(n659)
         );
  HS65_LH_FA1X4 U483 ( .A0(n1261), .B0(n663), .CI(n678), .CO(n660), .S0(n661)
         );
  HS65_LH_FA1X4 U484 ( .A0(n1229), .B0(n665), .CI(n680), .CO(n662), .S0(n663)
         );
  HS65_LH_FA1X4 U485 ( .A0(n1197), .B0(n667), .CI(n682), .CO(n664), .S0(n665)
         );
  HS65_LH_FA1X4 U486 ( .A0(n1165), .B0(n669), .CI(n684), .CO(n666), .S0(n667)
         );
  HS65_LH_FA1X4 U487 ( .A0(n1133), .B0(n671), .CI(n686), .CO(n668), .S0(n669)
         );
  HS65_LH_FA1X4 U488 ( .A0(n1101), .B0(n1069), .CI(n688), .CO(n670), .S0(n671)
         );
  HS65_LH_FA1X4 U489 ( .A0(n1358), .B0(n675), .CI(n690), .CO(n672), .S0(n673)
         );
  HS65_LH_FA1X4 U490 ( .A0(n1326), .B0(n677), .CI(n692), .CO(n674), .S0(n675)
         );
  HS65_LH_FA1X4 U491 ( .A0(n1294), .B0(n679), .CI(n694), .CO(n676), .S0(n677)
         );
  HS65_LH_FA1X4 U492 ( .A0(n1262), .B0(n681), .CI(n696), .CO(n678), .S0(n679)
         );
  HS65_LH_FA1X4 U493 ( .A0(n1230), .B0(n683), .CI(n698), .CO(n680), .S0(n681)
         );
  HS65_LH_FA1X4 U494 ( .A0(n1198), .B0(n685), .CI(n700), .CO(n682), .S0(n683)
         );
  HS65_LH_FA1X4 U495 ( .A0(n1166), .B0(n687), .CI(n702), .CO(n684), .S0(n685)
         );
  HS65_LH_FA1X4 U496 ( .A0(n1134), .B0(n689), .CI(n704), .CO(n686), .S0(n687)
         );
  HS65_LH_HA1X4 U497 ( .A0(n1102), .B0(n706), .CO(n688), .S0(n689) );
  HS65_LH_FA1X4 U498 ( .A0(n1359), .B0(n693), .CI(n708), .CO(n690), .S0(n691)
         );
  HS65_LH_FA1X4 U499 ( .A0(n1327), .B0(n695), .CI(n710), .CO(n692), .S0(n693)
         );
  HS65_LH_FA1X4 U500 ( .A0(n1295), .B0(n697), .CI(n712), .CO(n694), .S0(n695)
         );
  HS65_LH_FA1X4 U501 ( .A0(n1263), .B0(n699), .CI(n714), .CO(n696), .S0(n697)
         );
  HS65_LH_FA1X4 U502 ( .A0(n1231), .B0(n701), .CI(n716), .CO(n698), .S0(n699)
         );
  HS65_LH_FA1X4 U503 ( .A0(n1199), .B0(n703), .CI(n718), .CO(n700), .S0(n701)
         );
  HS65_LH_FA1X4 U504 ( .A0(n1167), .B0(n705), .CI(n720), .CO(n702), .S0(n703)
         );
  HS65_LH_FA1X4 U505 ( .A0(n1135), .B0(n707), .CI(n722), .CO(n704), .S0(n705)
         );
  HS65_LH_HA1X4 U506 ( .A0(n1103), .B0(n724), .CO(n706), .S0(n707) );
  HS65_LH_FA1X4 U507 ( .A0(n1360), .B0(n711), .CI(n726), .CO(n708), .S0(n709)
         );
  HS65_LH_FA1X4 U508 ( .A0(n1328), .B0(n713), .CI(n728), .CO(n710), .S0(n711)
         );
  HS65_LH_FA1X4 U509 ( .A0(n1296), .B0(n715), .CI(n730), .CO(n712), .S0(n713)
         );
  HS65_LH_FA1X4 U510 ( .A0(n1264), .B0(n717), .CI(n732), .CO(n714), .S0(n715)
         );
  HS65_LH_FA1X4 U511 ( .A0(n1232), .B0(n719), .CI(n734), .CO(n716), .S0(n717)
         );
  HS65_LH_FA1X4 U512 ( .A0(n1200), .B0(n721), .CI(n736), .CO(n718), .S0(n719)
         );
  HS65_LH_FA1X4 U513 ( .A0(n1168), .B0(n723), .CI(n738), .CO(n720), .S0(n721)
         );
  HS65_LH_FA1X4 U514 ( .A0(n1136), .B0(n725), .CI(n740), .CO(n722), .S0(n723)
         );
  HS65_LH_HA1X4 U515 ( .A0(n2645), .B0(n1104), .CO(n724), .S0(n725) );
  HS65_LH_FA1X4 U516 ( .A0(n1361), .B0(n729), .CI(n742), .CO(n726), .S0(n727)
         );
  HS65_LH_FA1X4 U517 ( .A0(n1329), .B0(n731), .CI(n744), .CO(n728), .S0(n729)
         );
  HS65_LH_FA1X4 U518 ( .A0(n1297), .B0(n733), .CI(n746), .CO(n730), .S0(n731)
         );
  HS65_LH_FA1X4 U519 ( .A0(n1265), .B0(n735), .CI(n748), .CO(n732), .S0(n733)
         );
  HS65_LH_FA1X4 U520 ( .A0(n1233), .B0(n737), .CI(n750), .CO(n734), .S0(n735)
         );
  HS65_LH_FA1X4 U521 ( .A0(n1201), .B0(n739), .CI(n752), .CO(n736), .S0(n737)
         );
  HS65_LH_FA1X4 U522 ( .A0(n1169), .B0(n741), .CI(n754), .CO(n738), .S0(n739)
         );
  HS65_LH_HA1X4 U523 ( .A0(n1137), .B0(n756), .CO(n740), .S0(n741) );
  HS65_LH_FA1X4 U524 ( .A0(n1362), .B0(n745), .CI(n758), .CO(n742), .S0(n743)
         );
  HS65_LH_FA1X4 U525 ( .A0(n1330), .B0(n747), .CI(n760), .CO(n744), .S0(n745)
         );
  HS65_LH_FA1X4 U526 ( .A0(n1298), .B0(n749), .CI(n762), .CO(n746), .S0(n747)
         );
  HS65_LH_FA1X4 U527 ( .A0(n1266), .B0(n751), .CI(n764), .CO(n748), .S0(n749)
         );
  HS65_LH_FA1X4 U528 ( .A0(n1234), .B0(n753), .CI(n766), .CO(n750), .S0(n751)
         );
  HS65_LH_FA1X4 U529 ( .A0(n1202), .B0(n755), .CI(n768), .CO(n752), .S0(n753)
         );
  HS65_LH_FA1X4 U530 ( .A0(n1170), .B0(n757), .CI(n770), .CO(n754), .S0(n755)
         );
  HS65_LH_HA1X4 U531 ( .A0(n1138), .B0(n772), .CO(n756), .S0(n757) );
  HS65_LH_FA1X4 U532 ( .A0(n1363), .B0(n761), .CI(n774), .CO(n758), .S0(n759)
         );
  HS65_LH_FA1X4 U533 ( .A0(n1331), .B0(n763), .CI(n776), .CO(n760), .S0(n761)
         );
  HS65_LH_FA1X4 U534 ( .A0(n1299), .B0(n765), .CI(n778), .CO(n762), .S0(n763)
         );
  HS65_LH_FA1X4 U535 ( .A0(n1267), .B0(n767), .CI(n780), .CO(n764), .S0(n765)
         );
  HS65_LH_FA1X4 U536 ( .A0(n1235), .B0(n769), .CI(n782), .CO(n766), .S0(n767)
         );
  HS65_LH_FA1X4 U537 ( .A0(n1203), .B0(n771), .CI(n784), .CO(n768), .S0(n769)
         );
  HS65_LH_FA1X4 U538 ( .A0(n1171), .B0(n773), .CI(n786), .CO(n770), .S0(n771)
         );
  HS65_LH_HA1X4 U539 ( .A0(n103), .B0(n1139), .CO(n772), .S0(n773) );
  HS65_LH_FA1X4 U540 ( .A0(n1364), .B0(n777), .CI(n788), .CO(n774), .S0(n775)
         );
  HS65_LH_FA1X4 U541 ( .A0(n1332), .B0(n779), .CI(n790), .CO(n776), .S0(n777)
         );
  HS65_LH_FA1X4 U542 ( .A0(n1300), .B0(n781), .CI(n792), .CO(n778), .S0(n779)
         );
  HS65_LH_FA1X4 U543 ( .A0(n1268), .B0(n783), .CI(n794), .CO(n780), .S0(n781)
         );
  HS65_LH_FA1X4 U544 ( .A0(n1236), .B0(n785), .CI(n796), .CO(n782), .S0(n783)
         );
  HS65_LH_FA1X4 U545 ( .A0(n1204), .B0(n787), .CI(n798), .CO(n784), .S0(n785)
         );
  HS65_LH_HA1X4 U546 ( .A0(n1172), .B0(n800), .CO(n786), .S0(n787) );
  HS65_LH_FA1X4 U547 ( .A0(n1365), .B0(n791), .CI(n802), .CO(n788), .S0(n789)
         );
  HS65_LH_FA1X4 U548 ( .A0(n1333), .B0(n793), .CI(n804), .CO(n790), .S0(n791)
         );
  HS65_LH_FA1X4 U549 ( .A0(n1301), .B0(n795), .CI(n806), .CO(n792), .S0(n793)
         );
  HS65_LH_FA1X4 U550 ( .A0(n1269), .B0(n797), .CI(n808), .CO(n794), .S0(n795)
         );
  HS65_LH_FA1X4 U551 ( .A0(n1237), .B0(n799), .CI(n810), .CO(n796), .S0(n797)
         );
  HS65_LH_FA1X4 U552 ( .A0(n1205), .B0(n801), .CI(n812), .CO(n798), .S0(n799)
         );
  HS65_LH_HA1X4 U553 ( .A0(n1173), .B0(n814), .CO(n800), .S0(n801) );
  HS65_LH_FA1X4 U554 ( .A0(n1366), .B0(n805), .CI(n816), .CO(n802), .S0(n803)
         );
  HS65_LH_FA1X4 U555 ( .A0(n1334), .B0(n807), .CI(n818), .CO(n804), .S0(n805)
         );
  HS65_LH_FA1X4 U556 ( .A0(n1302), .B0(n809), .CI(n820), .CO(n806), .S0(n807)
         );
  HS65_LH_FA1X4 U557 ( .A0(n1270), .B0(n811), .CI(n822), .CO(n808), .S0(n809)
         );
  HS65_LH_FA1X4 U558 ( .A0(n1238), .B0(n813), .CI(n824), .CO(n810), .S0(n811)
         );
  HS65_LH_FA1X4 U559 ( .A0(n1206), .B0(n815), .CI(n826), .CO(n812), .S0(n813)
         );
  HS65_LH_HA1X4 U560 ( .A0(n91), .B0(n1174), .CO(n814), .S0(n815) );
  HS65_LH_FA1X4 U561 ( .A0(n1367), .B0(n819), .CI(n828), .CO(n816), .S0(n817)
         );
  HS65_LH_FA1X4 U562 ( .A0(n1335), .B0(n821), .CI(n830), .CO(n818), .S0(n819)
         );
  HS65_LH_FA1X4 U563 ( .A0(n1303), .B0(n823), .CI(n832), .CO(n820), .S0(n821)
         );
  HS65_LH_FA1X4 U564 ( .A0(n1271), .B0(n825), .CI(n834), .CO(n822), .S0(n823)
         );
  HS65_LH_FA1X4 U565 ( .A0(n1239), .B0(n827), .CI(n836), .CO(n824), .S0(n825)
         );
  HS65_LH_HA1X4 U566 ( .A0(n1207), .B0(n838), .CO(n826), .S0(n827) );
  HS65_LH_FA1X4 U567 ( .A0(n1368), .B0(n831), .CI(n840), .CO(n828), .S0(n829)
         );
  HS65_LH_FA1X4 U568 ( .A0(n1336), .B0(n833), .CI(n842), .CO(n830), .S0(n831)
         );
  HS65_LH_FA1X4 U569 ( .A0(n1304), .B0(n835), .CI(n844), .CO(n832), .S0(n833)
         );
  HS65_LH_FA1X4 U570 ( .A0(n1272), .B0(n837), .CI(n846), .CO(n834), .S0(n835)
         );
  HS65_LH_FA1X4 U571 ( .A0(n1240), .B0(n839), .CI(n848), .CO(n836), .S0(n837)
         );
  HS65_LH_HA1X4 U572 ( .A0(n1208), .B0(n850), .CO(n838), .S0(n839) );
  HS65_LH_FA1X4 U573 ( .A0(n1369), .B0(n843), .CI(n852), .CO(n840), .S0(n841)
         );
  HS65_LH_FA1X4 U574 ( .A0(n1337), .B0(n845), .CI(n854), .CO(n842), .S0(n843)
         );
  HS65_LH_FA1X4 U575 ( .A0(n1305), .B0(n847), .CI(n856), .CO(n844), .S0(n845)
         );
  HS65_LH_FA1X4 U576 ( .A0(n1273), .B0(n849), .CI(n858), .CO(n846), .S0(n847)
         );
  HS65_LH_FA1X4 U577 ( .A0(n1241), .B0(n851), .CI(n860), .CO(n848), .S0(n849)
         );
  HS65_LH_HA1X4 U578 ( .A0(n79), .B0(n1209), .CO(n850), .S0(n851) );
  HS65_LH_FA1X4 U579 ( .A0(n1370), .B0(n855), .CI(n862), .CO(n852), .S0(n853)
         );
  HS65_LH_FA1X4 U580 ( .A0(n1338), .B0(n857), .CI(n864), .CO(n854), .S0(n855)
         );
  HS65_LH_FA1X4 U581 ( .A0(n1306), .B0(n859), .CI(n866), .CO(n856), .S0(n857)
         );
  HS65_LH_FA1X4 U582 ( .A0(n1274), .B0(n861), .CI(n868), .CO(n858), .S0(n859)
         );
  HS65_LH_HA1X4 U583 ( .A0(n1242), .B0(n870), .CO(n860), .S0(n861) );
  HS65_LH_FA1X4 U584 ( .A0(n1371), .B0(n865), .CI(n872), .CO(n862), .S0(n863)
         );
  HS65_LH_FA1X4 U585 ( .A0(n1339), .B0(n867), .CI(n874), .CO(n864), .S0(n865)
         );
  HS65_LH_FA1X4 U586 ( .A0(n1307), .B0(n869), .CI(n876), .CO(n866), .S0(n867)
         );
  HS65_LH_FA1X4 U587 ( .A0(n1275), .B0(n871), .CI(n878), .CO(n868), .S0(n869)
         );
  HS65_LH_HA1X4 U588 ( .A0(n1243), .B0(n880), .CO(n870), .S0(n871) );
  HS65_LH_FA1X4 U589 ( .A0(n1372), .B0(n875), .CI(n882), .CO(n872), .S0(n873)
         );
  HS65_LH_FA1X4 U590 ( .A0(n1340), .B0(n877), .CI(n884), .CO(n874), .S0(n875)
         );
  HS65_LH_FA1X4 U591 ( .A0(n1308), .B0(n879), .CI(n886), .CO(n876), .S0(n877)
         );
  HS65_LH_FA1X4 U592 ( .A0(n1276), .B0(n881), .CI(n888), .CO(n878), .S0(n879)
         );
  HS65_LH_HA1X4 U593 ( .A0(n67), .B0(n1244), .CO(n880), .S0(n881) );
  HS65_LH_FA1X4 U594 ( .A0(n1373), .B0(n885), .CI(n890), .CO(n882), .S0(n883)
         );
  HS65_LH_FA1X4 U595 ( .A0(n1341), .B0(n887), .CI(n892), .CO(n884), .S0(n885)
         );
  HS65_LH_FA1X4 U596 ( .A0(n1309), .B0(n889), .CI(n894), .CO(n886), .S0(n887)
         );
  HS65_LH_HA1X4 U597 ( .A0(n1277), .B0(n896), .CO(n888), .S0(n889) );
  HS65_LH_FA1X4 U598 ( .A0(n1374), .B0(n893), .CI(n898), .CO(n890), .S0(n891)
         );
  HS65_LH_FA1X4 U599 ( .A0(n1342), .B0(n895), .CI(n900), .CO(n892), .S0(n893)
         );
  HS65_LH_FA1X4 U600 ( .A0(n1310), .B0(n897), .CI(n902), .CO(n894), .S0(n895)
         );
  HS65_LH_HA1X4 U601 ( .A0(n1278), .B0(n904), .CO(n896), .S0(n897) );
  HS65_LH_FA1X4 U602 ( .A0(n1375), .B0(n901), .CI(n906), .CO(n898), .S0(n899)
         );
  HS65_LH_FA1X4 U603 ( .A0(n1343), .B0(n903), .CI(n908), .CO(n900), .S0(n901)
         );
  HS65_LH_FA1X4 U604 ( .A0(n1311), .B0(n905), .CI(n910), .CO(n902), .S0(n903)
         );
  HS65_LH_HA1X4 U605 ( .A0(n55), .B0(n1279), .CO(n904), .S0(n905) );
  HS65_LH_FA1X4 U606 ( .A0(n1376), .B0(n909), .CI(n912), .CO(n906), .S0(n907)
         );
  HS65_LH_FA1X4 U607 ( .A0(n1344), .B0(n911), .CI(n914), .CO(n908), .S0(n909)
         );
  HS65_LH_HA1X4 U608 ( .A0(n1312), .B0(n916), .CO(n910), .S0(n911) );
  HS65_LH_FA1X4 U609 ( .A0(n1377), .B0(n915), .CI(n918), .CO(n912), .S0(n913)
         );
  HS65_LH_FA1X4 U610 ( .A0(n1345), .B0(n917), .CI(n920), .CO(n914), .S0(n915)
         );
  HS65_LH_HA1X4 U611 ( .A0(n1313), .B0(n922), .CO(n916), .S0(n917) );
  HS65_LH_FA1X4 U612 ( .A0(n1378), .B0(n921), .CI(n924), .CO(n918), .S0(n919)
         );
  HS65_LH_FA1X4 U613 ( .A0(n1346), .B0(n923), .CI(n926), .CO(n920), .S0(n921)
         );
  HS65_LH_HA1X4 U614 ( .A0(n43), .B0(n1314), .CO(n922), .S0(n923) );
  HS65_LH_FA1X4 U615 ( .A0(n1379), .B0(n927), .CI(n928), .CO(n924), .S0(n925)
         );
  HS65_LH_HA1X4 U616 ( .A0(n1347), .B0(n930), .CO(n926), .S0(n927) );
  HS65_LH_FA1X4 U617 ( .A0(n1380), .B0(n931), .CI(n932), .CO(n928), .S0(n929)
         );
  HS65_LH_HA1X4 U618 ( .A0(n1348), .B0(n934), .CO(n930), .S0(n931) );
  HS65_LH_FA1X4 U619 ( .A0(n1381), .B0(n935), .CI(n936), .CO(n932), .S0(n933)
         );
  HS65_LH_HA1X4 U620 ( .A0(n31), .B0(n1349), .CO(n934), .S0(n935) );
  HS65_LH_HA1X4 U621 ( .A0(n1382), .B0(n938), .CO(n936), .S0(n937) );
  HS65_LH_HA1X4 U622 ( .A0(n1383), .B0(n940), .CO(n938), .S0(n939) );
  HS65_LH_HA1X4 U623 ( .A0(n19), .B0(n1384), .CO(n940), .S0(n941) );
  HS65_LH_HA1X4 U1907 ( .A0(n2626), .B0(n975), .CO(n1006), .S0(n1007) );
  HS65_LH_FA1X4 U1908 ( .A0(n2624), .B0(n2626), .CI(n976), .CO(n975), .S0(
        n1008) );
  HS65_LH_FA1X4 U1909 ( .A0(n2622), .B0(n2624), .CI(n977), .CO(n976), .S0(
        n1009) );
  HS65_LH_FA1X4 U1910 ( .A0(n2620), .B0(n2622), .CI(n978), .CO(n977), .S0(
        n1010) );
  HS65_LH_FA1X4 U1911 ( .A0(n2618), .B0(n2620), .CI(n979), .CO(n978), .S0(
        n1011) );
  HS65_LH_FA1X4 U1912 ( .A0(n2616), .B0(n2618), .CI(n980), .CO(n979), .S0(
        n1012) );
  HS65_LH_FA1X4 U1913 ( .A0(n2614), .B0(n2616), .CI(n981), .CO(n980), .S0(
        n1013) );
  HS65_LH_FA1X4 U1914 ( .A0(n2612), .B0(n2614), .CI(n982), .CO(n981), .S0(
        n1014) );
  HS65_LH_FA1X4 U1915 ( .A0(n2610), .B0(n2612), .CI(n983), .CO(n982), .S0(
        n1015) );
  HS65_LH_FA1X4 U1916 ( .A0(n2608), .B0(n2610), .CI(n984), .CO(n983), .S0(
        n1016) );
  HS65_LH_FA1X4 U1917 ( .A0(n2606), .B0(n2608), .CI(n985), .CO(n984), .S0(
        n1017) );
  HS65_LH_FA1X4 U1918 ( .A0(n2604), .B0(n2606), .CI(n986), .CO(n985), .S0(
        n1018) );
  HS65_LH_FA1X4 U1919 ( .A0(n2602), .B0(n2604), .CI(n987), .CO(n986), .S0(
        n1019) );
  HS65_LH_FA1X4 U1920 ( .A0(n2600), .B0(n2602), .CI(n988), .CO(n987), .S0(
        n1020) );
  HS65_LH_FA1X4 U1921 ( .A0(n2598), .B0(n2600), .CI(n989), .CO(n988), .S0(
        n1021) );
  HS65_LH_FA1X4 U1922 ( .A0(n2596), .B0(n2598), .CI(n990), .CO(n989), .S0(
        n1022) );
  HS65_LH_FA1X4 U1923 ( .A0(n2594), .B0(n2596), .CI(n991), .CO(n990), .S0(
        n1023) );
  HS65_LH_FA1X4 U1924 ( .A0(n2592), .B0(n2594), .CI(n992), .CO(n991), .S0(
        n1024) );
  HS65_LH_FA1X4 U1925 ( .A0(n2590), .B0(n2592), .CI(n993), .CO(n992), .S0(
        n1025) );
  HS65_LH_FA1X4 U1926 ( .A0(n2588), .B0(n2590), .CI(n994), .CO(n993), .S0(
        n1026) );
  HS65_LH_FA1X4 U1927 ( .A0(n2586), .B0(n2588), .CI(n995), .CO(n994), .S0(
        n1027) );
  HS65_LH_FA1X4 U1928 ( .A0(n2584), .B0(n2586), .CI(n996), .CO(n995), .S0(
        n1028) );
  HS65_LH_FA1X4 U1929 ( .A0(n2582), .B0(n2584), .CI(n997), .CO(n996), .S0(
        n1029) );
  HS65_LH_FA1X4 U1930 ( .A0(n2580), .B0(n2582), .CI(n998), .CO(n997), .S0(
        n1030) );
  HS65_LH_FA1X4 U1931 ( .A0(n2578), .B0(n2580), .CI(n999), .CO(n998), .S0(
        n1031) );
  HS65_LH_FA1X4 U1932 ( .A0(n2576), .B0(n2578), .CI(n1000), .CO(n999), .S0(
        n1032) );
  HS65_LH_FA1X4 U1933 ( .A0(n2574), .B0(n2576), .CI(n1001), .CO(n1000), .S0(
        n1033) );
  HS65_LH_FA1X4 U1934 ( .A0(n2572), .B0(n2574), .CI(n1002), .CO(n1001), .S0(
        n1034) );
  HS65_LH_FA1X4 U1935 ( .A0(n2570), .B0(n2572), .CI(n1003), .CO(n1002), .S0(
        n1035) );
  HS65_LH_FA1X4 U1936 ( .A0(n2568), .B0(n2570), .CI(n1004), .CO(n1003), .S0(
        n1036) );
  HS65_LH_FA1X4 U1937 ( .A0(n2566), .B0(n2568), .CI(n1005), .CO(n1004), .S0(
        n1037) );
  HS65_LH_IVX9 U1941 ( .A(n7), .Z(n2628) );
  HS65_LH_IVX9 U1942 ( .A(n1007), .Z(n2657) );
  HS65_LH_IVX9 U1943 ( .A(n419), .Z(n2654) );
  HS65_LH_IVX9 U1944 ( .A(n352), .Z(n2653) );
  HS65_LH_IVX9 U1945 ( .A(n309), .Z(n2652) );
  HS65_LH_IVX9 U1946 ( .A(n510), .Z(n2651) );
  HS65_LH_IVX9 U1947 ( .A(n462), .Z(n2650) );
  HS65_LH_IVX9 U1948 ( .A(n383), .Z(n2649) );
  HS65_LH_IVX9 U1949 ( .A(n328), .Z(n2648) );
  HS65_LH_IVX9 U1950 ( .A(n297), .Z(n2647) );
  HS65_LH_HA1X4 U1951 ( .A0(n2566), .B0(n2563), .CO(n1005), .S0(n1038) );
  HS65_LH_BFX9 U1952 ( .A(b[27]), .Z(n2618) );
  HS65_LH_BFX9 U1953 ( .A(b[3]), .Z(n2570) );
  HS65_LH_BFX9 U1954 ( .A(b[2]), .Z(n2568) );
  HS65_LH_BFX9 U1955 ( .A(b[20]), .Z(n2604) );
  HS65_LH_BFX9 U1956 ( .A(b[11]), .Z(n2586) );
  HS65_LH_BFX9 U1957 ( .A(b[4]), .Z(n2572) );
  HS65_LH_BFX9 U1958 ( .A(b[28]), .Z(n2620) );
  HS65_LH_BFX9 U1959 ( .A(n2655), .Z(n2418) );
  HS65_LH_BFX9 U1960 ( .A(n2655), .Z(n2417) );
  HS65_LH_BFX9 U1961 ( .A(n2656), .Z(n2421) );
  HS65_LH_BFX9 U1962 ( .A(n2656), .Z(n2420) );
  HS65_LH_BFX9 U1963 ( .A(b[31]), .Z(n2626) );
  HS65_LH_BFX9 U1964 ( .A(n2655), .Z(n2419) );
  HS65_LH_BFX9 U1965 ( .A(n2656), .Z(n2422) );
  HS65_LH_BFX9 U1966 ( .A(n2562), .Z(n2563) );
  HS65_LH_BFX9 U1967 ( .A(n2562), .Z(n2564) );
  HS65_LH_BFX9 U1968 ( .A(b[27]), .Z(n2619) );
  HS65_LH_BFX9 U1969 ( .A(b[2]), .Z(n2569) );
  HS65_LH_BFX9 U1970 ( .A(b[3]), .Z(n2571) );
  HS65_LH_BFX9 U1971 ( .A(n2445), .Z(n2446) );
  HS65_LH_BFX9 U1972 ( .A(n2458), .Z(n2459) );
  HS65_LH_BFX9 U1973 ( .A(n2484), .Z(n2485) );
  HS65_LH_BFX9 U1974 ( .A(n2497), .Z(n2498) );
  HS65_LH_BFX9 U1975 ( .A(n2510), .Z(n2511) );
  HS65_LH_BFX9 U1976 ( .A(n2536), .Z(n2537) );
  HS65_LH_BFX9 U1977 ( .A(n2549), .Z(n2550) );
  HS65_LH_BFX9 U1978 ( .A(b[20]), .Z(n2605) );
  HS65_LH_BFX9 U1979 ( .A(b[11]), .Z(n2587) );
  HS65_LH_BFX9 U1980 ( .A(b[4]), .Z(n2573) );
  HS65_LH_BFX9 U1981 ( .A(b[28]), .Z(n2621) );
  HS65_LH_BFX9 U1982 ( .A(n2471), .Z(n2472) );
  HS65_LH_BFX9 U1983 ( .A(n2523), .Z(n2524) );
  HS65_LH_BFX9 U1984 ( .A(n2433), .Z(n2430) );
  HS65_LH_BFX9 U1985 ( .A(n2433), .Z(n2431) );
  HS65_LH_BFX9 U1986 ( .A(b[31]), .Z(n2627) );
  HS65_LH_BFX9 U1987 ( .A(n2523), .Z(n2525) );
  HS65_LH_BFX9 U1988 ( .A(n2471), .Z(n2473) );
  HS65_LH_BFX9 U1989 ( .A(n2535), .Z(n2533) );
  HS65_LH_BFX9 U1990 ( .A(n2531), .Z(n2529) );
  HS65_LH_BFX9 U1991 ( .A(n2453), .Z(n2451) );
  HS65_LH_BFX9 U1992 ( .A(n2466), .Z(n2464) );
  HS65_LH_BFX9 U1993 ( .A(n2479), .Z(n2477) );
  HS65_LH_BFX9 U1994 ( .A(n2492), .Z(n2490) );
  HS65_LH_BFX9 U1995 ( .A(n2505), .Z(n2503) );
  HS65_LH_BFX9 U1996 ( .A(n2518), .Z(n2516) );
  HS65_LH_BFX9 U1997 ( .A(n2544), .Z(n2542) );
  HS65_LH_BFX9 U1998 ( .A(n2557), .Z(n2555) );
  HS65_LH_BFX9 U1999 ( .A(n2445), .Z(n2447) );
  HS65_LH_BFX9 U2000 ( .A(n2458), .Z(n2460) );
  HS65_LH_BFX9 U2001 ( .A(n2484), .Z(n2486) );
  HS65_LH_BFX9 U2002 ( .A(n2497), .Z(n2499) );
  HS65_LH_BFX9 U2003 ( .A(n2510), .Z(n2512) );
  HS65_LH_BFX9 U2004 ( .A(n2536), .Z(n2538) );
  HS65_LH_BFX9 U2005 ( .A(n2549), .Z(n2551) );
  HS65_LH_BFX9 U2006 ( .A(n2457), .Z(n2454) );
  HS65_LH_BFX9 U2007 ( .A(n2561), .Z(n2558) );
  HS65_LH_BFX9 U2008 ( .A(n2470), .Z(n2467) );
  HS65_LH_BFX9 U2009 ( .A(n2496), .Z(n2493) );
  HS65_LH_BFX9 U2010 ( .A(n2509), .Z(n2506) );
  HS65_LH_BFX9 U2011 ( .A(n2522), .Z(n2519) );
  HS65_LH_BFX9 U2012 ( .A(n2548), .Z(n2545) );
  HS65_LH_BFX9 U2013 ( .A(n2457), .Z(n2455) );
  HS65_LH_BFX9 U2014 ( .A(n2470), .Z(n2468) );
  HS65_LH_BFX9 U2015 ( .A(n2496), .Z(n2494) );
  HS65_LH_BFX9 U2016 ( .A(n2509), .Z(n2507) );
  HS65_LH_BFX9 U2017 ( .A(n2522), .Z(n2520) );
  HS65_LH_BFX9 U2018 ( .A(n2548), .Z(n2546) );
  HS65_LH_BFX9 U2019 ( .A(n2561), .Z(n2559) );
  HS65_LH_BFX9 U2020 ( .A(n2483), .Z(n2480) );
  HS65_LH_BFX9 U2021 ( .A(n2535), .Z(n2532) );
  HS65_LH_BFX9 U2022 ( .A(n2479), .Z(n2476) );
  HS65_LH_BFX9 U2023 ( .A(n2531), .Z(n2528) );
  HS65_LH_BFX9 U2024 ( .A(n2453), .Z(n2450) );
  HS65_LH_BFX9 U2025 ( .A(n2466), .Z(n2463) );
  HS65_LH_BFX9 U2026 ( .A(n2492), .Z(n2489) );
  HS65_LH_BFX9 U2027 ( .A(n2505), .Z(n2502) );
  HS65_LH_BFX9 U2028 ( .A(n2518), .Z(n2515) );
  HS65_LH_BFX9 U2029 ( .A(n2544), .Z(n2541) );
  HS65_LH_BFX9 U2030 ( .A(n2557), .Z(n2554) );
  HS65_LH_BFX9 U2031 ( .A(n2483), .Z(n2481) );
  HS65_LH_IVX9 U2032 ( .A(n2632), .Z(n2631) );
  HS65_LH_IVX9 U2033 ( .A(n2636), .Z(n2635) );
  HS65_LH_IVX9 U2034 ( .A(n31), .Z(n2632) );
  HS65_LH_IVX9 U2035 ( .A(n55), .Z(n2636) );
  HS65_LH_BFX9 U2036 ( .A(n2562), .Z(n2565) );
  HS65_LH_IVX9 U2037 ( .A(n2640), .Z(n2639) );
  HS65_LH_IVX9 U2038 ( .A(n79), .Z(n2640) );
  HS65_LH_IVX9 U2039 ( .A(n2634), .Z(n2633) );
  HS65_LH_IVX9 U2040 ( .A(n43), .Z(n2634) );
  HS65_LH_IVX9 U2041 ( .A(n2644), .Z(n2643) );
  HS65_LH_IVX9 U2042 ( .A(n103), .Z(n2644) );
  HS65_LH_IVX9 U2043 ( .A(n2630), .Z(n2629) );
  HS65_LH_IVX9 U2044 ( .A(n2638), .Z(n2637) );
  HS65_LH_IVX9 U2045 ( .A(n19), .Z(n2630) );
  HS65_LH_IVX9 U2046 ( .A(n67), .Z(n2638) );
  HS65_LH_IVX9 U2047 ( .A(n2646), .Z(n2645) );
  HS65_LH_IVX9 U2048 ( .A(n115), .Z(n2646) );
  HS65_LH_BFX9 U2049 ( .A(n2433), .Z(n2432) );
  HS65_LH_BFX9 U2050 ( .A(n2457), .Z(n2456) );
  HS65_LH_BFX9 U2051 ( .A(n2470), .Z(n2469) );
  HS65_LH_BFX9 U2052 ( .A(n2496), .Z(n2495) );
  HS65_LH_BFX9 U2053 ( .A(n2509), .Z(n2508) );
  HS65_LH_BFX9 U2054 ( .A(n2522), .Z(n2521) );
  HS65_LH_BFX9 U2055 ( .A(n2548), .Z(n2547) );
  HS65_LH_BFX9 U2056 ( .A(n2561), .Z(n2560) );
  HS65_LH_BFX9 U2057 ( .A(n2483), .Z(n2482) );
  HS65_LH_BFX9 U2058 ( .A(n2535), .Z(n2534) );
  HS65_LH_BFX9 U2059 ( .A(n2531), .Z(n2530) );
  HS65_LH_BFX9 U2060 ( .A(n2453), .Z(n2452) );
  HS65_LH_BFX9 U2061 ( .A(n2466), .Z(n2465) );
  HS65_LH_BFX9 U2062 ( .A(n2479), .Z(n2478) );
  HS65_LH_BFX9 U2063 ( .A(n2492), .Z(n2491) );
  HS65_LH_BFX9 U2064 ( .A(n2505), .Z(n2504) );
  HS65_LH_BFX9 U2065 ( .A(n2518), .Z(n2517) );
  HS65_LH_BFX9 U2066 ( .A(n2544), .Z(n2543) );
  HS65_LH_BFX9 U2067 ( .A(n2557), .Z(n2556) );
  HS65_LH_IVX9 U2068 ( .A(n2642), .Z(n2641) );
  HS65_LH_IVX9 U2069 ( .A(n91), .Z(n2642) );
  HS65_LH_IVX9 U2070 ( .A(n2449), .Z(n2448) );
  HS65_LH_IVX9 U2071 ( .A(n2462), .Z(n2461) );
  HS65_LH_IVX9 U2072 ( .A(n2475), .Z(n2474) );
  HS65_LH_IVX9 U2073 ( .A(n2488), .Z(n2487) );
  HS65_LH_IVX9 U2074 ( .A(n2501), .Z(n2500) );
  HS65_LH_IVX9 U2075 ( .A(n2514), .Z(n2513) );
  HS65_LH_IVX9 U2076 ( .A(n2527), .Z(n2526) );
  HS65_LH_IVX9 U2077 ( .A(n2540), .Z(n2539) );
  HS65_LH_IVX9 U2078 ( .A(n2553), .Z(n2552) );
  HS65_LH_IVX9 U2079 ( .A(n2662), .Z(n2655) );
  HS65_LH_IVX9 U2080 ( .A(n2702), .Z(n2656) );
  HS65_LH_BFX9 U2081 ( .A(n2712), .Z(n2457) );
  HS65_LH_BFX9 U2082 ( .A(n3056), .Z(n2561) );
  HS65_LH_BFX9 U2083 ( .A(n2755), .Z(n2470) );
  HS65_LH_BFX9 U2084 ( .A(n2798), .Z(n2483) );
  HS65_LH_BFX9 U2085 ( .A(n2841), .Z(n2496) );
  HS65_LH_BFX9 U2086 ( .A(n2884), .Z(n2509) );
  HS65_LH_BFX9 U2087 ( .A(n2927), .Z(n2522) );
  HS65_LH_BFX9 U2088 ( .A(n2970), .Z(n2535) );
  HS65_LH_BFX9 U2089 ( .A(n3013), .Z(n2548) );
  HS65_LH_BFX9 U2090 ( .A(n2710), .Z(n2453) );
  HS65_LH_BFX9 U2091 ( .A(n2753), .Z(n2466) );
  HS65_LH_BFX9 U2092 ( .A(n2839), .Z(n2492) );
  HS65_LH_BFX9 U2093 ( .A(n2882), .Z(n2505) );
  HS65_LH_BFX9 U2094 ( .A(n2925), .Z(n2518) );
  HS65_LH_BFX9 U2095 ( .A(n2968), .Z(n2531) );
  HS65_LH_BFX9 U2096 ( .A(n3011), .Z(n2544) );
  HS65_LH_BFX9 U2097 ( .A(n3054), .Z(n2557) );
  HS65_LH_BFX9 U2098 ( .A(n2796), .Z(n2479) );
  HS65_LH_BFX9 U2099 ( .A(n2661), .Z(n2433) );
  HS65_LH_IVX9 U2100 ( .A(n2708), .Z(n2449) );
  HS65_LH_IVX9 U2101 ( .A(n2751), .Z(n2462) );
  HS65_LH_IVX9 U2102 ( .A(n2794), .Z(n2475) );
  HS65_LH_IVX9 U2103 ( .A(n2837), .Z(n2488) );
  HS65_LH_IVX9 U2104 ( .A(n2880), .Z(n2501) );
  HS65_LH_IVX9 U2105 ( .A(n2923), .Z(n2514) );
  HS65_LH_IVX9 U2106 ( .A(n2966), .Z(n2527) );
  HS65_LH_IVX9 U2107 ( .A(n3009), .Z(n2540) );
  HS65_LH_IVX9 U2108 ( .A(n3052), .Z(n2553) );
  HS65_LH_BFX9 U2109 ( .A(b[0]), .Z(n2562) );
  HS65_LH_BFX9 U2110 ( .A(n2707), .Z(n2445) );
  HS65_LH_BFX9 U2111 ( .A(n2793), .Z(n2471) );
  HS65_LH_BFX9 U2112 ( .A(n2750), .Z(n2458) );
  HS65_LH_BFX9 U2113 ( .A(n2836), .Z(n2484) );
  HS65_LH_BFX9 U2114 ( .A(n2879), .Z(n2497) );
  HS65_LH_BFX9 U2115 ( .A(n2922), .Z(n2510) );
  HS65_LH_BFX9 U2116 ( .A(n2965), .Z(n2523) );
  HS65_LH_BFX9 U2117 ( .A(n3008), .Z(n2536) );
  HS65_LH_BFX9 U2118 ( .A(n3051), .Z(n2549) );
  HS65_LH_BFX9 U2119 ( .A(b[1]), .Z(n2566) );
  HS65_LH_BFX9 U2120 ( .A(b[19]), .Z(n2602) );
  HS65_LH_BFX9 U2121 ( .A(b[23]), .Z(n2610) );
  HS65_LH_BFX9 U2122 ( .A(b[25]), .Z(n2614) );
  HS65_LH_BFX9 U2123 ( .A(b[12]), .Z(n2588) );
  HS65_LH_BFX9 U2124 ( .A(b[13]), .Z(n2590) );
  HS65_LH_BFX9 U2125 ( .A(b[24]), .Z(n2612) );
  HS65_LH_BFX9 U2126 ( .A(b[26]), .Z(n2616) );
  HS65_LH_BFX9 U2127 ( .A(b[18]), .Z(n2600) );
  HS65_LH_BFX9 U2128 ( .A(b[5]), .Z(n2574) );
  HS65_LH_BFX9 U2129 ( .A(b[7]), .Z(n2578) );
  HS65_LH_BFX9 U2130 ( .A(b[15]), .Z(n2594) );
  HS65_LH_BFX9 U2131 ( .A(b[9]), .Z(n2582) );
  HS65_LH_BFX9 U2132 ( .A(b[17]), .Z(n2598) );
  HS65_LH_BFX9 U2133 ( .A(b[22]), .Z(n2608) );
  HS65_LH_BFX9 U2134 ( .A(b[21]), .Z(n2606) );
  HS65_LH_BFX9 U2135 ( .A(b[29]), .Z(n2622) );
  HS65_LH_BFX9 U2136 ( .A(b[30]), .Z(n2624) );
  HS65_LH_BFX9 U2137 ( .A(b[16]), .Z(n2596) );
  HS65_LH_BFX9 U2138 ( .A(b[6]), .Z(n2576) );
  HS65_LH_BFX9 U2139 ( .A(b[14]), .Z(n2592) );
  HS65_LH_BFX9 U2140 ( .A(b[8]), .Z(n2580) );
  HS65_LH_BFX9 U2141 ( .A(b[10]), .Z(n2584) );
  HS65_LH_BFX9 U2142 ( .A(n2425), .Z(n2423) );
  HS65_LH_BFX9 U2143 ( .A(b[19]), .Z(n2603) );
  HS65_LH_BFX9 U2144 ( .A(n2425), .Z(n2424) );
  HS65_LH_BFX9 U2145 ( .A(b[23]), .Z(n2611) );
  HS65_LH_BFX9 U2146 ( .A(n2436), .Z(n2434) );
  HS65_LH_BFX9 U2147 ( .A(n2440), .Z(n2437) );
  HS65_LH_BFX9 U2148 ( .A(b[25]), .Z(n2615) );
  HS65_LH_BFX9 U2149 ( .A(b[12]), .Z(n2589) );
  HS65_LH_BFX9 U2150 ( .A(b[13]), .Z(n2591) );
  HS65_LH_BFX9 U2151 ( .A(n2440), .Z(n2438) );
  HS65_LH_BFX9 U2152 ( .A(b[24]), .Z(n2613) );
  HS65_LH_BFX9 U2153 ( .A(b[26]), .Z(n2617) );
  HS65_LH_BFX9 U2154 ( .A(b[18]), .Z(n2601) );
  HS65_LH_BFX9 U2155 ( .A(b[5]), .Z(n2575) );
  HS65_LH_BFX9 U2156 ( .A(b[7]), .Z(n2579) );
  HS65_LH_BFX9 U2157 ( .A(b[15]), .Z(n2595) );
  HS65_LH_BFX9 U2158 ( .A(b[9]), .Z(n2583) );
  HS65_LH_BFX9 U2159 ( .A(b[21]), .Z(n2607) );
  HS65_LH_BFX9 U2160 ( .A(b[17]), .Z(n2599) );
  HS65_LH_BFX9 U2161 ( .A(b[22]), .Z(n2609) );
  HS65_LH_BFX9 U2162 ( .A(b[29]), .Z(n2623) );
  HS65_LH_BFX9 U2163 ( .A(n2436), .Z(n2435) );
  HS65_LH_BFX9 U2164 ( .A(b[1]), .Z(n2567) );
  HS65_LH_BFX9 U2165 ( .A(b[30]), .Z(n2625) );
  HS65_LH_BFX9 U2166 ( .A(b[14]), .Z(n2593) );
  HS65_LH_BFX9 U2167 ( .A(b[6]), .Z(n2577) );
  HS65_LH_BFX9 U2168 ( .A(b[8]), .Z(n2581) );
  HS65_LH_BFX9 U2169 ( .A(b[10]), .Z(n2585) );
  HS65_LH_BFX9 U2170 ( .A(b[16]), .Z(n2597) );
  HS65_LH_BFX9 U2171 ( .A(n2444), .Z(n2441) );
  HS65_LH_BFX9 U2172 ( .A(n2444), .Z(n2442) );
  HS65_LH_BFX9 U2173 ( .A(n2429), .Z(n2426) );
  HS65_LH_BFX9 U2174 ( .A(n2429), .Z(n2427) );
  HS65_LH_BFX9 U2175 ( .A(n2444), .Z(n2443) );
  HS65_LH_BFX9 U2176 ( .A(n2429), .Z(n2428) );
  HS65_LH_BFX9 U2177 ( .A(n2440), .Z(n2439) );
  HS65_LH_BFX9 U2178 ( .A(n2670), .Z(n2444) );
  HS65_LH_BFX9 U2179 ( .A(n2659), .Z(n2425) );
  HS65_LH_BFX9 U2180 ( .A(n2668), .Z(n2440) );
  HS65_LH_BFX9 U2181 ( .A(n2660), .Z(n2429) );
  HS65_LH_BFX9 U2182 ( .A(n2666), .Z(n2436) );
  HS65_LHS_XOR3X2 U2183 ( .A(n292), .B(n227), .C(n2658), .Z(product[63]) );
  HS65_LH_AO22X4 U2184 ( .A(n2627), .B(n2423), .C(n2419), .D(n1006), .Z(n2658)
         );
  HS65_LH_MX41X4 U2185 ( .D0(n1025), .S0(n2419), .D1(n2593), .S1(n2427), .D2(
        n2591), .S2(n2431), .D3(n2589), .S3(n2423), .Z(n419) );
  HS65_LH_MX41X4 U2186 ( .D0(n1019), .S0(n2419), .D1(n2601), .S1(n2423), .D2(
        n2603), .S2(n2430), .D3(n2605), .S3(n2426), .Z(n352) );
  HS65_LH_MX41X4 U2187 ( .D0(n1013), .S0(n2419), .D1(n2613), .S1(n2423), .D2(
        n2615), .S2(n2430), .D3(n2617), .S3(n2426), .Z(n309) );
  HS65_LH_OA12X4 U2188 ( .A(n2662), .B(n2657), .C(n2663), .Z(n292) );
  HS65_LH_OAI22X1 U2189 ( .A(n2625), .B(n2664), .C(n2423), .D(n2664), .Z(n2663) );
  HS65_LH_AND2X4 U2190 ( .A(n2626), .B(n2430), .Z(n2664) );
  HS65_LHS_XOR2X3 U2191 ( .A(n7), .B(n2665), .Z(n1419) );
  HS65_LH_AO22X4 U2192 ( .A(n2565), .B(n2434), .C(n2422), .D(n2564), .Z(n2665)
         );
  HS65_LHS_XOR2X3 U2193 ( .A(n7), .B(n2667), .Z(n1418) );
  HS65_LH_AO222X4 U2194 ( .A(n2564), .B(n2437), .C(n2434), .D(n2566), .E(n2422), .F(n1038), .Z(n2667) );
  HS65_LHS_XOR2X3 U2195 ( .A(n7), .B(n2669), .Z(n1417) );
  HS65_LH_MX41X4 U2196 ( .D0(n1037), .S0(n2422), .D1(n2442), .S1(n2564), .D2(
        n2439), .S2(n2566), .D3(n2569), .S3(n2434), .Z(n2669) );
  HS65_LHS_XOR2X3 U2197 ( .A(n7), .B(n2671), .Z(n1416) );
  HS65_LH_MX41X4 U2198 ( .D0(n1036), .S0(n2421), .D1(n2443), .S1(n2567), .D2(
        n2569), .S2(n2437), .D3(n2571), .S3(n2434), .Z(n2671) );
  HS65_LHS_XOR2X3 U2199 ( .A(n7), .B(n2672), .Z(n1415) );
  HS65_LH_MX41X4 U2200 ( .D0(n1035), .S0(n2422), .D1(n2443), .S1(n2569), .D2(
        n2571), .S2(n2437), .D3(n2573), .S3(n2434), .Z(n2672) );
  HS65_LHS_XOR2X3 U2201 ( .A(n7), .B(n2673), .Z(n1414) );
  HS65_LH_MX41X4 U2202 ( .D0(n1034), .S0(n2422), .D1(n2571), .S1(n2441), .D2(
        n2573), .S2(n2437), .D3(n2575), .S3(n2434), .Z(n2673) );
  HS65_LHS_XOR2X3 U2203 ( .A(n7), .B(n2674), .Z(n1413) );
  HS65_LH_MX41X4 U2204 ( .D0(n1033), .S0(n2421), .D1(n2573), .S1(n2441), .D2(
        n2575), .S2(n2437), .D3(n2577), .S3(n2434), .Z(n2674) );
  HS65_LHS_XOR2X3 U2205 ( .A(n7), .B(n2675), .Z(n1412) );
  HS65_LH_MX41X4 U2206 ( .D0(n1032), .S0(n2421), .D1(n2575), .S1(n2441), .D2(
        n2577), .S2(n2437), .D3(n2579), .S3(n2434), .Z(n2675) );
  HS65_LHS_XOR2X3 U2207 ( .A(n7), .B(n2676), .Z(n1411) );
  HS65_LH_MX41X4 U2208 ( .D0(n1031), .S0(n2421), .D1(n2577), .S1(n2441), .D2(
        n2579), .S2(n2437), .D3(n2581), .S3(n2434), .Z(n2676) );
  HS65_LHS_XOR2X3 U2209 ( .A(n7), .B(n2677), .Z(n1410) );
  HS65_LH_MX41X4 U2210 ( .D0(n1030), .S0(n2421), .D1(n2579), .S1(n2441), .D2(
        n2581), .S2(n2437), .D3(n2583), .S3(n2434), .Z(n2677) );
  HS65_LHS_XOR2X3 U2211 ( .A(n7), .B(n2678), .Z(n1409) );
  HS65_LH_MX41X4 U2212 ( .D0(n1029), .S0(n2421), .D1(n2581), .S1(n2441), .D2(
        n2583), .S2(n2437), .D3(n2585), .S3(n2434), .Z(n2678) );
  HS65_LHS_XOR2X3 U2213 ( .A(n7), .B(n2679), .Z(n1408) );
  HS65_LH_MX41X4 U2214 ( .D0(n1028), .S0(n2421), .D1(n2583), .S1(n2441), .D2(
        n2585), .S2(n2437), .D3(n2587), .S3(n2434), .Z(n2679) );
  HS65_LHS_XOR2X3 U2215 ( .A(n7), .B(n2680), .Z(n1407) );
  HS65_LH_MX41X4 U2216 ( .D0(n1027), .S0(n2421), .D1(n2585), .S1(n2441), .D2(
        n2587), .S2(n2437), .D3(n2435), .S3(n2589), .Z(n2680) );
  HS65_LHS_XOR2X3 U2217 ( .A(n7), .B(n2681), .Z(n1406) );
  HS65_LH_MX41X4 U2218 ( .D0(n1026), .S0(n2421), .D1(n2587), .S1(n2441), .D2(
        n2438), .S2(n2588), .D3(n2435), .S3(n2591), .Z(n2681) );
  HS65_LHS_XOR2X3 U2219 ( .A(n7), .B(n2682), .Z(n1405) );
  HS65_LH_MX41X4 U2220 ( .D0(n2422), .S0(n1025), .D1(n2442), .S1(n2589), .D2(
        n2438), .S2(n2590), .D3(n2435), .S3(n2593), .Z(n2682) );
  HS65_LHS_XOR2X3 U2221 ( .A(n7), .B(n2683), .Z(n1404) );
  HS65_LH_MX41X4 U2222 ( .D0(n1024), .S0(n2421), .D1(n2442), .S1(n2591), .D2(
        n2438), .S2(n2592), .D3(n2595), .S3(n2434), .Z(n2683) );
  HS65_LHS_XOR2X3 U2223 ( .A(n7), .B(n2684), .Z(n1403) );
  HS65_LH_MX41X4 U2224 ( .D0(n1023), .S0(n2421), .D1(n2442), .S1(n2593), .D2(
        n2595), .S2(n2437), .D3(n2597), .S3(n2434), .Z(n2684) );
  HS65_LHS_XOR2X3 U2225 ( .A(n7), .B(n2685), .Z(n1402) );
  HS65_LH_MX41X4 U2226 ( .D0(n1022), .S0(n2420), .D1(n2595), .S1(n2441), .D2(
        n2597), .S2(n2437), .D3(n2599), .S3(n2434), .Z(n2685) );
  HS65_LHS_XOR2X3 U2227 ( .A(n7), .B(n2686), .Z(n1401) );
  HS65_LH_MX41X4 U2228 ( .D0(n1021), .S0(n2420), .D1(n2597), .S1(n2441), .D2(
        n2599), .S2(n2437), .D3(n2435), .S3(n2601), .Z(n2686) );
  HS65_LHS_XOR2X3 U2229 ( .A(n7), .B(n2687), .Z(n1400) );
  HS65_LH_MX41X4 U2230 ( .D0(n1020), .S0(n2420), .D1(n2599), .S1(n2441), .D2(
        n2438), .S2(n2600), .D3(n2435), .S3(n2603), .Z(n2687) );
  HS65_LHS_XOR2X3 U2231 ( .A(n7), .B(n2688), .Z(n1399) );
  HS65_LH_MX41X4 U2232 ( .D0(n2422), .S0(n1019), .D1(n2442), .S1(n2601), .D2(
        n2438), .S2(n2602), .D3(n2435), .S3(n2605), .Z(n2688) );
  HS65_LHS_XOR2X3 U2233 ( .A(n7), .B(n2689), .Z(n1398) );
  HS65_LH_MX41X4 U2234 ( .D0(n1018), .S0(n2420), .D1(n2442), .S1(n2603), .D2(
        n2438), .S2(n2604), .D3(n2607), .S3(n2435), .Z(n2689) );
  HS65_LHS_XOR2X3 U2235 ( .A(n7), .B(n2690), .Z(n1397) );
  HS65_LH_MX41X4 U2236 ( .D0(n1017), .S0(n2420), .D1(n2442), .S1(n2605), .D2(
        n2607), .S2(n2438), .D3(n2609), .S3(n2434), .Z(n2690) );
  HS65_LHS_XOR2X3 U2237 ( .A(n7), .B(n2691), .Z(n1396) );
  HS65_LH_MX41X4 U2238 ( .D0(n1016), .S0(n2420), .D1(n2607), .S1(n2442), .D2(
        n2609), .S2(n2438), .D3(n2611), .S3(n2435), .Z(n2691) );
  HS65_LHS_XOR2X3 U2239 ( .A(n7), .B(n2692), .Z(n1395) );
  HS65_LH_MX41X4 U2240 ( .D0(n1015), .S0(n2421), .D1(n2609), .S1(n2442), .D2(
        n2611), .S2(n2438), .D3(n2435), .S3(n2613), .Z(n2692) );
  HS65_LHS_XOR2X3 U2241 ( .A(n7), .B(n2693), .Z(n1394) );
  HS65_LH_MX41X4 U2242 ( .D0(n1014), .S0(n2420), .D1(n2611), .S1(n2442), .D2(
        n2439), .S2(n2612), .D3(n2435), .S3(n2615), .Z(n2693) );
  HS65_LHS_XOR2X3 U2243 ( .A(n7), .B(n2694), .Z(n1393) );
  HS65_LH_MX41X4 U2244 ( .D0(n2422), .S0(n1013), .D1(n2443), .S1(n2613), .D2(
        n2438), .S2(n2614), .D3(n2435), .S3(n2617), .Z(n2694) );
  HS65_LHS_XOR2X3 U2245 ( .A(n7), .B(n2695), .Z(n1392) );
  HS65_LH_MX41X4 U2246 ( .D0(n1012), .S0(n2420), .D1(n2443), .S1(n2615), .D2(
        n2439), .S2(n2616), .D3(n2619), .S3(n2435), .Z(n2695) );
  HS65_LHS_XOR2X3 U2247 ( .A(n7), .B(n2696), .Z(n1391) );
  HS65_LH_MX41X4 U2248 ( .D0(n1011), .S0(n2420), .D1(n2443), .S1(n2617), .D2(
        n2619), .S2(n2438), .D3(n2621), .S3(n2435), .Z(n2696) );
  HS65_LHS_XOR2X3 U2249 ( .A(n7), .B(n2697), .Z(n1390) );
  HS65_LH_MX41X4 U2250 ( .D0(n1010), .S0(n2420), .D1(n2619), .S1(n2442), .D2(
        n2621), .S2(n2438), .D3(n2623), .S3(n2435), .Z(n2697) );
  HS65_LHS_XOR2X3 U2251 ( .A(n7), .B(n2698), .Z(n1389) );
  HS65_LH_MX41X4 U2252 ( .D0(n1009), .S0(n2420), .D1(n2621), .S1(n2442), .D2(
        n2623), .S2(n2438), .D3(n2625), .S3(n2435), .Z(n2698) );
  HS65_LHS_XOR2X3 U2253 ( .A(n7), .B(n2699), .Z(n1388) );
  HS65_LH_MX41X4 U2254 ( .D0(n1008), .S0(n2420), .D1(n2623), .S1(n2442), .D2(
        n2625), .S2(n2438), .D3(n2435), .S3(n2627), .Z(n2699) );
  HS65_LH_NOR2AX3 U2255 ( .A(a[0]), .B(n2700), .Z(n2666) );
  HS65_LHS_XOR2X3 U2256 ( .A(n7), .B(n2701), .Z(n1387) );
  HS65_LH_OAI12X2 U2257 ( .A(n2657), .B(n2702), .C(n2703), .Z(n2701) );
  HS65_LH_OAI22X1 U2258 ( .A(n2625), .B(n2704), .C(n2441), .D(n2704), .Z(n2703) );
  HS65_LH_AND2X4 U2259 ( .A(n2438), .B(n2626), .Z(n2704) );
  HS65_LH_NOR2AX3 U2260 ( .A(a[1]), .B(a[0]), .Z(n2668) );
  HS65_LHS_XOR2X3 U2261 ( .A(n2628), .B(n2705), .Z(n1386) );
  HS65_LH_AOI22X1 U2262 ( .A(n2422), .B(n1006), .C(n2443), .D(n2627), .Z(n2705) );
  HS65_LH_NOR3AX2 U2263 ( .A(n2700), .B(a[0]), .C(a[1]), .Z(n2670) );
  HS65_LH_NAND2X2 U2264 ( .A(a[0]), .B(n2700), .Z(n2702) );
  HS65_LHS_XOR2X3 U2265 ( .A(n7), .B(a[1]), .Z(n2700) );
  HS65_LHS_XOR2X3 U2266 ( .A(n2629), .B(n2706), .Z(n1384) );
  HS65_LH_AO22X4 U2267 ( .A(n2565), .B(n2446), .C(n2564), .D(n2708), .Z(n2706)
         );
  HS65_LHS_XOR2X3 U2268 ( .A(n2629), .B(n2709), .Z(n1383) );
  HS65_LH_AO222X4 U2269 ( .A(n2567), .B(n2446), .C(n2563), .D(n2450), .E(n1038), .F(n2708), .Z(n2709) );
  HS65_LHS_XOR2X3 U2270 ( .A(n2629), .B(n2711), .Z(n1382) );
  HS65_LH_MX41X4 U2271 ( .D0(n2708), .S0(n1037), .D1(n2455), .S1(n2564), .D2(
        n2450), .S2(n2566), .D3(n2446), .S3(n2569), .Z(n2711) );
  HS65_LHS_XOR2X3 U2272 ( .A(n2629), .B(n2713), .Z(n1381) );
  HS65_LH_MX41X4 U2273 ( .D0(n2448), .S0(n1036), .D1(n2454), .S1(n2567), .D2(
        n2450), .S2(n2568), .D3(n2446), .S3(n2571), .Z(n2713) );
  HS65_LHS_XOR2X3 U2274 ( .A(n2629), .B(n2714), .Z(n1380) );
  HS65_LH_MX41X4 U2275 ( .D0(n2708), .S0(n1035), .D1(n2454), .S1(n2569), .D2(
        n2450), .S2(n2570), .D3(n2446), .S3(n2573), .Z(n2714) );
  HS65_LHS_XOR2X3 U2276 ( .A(n2629), .B(n2715), .Z(n1379) );
  HS65_LH_MX41X4 U2277 ( .D0(n2448), .S0(n1034), .D1(n2454), .S1(n2571), .D2(
        n2450), .S2(n2572), .D3(n2446), .S3(n2575), .Z(n2715) );
  HS65_LHS_XOR2X3 U2278 ( .A(n2629), .B(n2716), .Z(n1378) );
  HS65_LH_MX41X4 U2279 ( .D0(n2708), .S0(n1033), .D1(n2454), .S1(n2573), .D2(
        n2450), .S2(n2574), .D3(n2446), .S3(n2577), .Z(n2716) );
  HS65_LHS_XOR2X3 U2280 ( .A(n19), .B(n2717), .Z(n1377) );
  HS65_LH_MX41X4 U2281 ( .D0(n2708), .S0(n1032), .D1(n2454), .S1(n2575), .D2(
        n2450), .S2(n2576), .D3(n2446), .S3(n2579), .Z(n2717) );
  HS65_LHS_XOR2X3 U2282 ( .A(n2629), .B(n2718), .Z(n1376) );
  HS65_LH_MX41X4 U2283 ( .D0(n2448), .S0(n1031), .D1(n2454), .S1(n2577), .D2(
        n2450), .S2(n2578), .D3(n2446), .S3(n2581), .Z(n2718) );
  HS65_LHS_XOR2X3 U2284 ( .A(n2629), .B(n2719), .Z(n1375) );
  HS65_LH_MX41X4 U2285 ( .D0(n2708), .S0(n1030), .D1(n2454), .S1(n2579), .D2(
        n2451), .S2(n2580), .D3(n2446), .S3(n2583), .Z(n2719) );
  HS65_LHS_XOR2X3 U2286 ( .A(n2629), .B(n2720), .Z(n1374) );
  HS65_LH_MX41X4 U2287 ( .D0(n2708), .S0(n1029), .D1(n2454), .S1(n2581), .D2(
        n2450), .S2(n2582), .D3(n2446), .S3(n2585), .Z(n2720) );
  HS65_LHS_XOR2X3 U2288 ( .A(n2629), .B(n2721), .Z(n1373) );
  HS65_LH_MX41X4 U2289 ( .D0(n2708), .S0(n1028), .D1(n2454), .S1(n2583), .D2(
        n2450), .S2(n2584), .D3(n2446), .S3(n2587), .Z(n2721) );
  HS65_LHS_XOR2X3 U2290 ( .A(n19), .B(n2722), .Z(n1372) );
  HS65_LH_MX41X4 U2291 ( .D0(n2708), .S0(n1027), .D1(n2454), .S1(n2585), .D2(
        n2450), .S2(n2586), .D3(n2446), .S3(n2589), .Z(n2722) );
  HS65_LHS_XOR2X3 U2292 ( .A(n19), .B(n2723), .Z(n1371) );
  HS65_LH_MX41X4 U2293 ( .D0(n2708), .S0(n1026), .D1(n2454), .S1(n2587), .D2(
        n2451), .S2(n2588), .D3(n2446), .S3(n2591), .Z(n2723) );
  HS65_LHS_XOR2X3 U2294 ( .A(n19), .B(n2724), .Z(n1370) );
  HS65_LH_MX41X4 U2295 ( .D0(n2708), .S0(n1025), .D1(n2454), .S1(n2589), .D2(
        n2451), .S2(n2590), .D3(n2446), .S3(n2592), .Z(n2724) );
  HS65_LHS_XOR2X3 U2296 ( .A(n19), .B(n2725), .Z(n1369) );
  HS65_LH_MX41X4 U2297 ( .D0(n2708), .S0(n1024), .D1(n2455), .S1(n2591), .D2(
        n2451), .S2(n2592), .D3(n2446), .S3(n2595), .Z(n2725) );
  HS65_LHS_XOR2X3 U2298 ( .A(n2629), .B(n2726), .Z(n1368) );
  HS65_LH_MX41X4 U2299 ( .D0(n2448), .S0(n1023), .D1(n2455), .S1(n2593), .D2(
        n2451), .S2(n2594), .D3(n2446), .S3(n2597), .Z(n2726) );
  HS65_LHS_XOR2X3 U2300 ( .A(n2629), .B(n2727), .Z(n1367) );
  HS65_LH_MX41X4 U2301 ( .D0(n2448), .S0(n1022), .D1(n2455), .S1(n2595), .D2(
        n2451), .S2(n2596), .D3(n2447), .S3(n2599), .Z(n2727) );
  HS65_LHS_XOR2X3 U2302 ( .A(n19), .B(n2728), .Z(n1366) );
  HS65_LH_MX41X4 U2303 ( .D0(n2448), .S0(n1021), .D1(n2455), .S1(n2597), .D2(
        n2451), .S2(n2598), .D3(n2447), .S3(n2600), .Z(n2728) );
  HS65_LHS_XOR2X3 U2304 ( .A(n2629), .B(n2729), .Z(n1365) );
  HS65_LH_MX41X4 U2305 ( .D0(n2448), .S0(n1020), .D1(n2455), .S1(n2599), .D2(
        n2451), .S2(n2600), .D3(n2447), .S3(n2602), .Z(n2729) );
  HS65_LHS_XOR2X3 U2306 ( .A(n19), .B(n2730), .Z(n1364) );
  HS65_LH_MX41X4 U2307 ( .D0(n2448), .S0(n1019), .D1(n2455), .S1(n2601), .D2(
        n2451), .S2(n2602), .D3(n2447), .S3(n2604), .Z(n2730) );
  HS65_LHS_XOR2X3 U2308 ( .A(n2629), .B(n2731), .Z(n1363) );
  HS65_LH_MX41X4 U2309 ( .D0(n2448), .S0(n1018), .D1(n2455), .S1(n2603), .D2(
        n2451), .S2(n2604), .D3(n2447), .S3(n2607), .Z(n2731) );
  HS65_LHS_XOR2X3 U2310 ( .A(n19), .B(n2732), .Z(n1362) );
  HS65_LH_MX41X4 U2311 ( .D0(n2448), .S0(n1017), .D1(n2455), .S1(n2605), .D2(
        n2451), .S2(n2606), .D3(n2447), .S3(n2609), .Z(n2732) );
  HS65_LHS_XOR2X3 U2312 ( .A(n19), .B(n2733), .Z(n1361) );
  HS65_LH_MX41X4 U2313 ( .D0(n2448), .S0(n1016), .D1(n2455), .S1(n2607), .D2(
        n2451), .S2(n2608), .D3(n2447), .S3(n2611), .Z(n2733) );
  HS65_LHS_XOR2X3 U2314 ( .A(n2629), .B(n2734), .Z(n1360) );
  HS65_LH_MX41X4 U2315 ( .D0(n2448), .S0(n1015), .D1(n2455), .S1(n2609), .D2(
        n2451), .S2(n2610), .D3(n2447), .S3(n2612), .Z(n2734) );
  HS65_LHS_XOR2X3 U2316 ( .A(n2629), .B(n2735), .Z(n1359) );
  HS65_LH_MX41X4 U2317 ( .D0(n2448), .S0(n1014), .D1(n2455), .S1(n2611), .D2(
        n2451), .S2(n2612), .D3(n2447), .S3(n2614), .Z(n2735) );
  HS65_LHS_XOR2X3 U2318 ( .A(n19), .B(n2736), .Z(n1358) );
  HS65_LH_MX41X4 U2319 ( .D0(n2448), .S0(n1013), .D1(n2455), .S1(n2613), .D2(
        n2452), .S2(n2614), .D3(n2447), .S3(n2616), .Z(n2736) );
  HS65_LHS_XOR2X3 U2320 ( .A(n19), .B(n2737), .Z(n1357) );
  HS65_LH_MX41X4 U2321 ( .D0(n2448), .S0(n1012), .D1(n2456), .S1(n2615), .D2(
        n2452), .S2(n2616), .D3(n2447), .S3(n2619), .Z(n2737) );
  HS65_LHS_XOR2X3 U2322 ( .A(n2629), .B(n2738), .Z(n1356) );
  HS65_LH_MX41X4 U2323 ( .D0(n2448), .S0(n1011), .D1(n2456), .S1(n2617), .D2(
        n2452), .S2(n2618), .D3(n2447), .S3(n2621), .Z(n2738) );
  HS65_LHS_XOR2X3 U2324 ( .A(n19), .B(n2739), .Z(n1355) );
  HS65_LH_MX41X4 U2325 ( .D0(n2448), .S0(n1010), .D1(n2456), .S1(n2619), .D2(
        n2452), .S2(n2620), .D3(n2447), .S3(n2623), .Z(n2739) );
  HS65_LHS_XOR2X3 U2326 ( .A(n19), .B(n2740), .Z(n1354) );
  HS65_LH_MX41X4 U2327 ( .D0(n2708), .S0(n1009), .D1(n2456), .S1(n2621), .D2(
        n2452), .S2(n2622), .D3(n2447), .S3(n2624), .Z(n2740) );
  HS65_LHS_XOR2X3 U2328 ( .A(n19), .B(n2741), .Z(n1353) );
  HS65_LH_MX41X4 U2329 ( .D0(n2708), .S0(n1008), .D1(n2456), .S1(n2623), .D2(
        n2450), .S2(n2624), .D3(n2447), .S3(n2627), .Z(n2741) );
  HS65_LH_AND2X4 U2330 ( .A(n2742), .B(n2743), .Z(n2707) );
  HS65_LHS_XOR2X3 U2331 ( .A(n19), .B(n2744), .Z(n1352) );
  HS65_LH_OAI12X2 U2332 ( .A(n2657), .B(n2449), .C(n2745), .Z(n2744) );
  HS65_LH_OAI22X1 U2333 ( .A(n2625), .B(n2746), .C(n2454), .D(n2746), .Z(n2745) );
  HS65_LH_AND2X4 U2334 ( .A(n2450), .B(n2626), .Z(n2746) );
  HS65_LH_NOR2X2 U2335 ( .A(n2742), .B(n2747), .Z(n2710) );
  HS65_LHS_XOR2X3 U2336 ( .A(n2630), .B(n2748), .Z(n1351) );
  HS65_LH_AOI22X1 U2337 ( .A(n2708), .B(n1006), .C(n2456), .D(n2627), .Z(n2748) );
  HS65_LH_NOR3AX2 U2338 ( .A(n2747), .B(n2743), .C(n2742), .Z(n2712) );
  HS65_LHS_XNOR2X3 U2339 ( .A(a[4]), .B(a[3]), .Z(n2747) );
  HS65_LH_NOR2AX3 U2340 ( .A(n2742), .B(n2743), .Z(n2708) );
  HS65_LHS_XNOR2X3 U2341 ( .A(n2629), .B(a[4]), .Z(n2743) );
  HS65_LHS_XOR2X3 U2342 ( .A(n7), .B(a[3]), .Z(n2742) );
  HS65_LHS_XOR2X3 U2343 ( .A(n2631), .B(n2749), .Z(n1349) );
  HS65_LH_AO22X4 U2344 ( .A(n2565), .B(n2459), .C(n2564), .D(n2751), .Z(n2749)
         );
  HS65_LHS_XOR2X3 U2345 ( .A(n2631), .B(n2752), .Z(n1348) );
  HS65_LH_AO222X4 U2346 ( .A(n2567), .B(n2459), .C(n2563), .D(n2463), .E(n1038), .F(n2751), .Z(n2752) );
  HS65_LHS_XOR2X3 U2347 ( .A(n2631), .B(n2754), .Z(n1347) );
  HS65_LH_MX41X4 U2348 ( .D0(n2751), .S0(n1037), .D1(n2468), .S1(n2564), .D2(
        n2463), .S2(n2566), .D3(n2459), .S3(n2569), .Z(n2754) );
  HS65_LHS_XOR2X3 U2349 ( .A(n2631), .B(n2756), .Z(n1346) );
  HS65_LH_MX41X4 U2350 ( .D0(n2461), .S0(n1036), .D1(n2467), .S1(n2566), .D2(
        n2463), .S2(n2568), .D3(n2459), .S3(n2571), .Z(n2756) );
  HS65_LHS_XOR2X3 U2351 ( .A(n2631), .B(n2757), .Z(n1345) );
  HS65_LH_MX41X4 U2352 ( .D0(n2751), .S0(n1035), .D1(n2467), .S1(n2569), .D2(
        n2463), .S2(n2570), .D3(n2459), .S3(n2573), .Z(n2757) );
  HS65_LHS_XOR2X3 U2353 ( .A(n2631), .B(n2758), .Z(n1344) );
  HS65_LH_MX41X4 U2354 ( .D0(n2461), .S0(n1034), .D1(n2467), .S1(n2571), .D2(
        n2463), .S2(n2572), .D3(n2459), .S3(n2575), .Z(n2758) );
  HS65_LHS_XOR2X3 U2355 ( .A(n2631), .B(n2759), .Z(n1343) );
  HS65_LH_MX41X4 U2356 ( .D0(n2751), .S0(n1033), .D1(n2467), .S1(n2573), .D2(
        n2463), .S2(n2574), .D3(n2459), .S3(n2577), .Z(n2759) );
  HS65_LHS_XOR2X3 U2357 ( .A(n31), .B(n2760), .Z(n1342) );
  HS65_LH_MX41X4 U2358 ( .D0(n2751), .S0(n1032), .D1(n2467), .S1(n2575), .D2(
        n2463), .S2(n2576), .D3(n2459), .S3(n2579), .Z(n2760) );
  HS65_LHS_XOR2X3 U2359 ( .A(n2631), .B(n2761), .Z(n1341) );
  HS65_LH_MX41X4 U2360 ( .D0(n2461), .S0(n1031), .D1(n2467), .S1(n2577), .D2(
        n2463), .S2(n2578), .D3(n2459), .S3(n2581), .Z(n2761) );
  HS65_LHS_XOR2X3 U2361 ( .A(n2631), .B(n2762), .Z(n1340) );
  HS65_LH_MX41X4 U2362 ( .D0(n2751), .S0(n1030), .D1(n2467), .S1(n2579), .D2(
        n2464), .S2(n2580), .D3(n2459), .S3(n2583), .Z(n2762) );
  HS65_LHS_XOR2X3 U2363 ( .A(n2631), .B(n2763), .Z(n1339) );
  HS65_LH_MX41X4 U2364 ( .D0(n2751), .S0(n1029), .D1(n2467), .S1(n2581), .D2(
        n2463), .S2(n2582), .D3(n2459), .S3(n2585), .Z(n2763) );
  HS65_LHS_XOR2X3 U2365 ( .A(n2631), .B(n2764), .Z(n1338) );
  HS65_LH_MX41X4 U2366 ( .D0(n2751), .S0(n1028), .D1(n2467), .S1(n2583), .D2(
        n2463), .S2(n2584), .D3(n2459), .S3(n2587), .Z(n2764) );
  HS65_LHS_XOR2X3 U2367 ( .A(n31), .B(n2765), .Z(n1337) );
  HS65_LH_MX41X4 U2368 ( .D0(n2751), .S0(n1027), .D1(n2467), .S1(n2585), .D2(
        n2463), .S2(n2586), .D3(n2459), .S3(n2589), .Z(n2765) );
  HS65_LHS_XOR2X3 U2369 ( .A(n31), .B(n2766), .Z(n1336) );
  HS65_LH_MX41X4 U2370 ( .D0(n2751), .S0(n1026), .D1(n2467), .S1(n2587), .D2(
        n2464), .S2(n2588), .D3(n2459), .S3(n2591), .Z(n2766) );
  HS65_LHS_XOR2X3 U2371 ( .A(n31), .B(n2767), .Z(n1335) );
  HS65_LH_MX41X4 U2372 ( .D0(n2751), .S0(n1025), .D1(n2467), .S1(n2589), .D2(
        n2464), .S2(n2590), .D3(n2459), .S3(n2593), .Z(n2767) );
  HS65_LHS_XOR2X3 U2373 ( .A(n31), .B(n2768), .Z(n1334) );
  HS65_LH_MX41X4 U2374 ( .D0(n2751), .S0(n1024), .D1(n2468), .S1(n2591), .D2(
        n2464), .S2(n2592), .D3(n2459), .S3(n2595), .Z(n2768) );
  HS65_LHS_XOR2X3 U2375 ( .A(n2631), .B(n2769), .Z(n1333) );
  HS65_LH_MX41X4 U2376 ( .D0(n2461), .S0(n1023), .D1(n2468), .S1(n2593), .D2(
        n2464), .S2(n2594), .D3(n2459), .S3(n2597), .Z(n2769) );
  HS65_LHS_XOR2X3 U2377 ( .A(n2631), .B(n2770), .Z(n1332) );
  HS65_LH_MX41X4 U2378 ( .D0(n2461), .S0(n1022), .D1(n2468), .S1(n2595), .D2(
        n2464), .S2(n2596), .D3(n2460), .S3(n2599), .Z(n2770) );
  HS65_LHS_XOR2X3 U2379 ( .A(n31), .B(n2771), .Z(n1331) );
  HS65_LH_MX41X4 U2380 ( .D0(n2461), .S0(n1021), .D1(n2468), .S1(n2597), .D2(
        n2464), .S2(n2598), .D3(n2460), .S3(n2601), .Z(n2771) );
  HS65_LHS_XOR2X3 U2381 ( .A(n2631), .B(n2772), .Z(n1330) );
  HS65_LH_MX41X4 U2382 ( .D0(n2461), .S0(n1020), .D1(n2468), .S1(n2599), .D2(
        n2464), .S2(n2600), .D3(n2460), .S3(n2603), .Z(n2772) );
  HS65_LHS_XOR2X3 U2383 ( .A(n31), .B(n2773), .Z(n1329) );
  HS65_LH_MX41X4 U2384 ( .D0(n2461), .S0(n1019), .D1(n2468), .S1(n2601), .D2(
        n2464), .S2(n2602), .D3(n2460), .S3(n2605), .Z(n2773) );
  HS65_LHS_XOR2X3 U2385 ( .A(n2631), .B(n2774), .Z(n1328) );
  HS65_LH_MX41X4 U2386 ( .D0(n2461), .S0(n1018), .D1(n2468), .S1(n2603), .D2(
        n2464), .S2(n2604), .D3(n2460), .S3(n2607), .Z(n2774) );
  HS65_LHS_XOR2X3 U2387 ( .A(n31), .B(n2775), .Z(n1327) );
  HS65_LH_MX41X4 U2388 ( .D0(n2461), .S0(n1017), .D1(n2468), .S1(n2605), .D2(
        n2464), .S2(n2606), .D3(n2460), .S3(n2609), .Z(n2775) );
  HS65_LHS_XOR2X3 U2389 ( .A(n31), .B(n2776), .Z(n1326) );
  HS65_LH_MX41X4 U2390 ( .D0(n2461), .S0(n1016), .D1(n2468), .S1(n2607), .D2(
        n2464), .S2(n2608), .D3(n2460), .S3(n2611), .Z(n2776) );
  HS65_LHS_XOR2X3 U2391 ( .A(n2631), .B(n2777), .Z(n1325) );
  HS65_LH_MX41X4 U2392 ( .D0(n2461), .S0(n1015), .D1(n2468), .S1(n2609), .D2(
        n2464), .S2(n2610), .D3(n2460), .S3(n2613), .Z(n2777) );
  HS65_LHS_XOR2X3 U2393 ( .A(n2631), .B(n2778), .Z(n1324) );
  HS65_LH_MX41X4 U2394 ( .D0(n2461), .S0(n1014), .D1(n2468), .S1(n2611), .D2(
        n2464), .S2(n2612), .D3(n2460), .S3(n2615), .Z(n2778) );
  HS65_LHS_XOR2X3 U2395 ( .A(n31), .B(n2779), .Z(n1323) );
  HS65_LH_MX41X4 U2396 ( .D0(n2461), .S0(n1013), .D1(n2468), .S1(n2613), .D2(
        n2465), .S2(n2614), .D3(n2460), .S3(n2617), .Z(n2779) );
  HS65_LHS_XOR2X3 U2397 ( .A(n31), .B(n2780), .Z(n1322) );
  HS65_LH_MX41X4 U2398 ( .D0(n2461), .S0(n1012), .D1(n2469), .S1(n2615), .D2(
        n2465), .S2(n2616), .D3(n2460), .S3(n2619), .Z(n2780) );
  HS65_LHS_XOR2X3 U2399 ( .A(n2631), .B(n2781), .Z(n1321) );
  HS65_LH_MX41X4 U2400 ( .D0(n2461), .S0(n1011), .D1(n2469), .S1(n2617), .D2(
        n2465), .S2(n2618), .D3(n2460), .S3(n2621), .Z(n2781) );
  HS65_LHS_XOR2X3 U2401 ( .A(n31), .B(n2782), .Z(n1320) );
  HS65_LH_MX41X4 U2402 ( .D0(n2461), .S0(n1010), .D1(n2469), .S1(n2619), .D2(
        n2465), .S2(n2620), .D3(n2460), .S3(n2623), .Z(n2782) );
  HS65_LHS_XOR2X3 U2403 ( .A(n31), .B(n2783), .Z(n1319) );
  HS65_LH_MX41X4 U2404 ( .D0(n2751), .S0(n1009), .D1(n2469), .S1(n2621), .D2(
        n2465), .S2(n2622), .D3(n2460), .S3(n2624), .Z(n2783) );
  HS65_LHS_XOR2X3 U2405 ( .A(n31), .B(n2784), .Z(n1318) );
  HS65_LH_MX41X4 U2406 ( .D0(n2751), .S0(n1008), .D1(n2469), .S1(n2623), .D2(
        n2463), .S2(n2624), .D3(n2460), .S3(n2627), .Z(n2784) );
  HS65_LH_AND2X4 U2407 ( .A(n2785), .B(n2786), .Z(n2750) );
  HS65_LHS_XOR2X3 U2408 ( .A(n31), .B(n2787), .Z(n1317) );
  HS65_LH_OAI12X2 U2409 ( .A(n2657), .B(n2462), .C(n2788), .Z(n2787) );
  HS65_LH_OAI22X1 U2410 ( .A(n2625), .B(n2789), .C(n2467), .D(n2789), .Z(n2788) );
  HS65_LH_AND2X4 U2411 ( .A(n2463), .B(n2626), .Z(n2789) );
  HS65_LH_NOR2X2 U2412 ( .A(n2785), .B(n2790), .Z(n2753) );
  HS65_LHS_XOR2X3 U2413 ( .A(n2632), .B(n2791), .Z(n1316) );
  HS65_LH_AOI22X1 U2414 ( .A(n2751), .B(n1006), .C(n2469), .D(n2627), .Z(n2791) );
  HS65_LH_NOR3AX2 U2415 ( .A(n2790), .B(n2786), .C(n2785), .Z(n2755) );
  HS65_LHS_XNOR2X3 U2416 ( .A(a[7]), .B(a[6]), .Z(n2790) );
  HS65_LH_NOR2AX3 U2417 ( .A(n2785), .B(n2786), .Z(n2751) );
  HS65_LHS_XNOR2X3 U2418 ( .A(n2631), .B(a[7]), .Z(n2786) );
  HS65_LHS_XOR2X3 U2419 ( .A(n2629), .B(a[6]), .Z(n2785) );
  HS65_LHS_XOR2X3 U2420 ( .A(n2633), .B(n2792), .Z(n1314) );
  HS65_LH_AO22X4 U2421 ( .A(n2565), .B(n2472), .C(n2564), .D(n2794), .Z(n2792)
         );
  HS65_LHS_XOR2X3 U2422 ( .A(n2633), .B(n2795), .Z(n1313) );
  HS65_LH_AO222X4 U2423 ( .A(n2567), .B(n2472), .C(n2563), .D(n2476), .E(n1038), .F(n2794), .Z(n2795) );
  HS65_LHS_XOR2X3 U2424 ( .A(n2633), .B(n2797), .Z(n1312) );
  HS65_LH_MX41X4 U2425 ( .D0(n2794), .S0(n1037), .D1(n2472), .S1(n2569), .D2(
        n2477), .S2(n2566), .D3(n2481), .S3(n2564), .Z(n2797) );
  HS65_LHS_XOR2X3 U2426 ( .A(n2633), .B(n2799), .Z(n1311) );
  HS65_LH_MX41X4 U2427 ( .D0(n2474), .S0(n1036), .D1(n2472), .S1(n2571), .D2(
        n2476), .S2(n2568), .D3(n2480), .S3(n2566), .Z(n2799) );
  HS65_LHS_XOR2X3 U2428 ( .A(n2633), .B(n2800), .Z(n1310) );
  HS65_LH_MX41X4 U2429 ( .D0(n2794), .S0(n1035), .D1(n2472), .S1(n2573), .D2(
        n2476), .S2(n2570), .D3(n2480), .S3(n2569), .Z(n2800) );
  HS65_LHS_XOR2X3 U2430 ( .A(n2633), .B(n2801), .Z(n1309) );
  HS65_LH_MX41X4 U2431 ( .D0(n2474), .S0(n1034), .D1(n2472), .S1(n2575), .D2(
        n2476), .S2(n2572), .D3(n2480), .S3(n2571), .Z(n2801) );
  HS65_LHS_XOR2X3 U2432 ( .A(n2633), .B(n2802), .Z(n1308) );
  HS65_LH_MX41X4 U2433 ( .D0(n2794), .S0(n1033), .D1(n2472), .S1(n2577), .D2(
        n2476), .S2(n2574), .D3(n2480), .S3(n2573), .Z(n2802) );
  HS65_LHS_XOR2X3 U2434 ( .A(n43), .B(n2803), .Z(n1307) );
  HS65_LH_MX41X4 U2435 ( .D0(n2794), .S0(n1032), .D1(n2472), .S1(n2579), .D2(
        n2476), .S2(n2576), .D3(n2480), .S3(n2575), .Z(n2803) );
  HS65_LHS_XOR2X3 U2436 ( .A(n2633), .B(n2804), .Z(n1306) );
  HS65_LH_MX41X4 U2437 ( .D0(n2474), .S0(n1031), .D1(n2472), .S1(n2581), .D2(
        n2476), .S2(n2578), .D3(n2480), .S3(n2577), .Z(n2804) );
  HS65_LHS_XOR2X3 U2438 ( .A(n2633), .B(n2805), .Z(n1305) );
  HS65_LH_MX41X4 U2439 ( .D0(n2794), .S0(n1030), .D1(n2472), .S1(n2583), .D2(
        n2477), .S2(n2580), .D3(n2480), .S3(n2579), .Z(n2805) );
  HS65_LHS_XOR2X3 U2440 ( .A(n2633), .B(n2806), .Z(n1304) );
  HS65_LH_MX41X4 U2441 ( .D0(n2794), .S0(n1029), .D1(n2472), .S1(n2585), .D2(
        n2476), .S2(n2582), .D3(n2480), .S3(n2581), .Z(n2806) );
  HS65_LHS_XOR2X3 U2442 ( .A(n2633), .B(n2807), .Z(n1303) );
  HS65_LH_MX41X4 U2443 ( .D0(n2794), .S0(n1028), .D1(n2472), .S1(n2587), .D2(
        n2477), .S2(n2584), .D3(n2480), .S3(n2583), .Z(n2807) );
  HS65_LHS_XOR2X3 U2444 ( .A(n43), .B(n2808), .Z(n1302) );
  HS65_LH_MX41X4 U2445 ( .D0(n2794), .S0(n1027), .D1(n2472), .S1(n2589), .D2(
        n2477), .S2(n2586), .D3(n2480), .S3(n2585), .Z(n2808) );
  HS65_LHS_XOR2X3 U2446 ( .A(n43), .B(n2809), .Z(n1301) );
  HS65_LH_MX41X4 U2447 ( .D0(n2794), .S0(n1026), .D1(n2472), .S1(n2591), .D2(
        n2477), .S2(n2588), .D3(n2480), .S3(n2587), .Z(n2809) );
  HS65_LHS_XOR2X3 U2448 ( .A(n43), .B(n2810), .Z(n1300) );
  HS65_LH_MX41X4 U2449 ( .D0(n2794), .S0(n1025), .D1(n2472), .S1(n2593), .D2(
        n2477), .S2(n2590), .D3(n2480), .S3(n2589), .Z(n2810) );
  HS65_LHS_XOR2X3 U2450 ( .A(n43), .B(n2811), .Z(n1299) );
  HS65_LH_MX41X4 U2451 ( .D0(n2794), .S0(n1024), .D1(n2476), .S1(n2593), .D2(
        n2473), .S2(n2594), .D3(n2481), .S3(n2591), .Z(n2811) );
  HS65_LHS_XOR2X3 U2452 ( .A(n2633), .B(n2812), .Z(n1298) );
  HS65_LH_MX41X4 U2453 ( .D0(n2474), .S0(n1023), .D1(n2476), .S1(n2595), .D2(
        n2473), .S2(n2596), .D3(n2481), .S3(n2593), .Z(n2812) );
  HS65_LHS_XOR2X3 U2454 ( .A(n2633), .B(n2813), .Z(n1297) );
  HS65_LH_MX41X4 U2455 ( .D0(n2474), .S0(n1022), .D1(n2473), .S1(n2599), .D2(
        n2477), .S2(n2596), .D3(n2481), .S3(n2595), .Z(n2813) );
  HS65_LHS_XOR2X3 U2456 ( .A(n43), .B(n2814), .Z(n1296) );
  HS65_LH_MX41X4 U2457 ( .D0(n2474), .S0(n1021), .D1(n2473), .S1(n2601), .D2(
        n2477), .S2(n2598), .D3(n2481), .S3(n2597), .Z(n2814) );
  HS65_LHS_XOR2X3 U2458 ( .A(n2633), .B(n2815), .Z(n1295) );
  HS65_LH_MX41X4 U2459 ( .D0(n2474), .S0(n1020), .D1(n2472), .S1(n2603), .D2(
        n2477), .S2(n2600), .D3(n2481), .S3(n2599), .Z(n2815) );
  HS65_LHS_XOR2X3 U2460 ( .A(n43), .B(n2816), .Z(n1294) );
  HS65_LH_MX41X4 U2461 ( .D0(n2474), .S0(n1019), .D1(n2473), .S1(n2605), .D2(
        n2477), .S2(n2602), .D3(n2481), .S3(n2601), .Z(n2816) );
  HS65_LHS_XOR2X3 U2462 ( .A(n2633), .B(n2817), .Z(n1293) );
  HS65_LH_MX41X4 U2463 ( .D0(n2474), .S0(n1018), .D1(n2473), .S1(n2607), .D2(
        n2477), .S2(n2604), .D3(n2481), .S3(n2603), .Z(n2817) );
  HS65_LHS_XOR2X3 U2464 ( .A(n43), .B(n2818), .Z(n1292) );
  HS65_LH_MX41X4 U2465 ( .D0(n2474), .S0(n1017), .D1(n2473), .S1(n2609), .D2(
        n2477), .S2(n2606), .D3(n2481), .S3(n2605), .Z(n2818) );
  HS65_LHS_XOR2X3 U2466 ( .A(n43), .B(n2819), .Z(n1291) );
  HS65_LH_MX41X4 U2467 ( .D0(n2474), .S0(n1016), .D1(n2473), .S1(n2611), .D2(
        n2477), .S2(n2608), .D3(n2481), .S3(n2607), .Z(n2819) );
  HS65_LHS_XOR2X3 U2468 ( .A(n2633), .B(n2820), .Z(n1290) );
  HS65_LH_MX41X4 U2469 ( .D0(n2474), .S0(n1015), .D1(n2473), .S1(n2613), .D2(
        n2477), .S2(n2610), .D3(n2481), .S3(n2609), .Z(n2820) );
  HS65_LHS_XOR2X3 U2470 ( .A(n2633), .B(n2821), .Z(n1289) );
  HS65_LH_MX41X4 U2471 ( .D0(n2474), .S0(n1014), .D1(n2473), .S1(n2615), .D2(
        n2478), .S2(n2612), .D3(n2481), .S3(n2611), .Z(n2821) );
  HS65_LHS_XOR2X3 U2472 ( .A(n43), .B(n2822), .Z(n1288) );
  HS65_LH_MX41X4 U2473 ( .D0(n2474), .S0(n1013), .D1(n2473), .S1(n2617), .D2(
        n2478), .S2(n2614), .D3(n2481), .S3(n2613), .Z(n2822) );
  HS65_LHS_XOR2X3 U2474 ( .A(n43), .B(n2823), .Z(n1287) );
  HS65_LH_MX41X4 U2475 ( .D0(n2474), .S0(n1012), .D1(n2473), .S1(n2619), .D2(
        n2478), .S2(n2616), .D3(n2482), .S3(n2615), .Z(n2823) );
  HS65_LHS_XOR2X3 U2476 ( .A(n2633), .B(n2824), .Z(n1286) );
  HS65_LH_MX41X4 U2477 ( .D0(n2474), .S0(n1011), .D1(n2473), .S1(n2621), .D2(
        n2478), .S2(n2618), .D3(n2482), .S3(n2617), .Z(n2824) );
  HS65_LHS_XOR2X3 U2478 ( .A(n43), .B(n2825), .Z(n1285) );
  HS65_LH_MX41X4 U2479 ( .D0(n2474), .S0(n1010), .D1(n2473), .S1(n2623), .D2(
        n2478), .S2(n2620), .D3(n2482), .S3(n2619), .Z(n2825) );
  HS65_LHS_XOR2X3 U2480 ( .A(n43), .B(n2826), .Z(n1284) );
  HS65_LH_MX41X4 U2481 ( .D0(n2794), .S0(n1009), .D1(n2473), .S1(n2624), .D2(
        n2476), .S2(n2622), .D3(n2482), .S3(n2621), .Z(n2826) );
  HS65_LHS_XOR2X3 U2482 ( .A(n43), .B(n2827), .Z(n1283) );
  HS65_LH_MX41X4 U2483 ( .D0(n2794), .S0(n1008), .D1(n2476), .S1(n2624), .D2(
        n2473), .S2(n2626), .D3(n2482), .S3(n2623), .Z(n2827) );
  HS65_LH_AND2X4 U2484 ( .A(n2828), .B(n2829), .Z(n2793) );
  HS65_LHS_XOR2X3 U2485 ( .A(n43), .B(n2830), .Z(n1282) );
  HS65_LH_OAI12X2 U2486 ( .A(n2657), .B(n2475), .C(n2831), .Z(n2830) );
  HS65_LH_OAI22X1 U2487 ( .A(n2625), .B(n2832), .C(n2480), .D(n2832), .Z(n2831) );
  HS65_LH_AND2X4 U2488 ( .A(n2476), .B(n2626), .Z(n2832) );
  HS65_LH_NOR2X2 U2489 ( .A(n2828), .B(n2833), .Z(n2796) );
  HS65_LHS_XOR2X3 U2490 ( .A(n2634), .B(n2834), .Z(n1281) );
  HS65_LH_AOI22X1 U2491 ( .A(n2794), .B(n1006), .C(n2482), .D(n2627), .Z(n2834) );
  HS65_LH_NOR3AX2 U2492 ( .A(n2833), .B(n2829), .C(n2828), .Z(n2798) );
  HS65_LHS_XNOR2X3 U2493 ( .A(a[9]), .B(a[10]), .Z(n2833) );
  HS65_LH_NOR2AX3 U2494 ( .A(n2828), .B(n2829), .Z(n2794) );
  HS65_LHS_XNOR2X3 U2495 ( .A(n2633), .B(a[10]), .Z(n2829) );
  HS65_LHS_XOR2X3 U2496 ( .A(n2631), .B(a[9]), .Z(n2828) );
  HS65_LHS_XOR2X3 U2497 ( .A(n2635), .B(n2835), .Z(n1279) );
  HS65_LH_AO22X4 U2498 ( .A(n2565), .B(n2485), .C(n2564), .D(n2837), .Z(n2835)
         );
  HS65_LHS_XOR2X3 U2499 ( .A(n2635), .B(n2838), .Z(n1278) );
  HS65_LH_AO222X4 U2500 ( .A(n2567), .B(n2485), .C(n2563), .D(n2489), .E(n1038), .F(n2837), .Z(n2838) );
  HS65_LHS_XOR2X3 U2501 ( .A(n2635), .B(n2840), .Z(n1277) );
  HS65_LH_MX41X4 U2502 ( .D0(n2837), .S0(n1037), .D1(n2494), .S1(n2563), .D2(
        n2489), .S2(n2566), .D3(n2485), .S3(n2569), .Z(n2840) );
  HS65_LHS_XOR2X3 U2503 ( .A(n2635), .B(n2842), .Z(n1276) );
  HS65_LH_MX41X4 U2504 ( .D0(n2487), .S0(n1036), .D1(n2493), .S1(n2566), .D2(
        n2489), .S2(n2568), .D3(n2485), .S3(n2571), .Z(n2842) );
  HS65_LHS_XOR2X3 U2505 ( .A(n2635), .B(n2843), .Z(n1275) );
  HS65_LH_MX41X4 U2506 ( .D0(n2837), .S0(n1035), .D1(n2493), .S1(n2569), .D2(
        n2489), .S2(n2570), .D3(n2485), .S3(n2573), .Z(n2843) );
  HS65_LHS_XOR2X3 U2507 ( .A(n2635), .B(n2844), .Z(n1274) );
  HS65_LH_MX41X4 U2508 ( .D0(n2487), .S0(n1034), .D1(n2493), .S1(n2571), .D2(
        n2489), .S2(n2572), .D3(n2485), .S3(n2575), .Z(n2844) );
  HS65_LHS_XOR2X3 U2509 ( .A(n2635), .B(n2845), .Z(n1273) );
  HS65_LH_MX41X4 U2510 ( .D0(n2837), .S0(n1033), .D1(n2493), .S1(n2573), .D2(
        n2489), .S2(n2574), .D3(n2485), .S3(n2577), .Z(n2845) );
  HS65_LHS_XOR2X3 U2511 ( .A(n55), .B(n2846), .Z(n1272) );
  HS65_LH_MX41X4 U2512 ( .D0(n2837), .S0(n1032), .D1(n2493), .S1(n2575), .D2(
        n2489), .S2(n2576), .D3(n2485), .S3(n2579), .Z(n2846) );
  HS65_LHS_XOR2X3 U2513 ( .A(n2635), .B(n2847), .Z(n1271) );
  HS65_LH_MX41X4 U2514 ( .D0(n2487), .S0(n1031), .D1(n2493), .S1(n2577), .D2(
        n2489), .S2(n2578), .D3(n2485), .S3(n2581), .Z(n2847) );
  HS65_LHS_XOR2X3 U2515 ( .A(n2635), .B(n2848), .Z(n1270) );
  HS65_LH_MX41X4 U2516 ( .D0(n2837), .S0(n1030), .D1(n2493), .S1(n2579), .D2(
        n2490), .S2(n2580), .D3(n2485), .S3(n2583), .Z(n2848) );
  HS65_LHS_XOR2X3 U2517 ( .A(n2635), .B(n2849), .Z(n1269) );
  HS65_LH_MX41X4 U2518 ( .D0(n2837), .S0(n1029), .D1(n2493), .S1(n2581), .D2(
        n2489), .S2(n2582), .D3(n2485), .S3(n2585), .Z(n2849) );
  HS65_LHS_XOR2X3 U2519 ( .A(n2635), .B(n2850), .Z(n1268) );
  HS65_LH_MX41X4 U2520 ( .D0(n2837), .S0(n1028), .D1(n2493), .S1(n2583), .D2(
        n2489), .S2(n2584), .D3(n2485), .S3(n2587), .Z(n2850) );
  HS65_LHS_XOR2X3 U2521 ( .A(n55), .B(n2851), .Z(n1267) );
  HS65_LH_MX41X4 U2522 ( .D0(n2837), .S0(n1027), .D1(n2493), .S1(n2585), .D2(
        n2489), .S2(n2586), .D3(n2485), .S3(n2589), .Z(n2851) );
  HS65_LHS_XOR2X3 U2523 ( .A(n55), .B(n2852), .Z(n1266) );
  HS65_LH_MX41X4 U2524 ( .D0(n2837), .S0(n1026), .D1(n2493), .S1(n2587), .D2(
        n2490), .S2(n2588), .D3(n2485), .S3(n2591), .Z(n2852) );
  HS65_LHS_XOR2X3 U2525 ( .A(n55), .B(n2853), .Z(n1265) );
  HS65_LH_MX41X4 U2526 ( .D0(n2837), .S0(n1025), .D1(n2493), .S1(n2589), .D2(
        n2490), .S2(n2590), .D3(n2485), .S3(n2593), .Z(n2853) );
  HS65_LHS_XOR2X3 U2527 ( .A(n55), .B(n2854), .Z(n1264) );
  HS65_LH_MX41X4 U2528 ( .D0(n2837), .S0(n1024), .D1(n2494), .S1(n2591), .D2(
        n2490), .S2(n2592), .D3(n2485), .S3(n2595), .Z(n2854) );
  HS65_LHS_XOR2X3 U2529 ( .A(n2635), .B(n2855), .Z(n1263) );
  HS65_LH_MX41X4 U2530 ( .D0(n2487), .S0(n1023), .D1(n2494), .S1(n2593), .D2(
        n2490), .S2(n2594), .D3(n2485), .S3(n2597), .Z(n2855) );
  HS65_LHS_XOR2X3 U2531 ( .A(n2635), .B(n2856), .Z(n1262) );
  HS65_LH_MX41X4 U2532 ( .D0(n2487), .S0(n1022), .D1(n2494), .S1(n2595), .D2(
        n2490), .S2(n2596), .D3(n2486), .S3(n2599), .Z(n2856) );
  HS65_LHS_XOR2X3 U2533 ( .A(n55), .B(n2857), .Z(n1261) );
  HS65_LH_MX41X4 U2534 ( .D0(n2487), .S0(n1021), .D1(n2494), .S1(n2597), .D2(
        n2490), .S2(n2598), .D3(n2486), .S3(n2601), .Z(n2857) );
  HS65_LHS_XOR2X3 U2535 ( .A(n2635), .B(n2858), .Z(n1260) );
  HS65_LH_MX41X4 U2536 ( .D0(n2487), .S0(n1020), .D1(n2494), .S1(n2599), .D2(
        n2490), .S2(n2600), .D3(n2486), .S3(n2603), .Z(n2858) );
  HS65_LHS_XOR2X3 U2537 ( .A(n55), .B(n2859), .Z(n1259) );
  HS65_LH_MX41X4 U2538 ( .D0(n2487), .S0(n1019), .D1(n2494), .S1(n2601), .D2(
        n2490), .S2(n2602), .D3(n2486), .S3(n2605), .Z(n2859) );
  HS65_LHS_XOR2X3 U2539 ( .A(n2635), .B(n2860), .Z(n1258) );
  HS65_LH_MX41X4 U2540 ( .D0(n2487), .S0(n1018), .D1(n2494), .S1(n2603), .D2(
        n2490), .S2(n2604), .D3(n2486), .S3(n2607), .Z(n2860) );
  HS65_LHS_XOR2X3 U2541 ( .A(n55), .B(n2861), .Z(n1257) );
  HS65_LH_MX41X4 U2542 ( .D0(n2487), .S0(n1017), .D1(n2494), .S1(n2605), .D2(
        n2490), .S2(n2606), .D3(n2486), .S3(n2609), .Z(n2861) );
  HS65_LHS_XOR2X3 U2543 ( .A(n55), .B(n2862), .Z(n1256) );
  HS65_LH_MX41X4 U2544 ( .D0(n2487), .S0(n1016), .D1(n2494), .S1(n2607), .D2(
        n2490), .S2(n2608), .D3(n2486), .S3(n2611), .Z(n2862) );
  HS65_LHS_XOR2X3 U2545 ( .A(n2635), .B(n2863), .Z(n1255) );
  HS65_LH_MX41X4 U2546 ( .D0(n2487), .S0(n1015), .D1(n2494), .S1(n2609), .D2(
        n2490), .S2(n2610), .D3(n2486), .S3(n2613), .Z(n2863) );
  HS65_LHS_XOR2X3 U2547 ( .A(n2635), .B(n2864), .Z(n1254) );
  HS65_LH_MX41X4 U2548 ( .D0(n2487), .S0(n1014), .D1(n2494), .S1(n2611), .D2(
        n2490), .S2(n2612), .D3(n2486), .S3(n2615), .Z(n2864) );
  HS65_LHS_XOR2X3 U2549 ( .A(n55), .B(n2865), .Z(n1253) );
  HS65_LH_MX41X4 U2550 ( .D0(n2487), .S0(n1013), .D1(n2494), .S1(n2613), .D2(
        n2491), .S2(n2614), .D3(n2486), .S3(n2617), .Z(n2865) );
  HS65_LHS_XOR2X3 U2551 ( .A(n55), .B(n2866), .Z(n1252) );
  HS65_LH_MX41X4 U2552 ( .D0(n2487), .S0(n1012), .D1(n2495), .S1(n2615), .D2(
        n2491), .S2(n2616), .D3(n2486), .S3(n2619), .Z(n2866) );
  HS65_LHS_XOR2X3 U2553 ( .A(n2635), .B(n2867), .Z(n1251) );
  HS65_LH_MX41X4 U2554 ( .D0(n2487), .S0(n1011), .D1(n2495), .S1(n2617), .D2(
        n2491), .S2(n2618), .D3(n2486), .S3(n2621), .Z(n2867) );
  HS65_LHS_XOR2X3 U2555 ( .A(n55), .B(n2868), .Z(n1250) );
  HS65_LH_MX41X4 U2556 ( .D0(n2487), .S0(n1010), .D1(n2495), .S1(n2619), .D2(
        n2491), .S2(n2620), .D3(n2486), .S3(n2623), .Z(n2868) );
  HS65_LHS_XOR2X3 U2557 ( .A(n55), .B(n2869), .Z(n1249) );
  HS65_LH_MX41X4 U2558 ( .D0(n2837), .S0(n1009), .D1(n2495), .S1(n2621), .D2(
        n2491), .S2(n2622), .D3(n2486), .S3(n2624), .Z(n2869) );
  HS65_LHS_XOR2X3 U2559 ( .A(n55), .B(n2870), .Z(n1248) );
  HS65_LH_MX41X4 U2560 ( .D0(n2837), .S0(n1008), .D1(n2495), .S1(n2623), .D2(
        n2489), .S2(n2624), .D3(n2486), .S3(n2627), .Z(n2870) );
  HS65_LH_AND2X4 U2561 ( .A(n2871), .B(n2872), .Z(n2836) );
  HS65_LHS_XOR2X3 U2562 ( .A(n55), .B(n2873), .Z(n1247) );
  HS65_LH_OAI12X2 U2563 ( .A(n2657), .B(n2488), .C(n2874), .Z(n2873) );
  HS65_LH_OAI22X1 U2564 ( .A(n2625), .B(n2875), .C(n2493), .D(n2875), .Z(n2874) );
  HS65_LH_AND2X4 U2565 ( .A(n2489), .B(n2626), .Z(n2875) );
  HS65_LH_NOR2X2 U2566 ( .A(n2871), .B(n2876), .Z(n2839) );
  HS65_LHS_XOR2X3 U2567 ( .A(n2636), .B(n2877), .Z(n1246) );
  HS65_LH_AOI22X1 U2568 ( .A(n2837), .B(n1006), .C(n2495), .D(n2627), .Z(n2877) );
  HS65_LH_NOR3AX2 U2569 ( .A(n2876), .B(n2872), .C(n2871), .Z(n2841) );
  HS65_LHS_XNOR2X3 U2570 ( .A(a[13]), .B(a[12]), .Z(n2876) );
  HS65_LH_NOR2AX3 U2571 ( .A(n2871), .B(n2872), .Z(n2837) );
  HS65_LHS_XNOR2X3 U2572 ( .A(n2635), .B(a[13]), .Z(n2872) );
  HS65_LHS_XOR2X3 U2573 ( .A(n2633), .B(a[12]), .Z(n2871) );
  HS65_LHS_XOR2X3 U2574 ( .A(n2637), .B(n2878), .Z(n1244) );
  HS65_LH_AO22X4 U2575 ( .A(n2564), .B(n2498), .C(n2564), .D(n2880), .Z(n2878)
         );
  HS65_LHS_XOR2X3 U2576 ( .A(n2637), .B(n2881), .Z(n1243) );
  HS65_LH_AO222X4 U2577 ( .A(n2567), .B(n2498), .C(n2563), .D(n2502), .E(n1038), .F(n2880), .Z(n2881) );
  HS65_LHS_XOR2X3 U2578 ( .A(n2637), .B(n2883), .Z(n1242) );
  HS65_LH_MX41X4 U2579 ( .D0(n2880), .S0(n1037), .D1(n2507), .S1(n2563), .D2(
        n2502), .S2(n2566), .D3(n2498), .S3(n2569), .Z(n2883) );
  HS65_LHS_XOR2X3 U2580 ( .A(n2637), .B(n2885), .Z(n1241) );
  HS65_LH_MX41X4 U2581 ( .D0(n2500), .S0(n1036), .D1(n2506), .S1(n2566), .D2(
        n2502), .S2(n2568), .D3(n2498), .S3(n2571), .Z(n2885) );
  HS65_LHS_XOR2X3 U2582 ( .A(n2637), .B(n2886), .Z(n1240) );
  HS65_LH_MX41X4 U2583 ( .D0(n2880), .S0(n1035), .D1(n2506), .S1(n2568), .D2(
        n2502), .S2(n2570), .D3(n2498), .S3(n2573), .Z(n2886) );
  HS65_LHS_XOR2X3 U2584 ( .A(n2637), .B(n2887), .Z(n1239) );
  HS65_LH_MX41X4 U2585 ( .D0(n2500), .S0(n1034), .D1(n2506), .S1(n2570), .D2(
        n2502), .S2(n2572), .D3(n2498), .S3(n2575), .Z(n2887) );
  HS65_LHS_XOR2X3 U2586 ( .A(n2637), .B(n2888), .Z(n1238) );
  HS65_LH_MX41X4 U2587 ( .D0(n2880), .S0(n1033), .D1(n2506), .S1(n2572), .D2(
        n2502), .S2(n2574), .D3(n2498), .S3(n2577), .Z(n2888) );
  HS65_LHS_XOR2X3 U2588 ( .A(n67), .B(n2889), .Z(n1237) );
  HS65_LH_MX41X4 U2589 ( .D0(n2880), .S0(n1032), .D1(n2506), .S1(n2574), .D2(
        n2502), .S2(n2576), .D3(n2498), .S3(n2579), .Z(n2889) );
  HS65_LHS_XOR2X3 U2590 ( .A(n2637), .B(n2890), .Z(n1236) );
  HS65_LH_MX41X4 U2591 ( .D0(n2500), .S0(n1031), .D1(n2506), .S1(n2576), .D2(
        n2502), .S2(n2578), .D3(n2498), .S3(n2581), .Z(n2890) );
  HS65_LHS_XOR2X3 U2592 ( .A(n2637), .B(n2891), .Z(n1235) );
  HS65_LH_MX41X4 U2593 ( .D0(n2880), .S0(n1030), .D1(n2506), .S1(n2578), .D2(
        n2503), .S2(n2580), .D3(n2498), .S3(n2583), .Z(n2891) );
  HS65_LHS_XOR2X3 U2594 ( .A(n2637), .B(n2892), .Z(n1234) );
  HS65_LH_MX41X4 U2595 ( .D0(n2880), .S0(n1029), .D1(n2506), .S1(n2580), .D2(
        n2502), .S2(n2582), .D3(n2498), .S3(n2585), .Z(n2892) );
  HS65_LHS_XOR2X3 U2596 ( .A(n2637), .B(n2893), .Z(n1233) );
  HS65_LH_MX41X4 U2597 ( .D0(n2880), .S0(n1028), .D1(n2506), .S1(n2582), .D2(
        n2502), .S2(n2584), .D3(n2498), .S3(n2587), .Z(n2893) );
  HS65_LHS_XOR2X3 U2598 ( .A(n67), .B(n2894), .Z(n1232) );
  HS65_LH_MX41X4 U2599 ( .D0(n2880), .S0(n1027), .D1(n2506), .S1(n2584), .D2(
        n2502), .S2(n2586), .D3(n2498), .S3(n2589), .Z(n2894) );
  HS65_LHS_XOR2X3 U2600 ( .A(n67), .B(n2895), .Z(n1231) );
  HS65_LH_MX41X4 U2601 ( .D0(n2880), .S0(n1026), .D1(n2506), .S1(n2586), .D2(
        n2503), .S2(n2588), .D3(n2498), .S3(n2591), .Z(n2895) );
  HS65_LHS_XOR2X3 U2602 ( .A(n67), .B(n2896), .Z(n1230) );
  HS65_LH_MX41X4 U2603 ( .D0(n2880), .S0(n1025), .D1(n2506), .S1(n2589), .D2(
        n2503), .S2(n2590), .D3(n2498), .S3(n2593), .Z(n2896) );
  HS65_LHS_XOR2X3 U2604 ( .A(n67), .B(n2897), .Z(n1229) );
  HS65_LH_MX41X4 U2605 ( .D0(n2880), .S0(n1024), .D1(n2507), .S1(n2591), .D2(
        n2503), .S2(n2592), .D3(n2498), .S3(n2595), .Z(n2897) );
  HS65_LHS_XOR2X3 U2606 ( .A(n2637), .B(n2898), .Z(n1228) );
  HS65_LH_MX41X4 U2607 ( .D0(n2500), .S0(n1023), .D1(n2507), .S1(n2593), .D2(
        n2503), .S2(n2594), .D3(n2498), .S3(n2597), .Z(n2898) );
  HS65_LHS_XOR2X3 U2608 ( .A(n2637), .B(n2899), .Z(n1227) );
  HS65_LH_MX41X4 U2609 ( .D0(n2500), .S0(n1022), .D1(n2507), .S1(n2594), .D2(
        n2503), .S2(n2596), .D3(n2499), .S3(n2599), .Z(n2899) );
  HS65_LHS_XOR2X3 U2610 ( .A(n67), .B(n2900), .Z(n1226) );
  HS65_LH_MX41X4 U2611 ( .D0(n2500), .S0(n1021), .D1(n2507), .S1(n2597), .D2(
        n2503), .S2(n2598), .D3(n2499), .S3(n2601), .Z(n2900) );
  HS65_LHS_XOR2X3 U2612 ( .A(n2637), .B(n2901), .Z(n1225) );
  HS65_LH_MX41X4 U2613 ( .D0(n2500), .S0(n1020), .D1(n2507), .S1(n2598), .D2(
        n2503), .S2(n2600), .D3(n2499), .S3(n2603), .Z(n2901) );
  HS65_LHS_XOR2X3 U2614 ( .A(n67), .B(n2902), .Z(n1224) );
  HS65_LH_MX41X4 U2615 ( .D0(n2500), .S0(n1019), .D1(n2507), .S1(n2601), .D2(
        n2503), .S2(n2602), .D3(n2499), .S3(n2605), .Z(n2902) );
  HS65_LHS_XOR2X3 U2616 ( .A(n2637), .B(n2903), .Z(n1223) );
  HS65_LH_MX41X4 U2617 ( .D0(n2500), .S0(n1018), .D1(n2507), .S1(n2603), .D2(
        n2503), .S2(n2604), .D3(n2499), .S3(n2607), .Z(n2903) );
  HS65_LHS_XOR2X3 U2618 ( .A(n67), .B(n2904), .Z(n1222) );
  HS65_LH_MX41X4 U2619 ( .D0(n2500), .S0(n1017), .D1(n2507), .S1(n2605), .D2(
        n2503), .S2(n2606), .D3(n2499), .S3(n2609), .Z(n2904) );
  HS65_LHS_XOR2X3 U2620 ( .A(n67), .B(n2905), .Z(n1221) );
  HS65_LH_MX41X4 U2621 ( .D0(n2500), .S0(n1016), .D1(n2507), .S1(n2606), .D2(
        n2503), .S2(n2608), .D3(n2499), .S3(n2611), .Z(n2905) );
  HS65_LHS_XOR2X3 U2622 ( .A(n2637), .B(n2906), .Z(n1220) );
  HS65_LH_MX41X4 U2623 ( .D0(n2500), .S0(n1015), .D1(n2507), .S1(n2608), .D2(
        n2503), .S2(n2610), .D3(n2499), .S3(n2613), .Z(n2906) );
  HS65_LHS_XOR2X3 U2624 ( .A(n2637), .B(n2907), .Z(n1219) );
  HS65_LH_MX41X4 U2625 ( .D0(n2500), .S0(n1014), .D1(n2507), .S1(n2610), .D2(
        n2503), .S2(n2612), .D3(n2499), .S3(n2615), .Z(n2907) );
  HS65_LHS_XOR2X3 U2626 ( .A(n67), .B(n2908), .Z(n1218) );
  HS65_LH_MX41X4 U2627 ( .D0(n2500), .S0(n1013), .D1(n2507), .S1(n2613), .D2(
        n2504), .S2(n2614), .D3(n2499), .S3(n2617), .Z(n2908) );
  HS65_LHS_XOR2X3 U2628 ( .A(n67), .B(n2909), .Z(n1217) );
  HS65_LH_MX41X4 U2629 ( .D0(n2500), .S0(n1012), .D1(n2508), .S1(n2615), .D2(
        n2504), .S2(n2616), .D3(n2499), .S3(n2619), .Z(n2909) );
  HS65_LHS_XOR2X3 U2630 ( .A(n2637), .B(n2910), .Z(n1216) );
  HS65_LH_MX41X4 U2631 ( .D0(n2500), .S0(n1011), .D1(n2508), .S1(n2617), .D2(
        n2504), .S2(n2618), .D3(n2499), .S3(n2621), .Z(n2910) );
  HS65_LHS_XOR2X3 U2632 ( .A(n67), .B(n2911), .Z(n1215) );
  HS65_LH_MX41X4 U2633 ( .D0(n2500), .S0(n1010), .D1(n2508), .S1(n2618), .D2(
        n2504), .S2(n2620), .D3(n2499), .S3(n2623), .Z(n2911) );
  HS65_LHS_XOR2X3 U2634 ( .A(n67), .B(n2912), .Z(n1214) );
  HS65_LH_MX41X4 U2635 ( .D0(n2880), .S0(n1009), .D1(n2508), .S1(n2620), .D2(
        n2504), .S2(n2622), .D3(n2499), .S3(n2624), .Z(n2912) );
  HS65_LHS_XOR2X3 U2636 ( .A(n67), .B(n2913), .Z(n1213) );
  HS65_LH_MX41X4 U2637 ( .D0(n2880), .S0(n1008), .D1(n2508), .S1(n2622), .D2(
        n2502), .S2(n2624), .D3(n2499), .S3(n2626), .Z(n2913) );
  HS65_LH_AND2X4 U2638 ( .A(n2914), .B(n2915), .Z(n2879) );
  HS65_LHS_XOR2X3 U2639 ( .A(n67), .B(n2916), .Z(n1212) );
  HS65_LH_OAI12X2 U2640 ( .A(n2657), .B(n2501), .C(n2917), .Z(n2916) );
  HS65_LH_OAI22X1 U2641 ( .A(n2625), .B(n2918), .C(n2506), .D(n2918), .Z(n2917) );
  HS65_LH_AND2X4 U2642 ( .A(n2502), .B(n2626), .Z(n2918) );
  HS65_LH_NOR2X2 U2643 ( .A(n2914), .B(n2919), .Z(n2882) );
  HS65_LHS_XOR2X3 U2644 ( .A(n2638), .B(n2920), .Z(n1211) );
  HS65_LH_AOI22X1 U2645 ( .A(n2880), .B(n1006), .C(n2508), .D(n2627), .Z(n2920) );
  HS65_LH_NOR3AX2 U2646 ( .A(n2919), .B(n2915), .C(n2914), .Z(n2884) );
  HS65_LHS_XNOR2X3 U2647 ( .A(a[16]), .B(a[15]), .Z(n2919) );
  HS65_LH_NOR2AX3 U2648 ( .A(n2914), .B(n2915), .Z(n2880) );
  HS65_LHS_XNOR2X3 U2649 ( .A(n2637), .B(a[16]), .Z(n2915) );
  HS65_LHS_XOR2X3 U2650 ( .A(n2635), .B(a[15]), .Z(n2914) );
  HS65_LHS_XOR2X3 U2651 ( .A(n2639), .B(n2921), .Z(n1209) );
  HS65_LH_AO22X4 U2652 ( .A(n2565), .B(n2511), .C(n2564), .D(n2923), .Z(n2921)
         );
  HS65_LHS_XOR2X3 U2653 ( .A(n2639), .B(n2924), .Z(n1208) );
  HS65_LH_AO222X4 U2654 ( .A(n2567), .B(n2511), .C(n2563), .D(n2515), .E(n1038), .F(n2923), .Z(n2924) );
  HS65_LHS_XOR2X3 U2655 ( .A(n2639), .B(n2926), .Z(n1207) );
  HS65_LH_MX41X4 U2656 ( .D0(n2923), .S0(n1037), .D1(n2520), .S1(n2564), .D2(
        n2515), .S2(n2566), .D3(n2511), .S3(n2568), .Z(n2926) );
  HS65_LHS_XOR2X3 U2657 ( .A(n2639), .B(n2928), .Z(n1206) );
  HS65_LH_MX41X4 U2658 ( .D0(n2513), .S0(n1036), .D1(n2519), .S1(n2566), .D2(
        n2515), .S2(n2568), .D3(n2511), .S3(n2570), .Z(n2928) );
  HS65_LHS_XOR2X3 U2659 ( .A(n2639), .B(n2929), .Z(n1205) );
  HS65_LH_MX41X4 U2660 ( .D0(n2923), .S0(n1035), .D1(n2519), .S1(n2568), .D2(
        n2515), .S2(n2570), .D3(n2511), .S3(n2572), .Z(n2929) );
  HS65_LHS_XOR2X3 U2661 ( .A(n2639), .B(n2930), .Z(n1204) );
  HS65_LH_MX41X4 U2662 ( .D0(n2513), .S0(n1034), .D1(n2519), .S1(n2570), .D2(
        n2515), .S2(n2572), .D3(n2511), .S3(n2574), .Z(n2930) );
  HS65_LHS_XOR2X3 U2663 ( .A(n2639), .B(n2931), .Z(n1203) );
  HS65_LH_MX41X4 U2664 ( .D0(n2923), .S0(n1033), .D1(n2519), .S1(n2572), .D2(
        n2515), .S2(n2574), .D3(n2511), .S3(n2576), .Z(n2931) );
  HS65_LHS_XOR2X3 U2665 ( .A(n79), .B(n2932), .Z(n1202) );
  HS65_LH_MX41X4 U2666 ( .D0(n2923), .S0(n1032), .D1(n2519), .S1(n2574), .D2(
        n2515), .S2(n2576), .D3(n2511), .S3(n2578), .Z(n2932) );
  HS65_LHS_XOR2X3 U2667 ( .A(n2639), .B(n2933), .Z(n1201) );
  HS65_LH_MX41X4 U2668 ( .D0(n2513), .S0(n1031), .D1(n2519), .S1(n2576), .D2(
        n2515), .S2(n2578), .D3(n2511), .S3(n2580), .Z(n2933) );
  HS65_LHS_XOR2X3 U2669 ( .A(n2639), .B(n2934), .Z(n1200) );
  HS65_LH_MX41X4 U2670 ( .D0(n2923), .S0(n1030), .D1(n2519), .S1(n2578), .D2(
        n2516), .S2(n2580), .D3(n2511), .S3(n2582), .Z(n2934) );
  HS65_LHS_XOR2X3 U2671 ( .A(n2639), .B(n2935), .Z(n1199) );
  HS65_LH_MX41X4 U2672 ( .D0(n2923), .S0(n1029), .D1(n2519), .S1(n2580), .D2(
        n2515), .S2(n2582), .D3(n2511), .S3(n2584), .Z(n2935) );
  HS65_LHS_XOR2X3 U2673 ( .A(n2639), .B(n2936), .Z(n1198) );
  HS65_LH_MX41X4 U2674 ( .D0(n2923), .S0(n1028), .D1(n2519), .S1(n2582), .D2(
        n2515), .S2(n2584), .D3(n2511), .S3(n2586), .Z(n2936) );
  HS65_LHS_XOR2X3 U2675 ( .A(n79), .B(n2937), .Z(n1197) );
  HS65_LH_MX41X4 U2676 ( .D0(n2923), .S0(n1027), .D1(n2519), .S1(n2584), .D2(
        n2515), .S2(n2586), .D3(n2511), .S3(n2589), .Z(n2937) );
  HS65_LHS_XOR2X3 U2677 ( .A(n79), .B(n2938), .Z(n1196) );
  HS65_LH_MX41X4 U2678 ( .D0(n2923), .S0(n1026), .D1(n2519), .S1(n2586), .D2(
        n2516), .S2(n2588), .D3(n2511), .S3(n2591), .Z(n2938) );
  HS65_LHS_XOR2X3 U2679 ( .A(n79), .B(n2939), .Z(n1195) );
  HS65_LH_MX41X4 U2680 ( .D0(n2923), .S0(n1025), .D1(n2519), .S1(n2588), .D2(
        n2516), .S2(n2590), .D3(n2511), .S3(n2592), .Z(n2939) );
  HS65_LHS_XOR2X3 U2681 ( .A(n79), .B(n2940), .Z(n1194) );
  HS65_LH_MX41X4 U2682 ( .D0(n2923), .S0(n1024), .D1(n2520), .S1(n2590), .D2(
        n2516), .S2(n2592), .D3(n2511), .S3(n2594), .Z(n2940) );
  HS65_LHS_XOR2X3 U2683 ( .A(n2639), .B(n2941), .Z(n1193) );
  HS65_LH_MX41X4 U2684 ( .D0(n2513), .S0(n1023), .D1(n2520), .S1(n2592), .D2(
        n2516), .S2(n2594), .D3(n2511), .S3(n2596), .Z(n2941) );
  HS65_LHS_XOR2X3 U2685 ( .A(n2639), .B(n2942), .Z(n1192) );
  HS65_LH_MX41X4 U2686 ( .D0(n2513), .S0(n1022), .D1(n2520), .S1(n2594), .D2(
        n2516), .S2(n2596), .D3(n2512), .S3(n2598), .Z(n2942) );
  HS65_LHS_XOR2X3 U2687 ( .A(n79), .B(n2943), .Z(n1191) );
  HS65_LH_MX41X4 U2688 ( .D0(n2513), .S0(n1021), .D1(n2520), .S1(n2596), .D2(
        n2516), .S2(n2598), .D3(n2512), .S3(n2601), .Z(n2943) );
  HS65_LHS_XOR2X3 U2689 ( .A(n2639), .B(n2944), .Z(n1190) );
  HS65_LH_MX41X4 U2690 ( .D0(n2513), .S0(n1020), .D1(n2520), .S1(n2598), .D2(
        n2516), .S2(n2600), .D3(n2512), .S3(n2603), .Z(n2944) );
  HS65_LHS_XOR2X3 U2691 ( .A(n79), .B(n2945), .Z(n1189) );
  HS65_LH_MX41X4 U2692 ( .D0(n2513), .S0(n1019), .D1(n2520), .S1(n2600), .D2(
        n2516), .S2(n2602), .D3(n2512), .S3(n2605), .Z(n2945) );
  HS65_LHS_XOR2X3 U2693 ( .A(n2639), .B(n2946), .Z(n1188) );
  HS65_LH_MX41X4 U2694 ( .D0(n2513), .S0(n1018), .D1(n2520), .S1(n2602), .D2(
        n2516), .S2(n2604), .D3(n2512), .S3(n2606), .Z(n2946) );
  HS65_LHS_XOR2X3 U2695 ( .A(n79), .B(n2947), .Z(n1187) );
  HS65_LH_MX41X4 U2696 ( .D0(n2513), .S0(n1017), .D1(n2520), .S1(n2604), .D2(
        n2516), .S2(n2606), .D3(n2512), .S3(n2608), .Z(n2947) );
  HS65_LHS_XOR2X3 U2697 ( .A(n79), .B(n2948), .Z(n1186) );
  HS65_LH_MX41X4 U2698 ( .D0(n2513), .S0(n1016), .D1(n2520), .S1(n2606), .D2(
        n2516), .S2(n2608), .D3(n2512), .S3(n2610), .Z(n2948) );
  HS65_LHS_XOR2X3 U2699 ( .A(n2639), .B(n2949), .Z(n1185) );
  HS65_LH_MX41X4 U2700 ( .D0(n2513), .S0(n1015), .D1(n2520), .S1(n2608), .D2(
        n2516), .S2(n2610), .D3(n2512), .S3(n2613), .Z(n2949) );
  HS65_LHS_XOR2X3 U2701 ( .A(n2639), .B(n2950), .Z(n1184) );
  HS65_LH_MX41X4 U2702 ( .D0(n2513), .S0(n1014), .D1(n2520), .S1(n2610), .D2(
        n2516), .S2(n2612), .D3(n2512), .S3(n2615), .Z(n2950) );
  HS65_LHS_XOR2X3 U2703 ( .A(n79), .B(n2951), .Z(n1183) );
  HS65_LH_MX41X4 U2704 ( .D0(n2513), .S0(n1013), .D1(n2520), .S1(n2612), .D2(
        n2517), .S2(n2614), .D3(n2512), .S3(n2617), .Z(n2951) );
  HS65_LHS_XOR2X3 U2705 ( .A(n79), .B(n2952), .Z(n1182) );
  HS65_LH_MX41X4 U2706 ( .D0(n2513), .S0(n1012), .D1(n2521), .S1(n2614), .D2(
        n2517), .S2(n2616), .D3(n2512), .S3(n2618), .Z(n2952) );
  HS65_LHS_XOR2X3 U2707 ( .A(n2639), .B(n2953), .Z(n1181) );
  HS65_LH_MX41X4 U2708 ( .D0(n2513), .S0(n1011), .D1(n2521), .S1(n2616), .D2(
        n2517), .S2(n2618), .D3(n2512), .S3(n2620), .Z(n2953) );
  HS65_LHS_XOR2X3 U2709 ( .A(n79), .B(n2954), .Z(n1180) );
  HS65_LH_MX41X4 U2710 ( .D0(n2513), .S0(n1010), .D1(n2521), .S1(n2618), .D2(
        n2517), .S2(n2620), .D3(n2512), .S3(n2622), .Z(n2954) );
  HS65_LHS_XOR2X3 U2711 ( .A(n79), .B(n2955), .Z(n1179) );
  HS65_LH_MX41X4 U2712 ( .D0(n2923), .S0(n1009), .D1(n2521), .S1(n2620), .D2(
        n2517), .S2(n2622), .D3(n2512), .S3(n2624), .Z(n2955) );
  HS65_LHS_XOR2X3 U2713 ( .A(n79), .B(n2956), .Z(n1178) );
  HS65_LH_MX41X4 U2714 ( .D0(n2923), .S0(n1008), .D1(n2521), .S1(n2622), .D2(
        n2515), .S2(n2624), .D3(n2512), .S3(n2626), .Z(n2956) );
  HS65_LH_AND2X4 U2715 ( .A(n2957), .B(n2958), .Z(n2922) );
  HS65_LHS_XOR2X3 U2716 ( .A(n79), .B(n2959), .Z(n1177) );
  HS65_LH_OAI12X2 U2717 ( .A(n2657), .B(n2514), .C(n2960), .Z(n2959) );
  HS65_LH_OAI22X1 U2718 ( .A(n2625), .B(n2961), .C(n2519), .D(n2961), .Z(n2960) );
  HS65_LH_AND2X4 U2719 ( .A(n2515), .B(n2626), .Z(n2961) );
  HS65_LH_NOR2X2 U2720 ( .A(n2957), .B(n2962), .Z(n2925) );
  HS65_LHS_XOR2X3 U2721 ( .A(n2640), .B(n2963), .Z(n1176) );
  HS65_LH_AOI22X1 U2722 ( .A(n2923), .B(n1006), .C(n2521), .D(n2627), .Z(n2963) );
  HS65_LH_NOR3AX2 U2723 ( .A(n2962), .B(n2958), .C(n2957), .Z(n2927) );
  HS65_LHS_XNOR2X3 U2724 ( .A(a[19]), .B(a[18]), .Z(n2962) );
  HS65_LH_NOR2AX3 U2725 ( .A(n2957), .B(n2958), .Z(n2923) );
  HS65_LHS_XNOR2X3 U2726 ( .A(n2639), .B(a[19]), .Z(n2958) );
  HS65_LHS_XOR2X3 U2727 ( .A(n2637), .B(a[18]), .Z(n2957) );
  HS65_LHS_XOR2X3 U2728 ( .A(n2641), .B(n2964), .Z(n1174) );
  HS65_LH_AO22X4 U2729 ( .A(n2565), .B(n2524), .C(n2564), .D(n2966), .Z(n2964)
         );
  HS65_LHS_XOR2X3 U2730 ( .A(n2641), .B(n2967), .Z(n1173) );
  HS65_LH_AO222X4 U2731 ( .A(n2567), .B(n2524), .C(n2563), .D(n2528), .E(n1038), .F(n2966), .Z(n2967) );
  HS65_LHS_XOR2X3 U2732 ( .A(n2641), .B(n2969), .Z(n1172) );
  HS65_LH_MX41X4 U2733 ( .D0(n2966), .S0(n1037), .D1(n2524), .S1(n2568), .D2(
        n2533), .S2(n2563), .D3(n2528), .S3(n2566), .Z(n2969) );
  HS65_LHS_XOR2X3 U2734 ( .A(n2641), .B(n2971), .Z(n1171) );
  HS65_LH_MX41X4 U2735 ( .D0(n2526), .S0(n1036), .D1(n2524), .S1(n2570), .D2(
        n2532), .S2(n2566), .D3(n2528), .S3(n2568), .Z(n2971) );
  HS65_LHS_XOR2X3 U2736 ( .A(n2641), .B(n2972), .Z(n1170) );
  HS65_LH_MX41X4 U2737 ( .D0(n2966), .S0(n1035), .D1(n2524), .S1(n2572), .D2(
        n2532), .S2(n2568), .D3(n2528), .S3(n2570), .Z(n2972) );
  HS65_LHS_XOR2X3 U2738 ( .A(n2641), .B(n2973), .Z(n1169) );
  HS65_LH_MX41X4 U2739 ( .D0(n2526), .S0(n1034), .D1(n2524), .S1(n2574), .D2(
        n2532), .S2(n2570), .D3(n2528), .S3(n2572), .Z(n2973) );
  HS65_LHS_XOR2X3 U2740 ( .A(n2641), .B(n2974), .Z(n1168) );
  HS65_LH_MX41X4 U2741 ( .D0(n2966), .S0(n1033), .D1(n2524), .S1(n2576), .D2(
        n2532), .S2(n2572), .D3(n2528), .S3(n2574), .Z(n2974) );
  HS65_LHS_XOR2X3 U2742 ( .A(n91), .B(n2975), .Z(n1167) );
  HS65_LH_MX41X4 U2743 ( .D0(n2966), .S0(n1032), .D1(n2524), .S1(n2578), .D2(
        n2532), .S2(n2574), .D3(n2528), .S3(n2576), .Z(n2975) );
  HS65_LHS_XOR2X3 U2744 ( .A(n2641), .B(n2976), .Z(n1166) );
  HS65_LH_MX41X4 U2745 ( .D0(n2526), .S0(n1031), .D1(n2524), .S1(n2580), .D2(
        n2532), .S2(n2576), .D3(n2528), .S3(n2578), .Z(n2976) );
  HS65_LHS_XOR2X3 U2746 ( .A(n2641), .B(n2977), .Z(n1165) );
  HS65_LH_MX41X4 U2747 ( .D0(n2966), .S0(n1030), .D1(n2524), .S1(n2582), .D2(
        n2532), .S2(n2578), .D3(n2529), .S3(n2580), .Z(n2977) );
  HS65_LHS_XOR2X3 U2748 ( .A(n2641), .B(n2978), .Z(n1164) );
  HS65_LH_MX41X4 U2749 ( .D0(n2966), .S0(n1029), .D1(n2524), .S1(n2584), .D2(
        n2532), .S2(n2580), .D3(n2528), .S3(n2582), .Z(n2978) );
  HS65_LHS_XOR2X3 U2750 ( .A(n2641), .B(n2979), .Z(n1163) );
  HS65_LH_MX41X4 U2751 ( .D0(n2966), .S0(n1028), .D1(n2524), .S1(n2586), .D2(
        n2532), .S2(n2582), .D3(n2528), .S3(n2584), .Z(n2979) );
  HS65_LHS_XOR2X3 U2752 ( .A(n91), .B(n2980), .Z(n1162) );
  HS65_LH_MX41X4 U2753 ( .D0(n2966), .S0(n1027), .D1(n2524), .S1(n2588), .D2(
        n2532), .S2(n2584), .D3(n2528), .S3(n2586), .Z(n2980) );
  HS65_LHS_XOR2X3 U2754 ( .A(n91), .B(n2981), .Z(n1161) );
  HS65_LH_MX41X4 U2755 ( .D0(n2966), .S0(n1026), .D1(n2524), .S1(n2590), .D2(
        n2532), .S2(n2586), .D3(n2529), .S3(n2588), .Z(n2981) );
  HS65_LHS_XOR2X3 U2756 ( .A(n91), .B(n2982), .Z(n1160) );
  HS65_LH_MX41X4 U2757 ( .D0(n2966), .S0(n1025), .D1(n2524), .S1(n2592), .D2(
        n2532), .S2(n2588), .D3(n2529), .S3(n2590), .Z(n2982) );
  HS65_LHS_XOR2X3 U2758 ( .A(n91), .B(n2983), .Z(n1159) );
  HS65_LH_MX41X4 U2759 ( .D0(n2966), .S0(n1024), .D1(n2524), .S1(n2594), .D2(
        n2533), .S2(n2590), .D3(n2529), .S3(n2592), .Z(n2983) );
  HS65_LHS_XOR2X3 U2760 ( .A(n2641), .B(n2984), .Z(n1158) );
  HS65_LH_MX41X4 U2761 ( .D0(n2526), .S0(n1023), .D1(n2525), .S1(n2596), .D2(
        n2533), .S2(n2592), .D3(n2529), .S3(n2594), .Z(n2984) );
  HS65_LHS_XOR2X3 U2762 ( .A(n2641), .B(n2985), .Z(n1157) );
  HS65_LH_MX41X4 U2763 ( .D0(n2526), .S0(n1022), .D1(n2525), .S1(n2598), .D2(
        n2533), .S2(n2594), .D3(n2529), .S3(n2596), .Z(n2985) );
  HS65_LHS_XOR2X3 U2764 ( .A(n91), .B(n2986), .Z(n1156) );
  HS65_LH_MX41X4 U2765 ( .D0(n2526), .S0(n1021), .D1(n2525), .S1(n2600), .D2(
        n2533), .S2(n2596), .D3(n2529), .S3(n2598), .Z(n2986) );
  HS65_LHS_XOR2X3 U2766 ( .A(n2641), .B(n2987), .Z(n1155) );
  HS65_LH_MX41X4 U2767 ( .D0(n2526), .S0(n1020), .D1(n2525), .S1(n2602), .D2(
        n2533), .S2(n2598), .D3(n2529), .S3(n2600), .Z(n2987) );
  HS65_LHS_XOR2X3 U2768 ( .A(n91), .B(n2988), .Z(n1154) );
  HS65_LH_MX41X4 U2769 ( .D0(n2526), .S0(n1019), .D1(n2525), .S1(n2604), .D2(
        n2533), .S2(n2600), .D3(n2529), .S3(n2602), .Z(n2988) );
  HS65_LHS_XOR2X3 U2770 ( .A(n2641), .B(n2989), .Z(n1153) );
  HS65_LH_MX41X4 U2771 ( .D0(n2526), .S0(n1018), .D1(n2525), .S1(n2606), .D2(
        n2533), .S2(n2602), .D3(n2529), .S3(n2604), .Z(n2989) );
  HS65_LHS_XOR2X3 U2772 ( .A(n91), .B(n2990), .Z(n1152) );
  HS65_LH_MX41X4 U2773 ( .D0(n2526), .S0(n1017), .D1(n2525), .S1(n2608), .D2(
        n2533), .S2(n2604), .D3(n2529), .S3(n2606), .Z(n2990) );
  HS65_LHS_XOR2X3 U2774 ( .A(n91), .B(n2991), .Z(n1151) );
  HS65_LH_MX41X4 U2775 ( .D0(n2526), .S0(n1016), .D1(n2525), .S1(n2610), .D2(
        n2533), .S2(n2606), .D3(n2529), .S3(n2608), .Z(n2991) );
  HS65_LHS_XOR2X3 U2776 ( .A(n2641), .B(n2992), .Z(n1150) );
  HS65_LH_MX41X4 U2777 ( .D0(n2526), .S0(n1015), .D1(n2525), .S1(n2612), .D2(
        n2533), .S2(n2608), .D3(n2529), .S3(n2610), .Z(n2992) );
  HS65_LHS_XOR2X3 U2778 ( .A(n2641), .B(n2993), .Z(n1149) );
  HS65_LH_MX41X4 U2779 ( .D0(n2526), .S0(n1014), .D1(n2525), .S1(n2614), .D2(
        n2533), .S2(n2610), .D3(n2529), .S3(n2612), .Z(n2993) );
  HS65_LHS_XOR2X3 U2780 ( .A(n91), .B(n2994), .Z(n1148) );
  HS65_LH_MX41X4 U2781 ( .D0(n2526), .S0(n1013), .D1(n2525), .S1(n2616), .D2(
        n2533), .S2(n2612), .D3(n2530), .S3(n2614), .Z(n2994) );
  HS65_LHS_XOR2X3 U2782 ( .A(n91), .B(n2995), .Z(n1147) );
  HS65_LH_MX41X4 U2783 ( .D0(n2526), .S0(n1012), .D1(n2525), .S1(n2618), .D2(
        n2533), .S2(n2614), .D3(n2530), .S3(n2616), .Z(n2995) );
  HS65_LHS_XOR2X3 U2784 ( .A(n2641), .B(n2996), .Z(n1146) );
  HS65_LH_MX41X4 U2785 ( .D0(n2526), .S0(n1011), .D1(n2525), .S1(n2620), .D2(
        n2534), .S2(n2616), .D3(n2530), .S3(n2618), .Z(n2996) );
  HS65_LHS_XOR2X3 U2786 ( .A(n91), .B(n2997), .Z(n1145) );
  HS65_LH_MX41X4 U2787 ( .D0(n2526), .S0(n1010), .D1(n2525), .S1(n2622), .D2(
        n2534), .S2(n2618), .D3(n2530), .S3(n2620), .Z(n2997) );
  HS65_LHS_XOR2X3 U2788 ( .A(n91), .B(n2998), .Z(n1144) );
  HS65_LH_MX41X4 U2789 ( .D0(n2966), .S0(n1009), .D1(n2525), .S1(n2624), .D2(
        n2534), .S2(n2620), .D3(n2530), .S3(n2622), .Z(n2998) );
  HS65_LHS_XOR2X3 U2790 ( .A(n91), .B(n2999), .Z(n1143) );
  HS65_LH_MX41X4 U2791 ( .D0(n2966), .S0(n1008), .D1(n2525), .S1(n2626), .D2(
        n2534), .S2(n2622), .D3(n2528), .S3(n2624), .Z(n2999) );
  HS65_LH_AND2X4 U2792 ( .A(n3000), .B(n3001), .Z(n2965) );
  HS65_LHS_XOR2X3 U2793 ( .A(n91), .B(n3002), .Z(n1142) );
  HS65_LH_OAI12X2 U2794 ( .A(n2657), .B(n2527), .C(n3003), .Z(n3002) );
  HS65_LH_OAI22X1 U2795 ( .A(n2625), .B(n3004), .C(n2532), .D(n3004), .Z(n3003) );
  HS65_LH_AND2X4 U2796 ( .A(n2528), .B(n2626), .Z(n3004) );
  HS65_LH_NOR2X2 U2797 ( .A(n3000), .B(n3005), .Z(n2968) );
  HS65_LHS_XOR2X3 U2798 ( .A(n2642), .B(n3006), .Z(n1141) );
  HS65_LH_AOI22X1 U2799 ( .A(n2966), .B(n1006), .C(n2534), .D(n2627), .Z(n3006) );
  HS65_LH_NOR3AX2 U2800 ( .A(n3005), .B(n3001), .C(n3000), .Z(n2970) );
  HS65_LHS_XNOR2X3 U2801 ( .A(a[22]), .B(a[21]), .Z(n3005) );
  HS65_LH_NOR2AX3 U2802 ( .A(n3000), .B(n3001), .Z(n2966) );
  HS65_LHS_XNOR2X3 U2803 ( .A(n2641), .B(a[22]), .Z(n3001) );
  HS65_LHS_XOR2X3 U2804 ( .A(n2639), .B(a[21]), .Z(n3000) );
  HS65_LHS_XOR2X3 U2805 ( .A(n2643), .B(n3007), .Z(n1139) );
  HS65_LH_AO22X4 U2806 ( .A(n2565), .B(n2537), .C(n2564), .D(n3009), .Z(n3007)
         );
  HS65_LHS_XOR2X3 U2807 ( .A(n2643), .B(n3010), .Z(n1138) );
  HS65_LH_AO222X4 U2808 ( .A(n2567), .B(n2537), .C(n2563), .D(n2541), .E(n1038), .F(n3009), .Z(n3010) );
  HS65_LHS_XOR2X3 U2809 ( .A(n2643), .B(n3012), .Z(n1137) );
  HS65_LH_MX41X4 U2810 ( .D0(n3009), .S0(n1037), .D1(n2546), .S1(n2563), .D2(
        n2541), .S2(n2566), .D3(n2537), .S3(n2568), .Z(n3012) );
  HS65_LHS_XOR2X3 U2811 ( .A(n2643), .B(n3014), .Z(n1136) );
  HS65_LH_MX41X4 U2812 ( .D0(n2539), .S0(n1036), .D1(n2545), .S1(n2567), .D2(
        n2541), .S2(n2568), .D3(n2537), .S3(n2570), .Z(n3014) );
  HS65_LHS_XOR2X3 U2813 ( .A(n2643), .B(n3015), .Z(n1135) );
  HS65_LH_MX41X4 U2814 ( .D0(n3009), .S0(n1035), .D1(n2545), .S1(n2568), .D2(
        n2541), .S2(n2570), .D3(n2537), .S3(n2572), .Z(n3015) );
  HS65_LHS_XOR2X3 U2815 ( .A(n2643), .B(n3016), .Z(n1134) );
  HS65_LH_MX41X4 U2816 ( .D0(n2539), .S0(n1034), .D1(n2545), .S1(n2570), .D2(
        n2541), .S2(n2572), .D3(n2537), .S3(n2574), .Z(n3016) );
  HS65_LHS_XOR2X3 U2817 ( .A(n2643), .B(n3017), .Z(n1133) );
  HS65_LH_MX41X4 U2818 ( .D0(n3009), .S0(n1033), .D1(n2545), .S1(n2572), .D2(
        n2541), .S2(n2574), .D3(n2537), .S3(n2576), .Z(n3017) );
  HS65_LHS_XOR2X3 U2819 ( .A(n103), .B(n3018), .Z(n1132) );
  HS65_LH_MX41X4 U2820 ( .D0(n3009), .S0(n1032), .D1(n2545), .S1(n2574), .D2(
        n2541), .S2(n2576), .D3(n2537), .S3(n2578), .Z(n3018) );
  HS65_LHS_XOR2X3 U2821 ( .A(n2643), .B(n3019), .Z(n1131) );
  HS65_LH_MX41X4 U2822 ( .D0(n2539), .S0(n1031), .D1(n2545), .S1(n2576), .D2(
        n2541), .S2(n2578), .D3(n2537), .S3(n2580), .Z(n3019) );
  HS65_LHS_XOR2X3 U2823 ( .A(n2643), .B(n3020), .Z(n1130) );
  HS65_LH_MX41X4 U2824 ( .D0(n3009), .S0(n1030), .D1(n2545), .S1(n2578), .D2(
        n2542), .S2(n2580), .D3(n2537), .S3(n2582), .Z(n3020) );
  HS65_LHS_XOR2X3 U2825 ( .A(n2643), .B(n3021), .Z(n1129) );
  HS65_LH_MX41X4 U2826 ( .D0(n3009), .S0(n1029), .D1(n2545), .S1(n2580), .D2(
        n2541), .S2(n2582), .D3(n2537), .S3(n2584), .Z(n3021) );
  HS65_LHS_XOR2X3 U2827 ( .A(n2643), .B(n3022), .Z(n1128) );
  HS65_LH_MX41X4 U2828 ( .D0(n3009), .S0(n1028), .D1(n2545), .S1(n2582), .D2(
        n2541), .S2(n2584), .D3(n2537), .S3(n2586), .Z(n3022) );
  HS65_LHS_XOR2X3 U2829 ( .A(n103), .B(n3023), .Z(n1127) );
  HS65_LH_MX41X4 U2830 ( .D0(n3009), .S0(n1027), .D1(n2545), .S1(n2584), .D2(
        n2541), .S2(n2586), .D3(n2537), .S3(n2588), .Z(n3023) );
  HS65_LHS_XOR2X3 U2831 ( .A(n103), .B(n3024), .Z(n1126) );
  HS65_LH_MX41X4 U2832 ( .D0(n3009), .S0(n1026), .D1(n2545), .S1(n2586), .D2(
        n2542), .S2(n2588), .D3(n2537), .S3(n2590), .Z(n3024) );
  HS65_LHS_XOR2X3 U2833 ( .A(n103), .B(n3025), .Z(n1125) );
  HS65_LH_MX41X4 U2834 ( .D0(n3009), .S0(n1025), .D1(n2545), .S1(n2588), .D2(
        n2542), .S2(n2590), .D3(n2537), .S3(n2592), .Z(n3025) );
  HS65_LHS_XOR2X3 U2835 ( .A(n103), .B(n3026), .Z(n1124) );
  HS65_LH_MX41X4 U2836 ( .D0(n3009), .S0(n1024), .D1(n2546), .S1(n2590), .D2(
        n2542), .S2(n2592), .D3(n2537), .S3(n2594), .Z(n3026) );
  HS65_LHS_XOR2X3 U2837 ( .A(n2643), .B(n3027), .Z(n1123) );
  HS65_LH_MX41X4 U2838 ( .D0(n2539), .S0(n1023), .D1(n2546), .S1(n2592), .D2(
        n2542), .S2(n2594), .D3(n2537), .S3(n2596), .Z(n3027) );
  HS65_LHS_XOR2X3 U2839 ( .A(n2643), .B(n3028), .Z(n1122) );
  HS65_LH_MX41X4 U2840 ( .D0(n2539), .S0(n1022), .D1(n2546), .S1(n2594), .D2(
        n2542), .S2(n2596), .D3(n2538), .S3(n2598), .Z(n3028) );
  HS65_LHS_XOR2X3 U2841 ( .A(n103), .B(n3029), .Z(n1121) );
  HS65_LH_MX41X4 U2842 ( .D0(n2539), .S0(n1021), .D1(n2546), .S1(n2596), .D2(
        n2542), .S2(n2598), .D3(n2538), .S3(n2600), .Z(n3029) );
  HS65_LHS_XOR2X3 U2843 ( .A(n2643), .B(n3030), .Z(n1120) );
  HS65_LH_MX41X4 U2844 ( .D0(n2539), .S0(n1020), .D1(n2546), .S1(n2598), .D2(
        n2542), .S2(n2600), .D3(n2538), .S3(n2602), .Z(n3030) );
  HS65_LHS_XOR2X3 U2845 ( .A(n103), .B(n3031), .Z(n1119) );
  HS65_LH_MX41X4 U2846 ( .D0(n2539), .S0(n1019), .D1(n2546), .S1(n2600), .D2(
        n2542), .S2(n2602), .D3(n2538), .S3(n2604), .Z(n3031) );
  HS65_LHS_XOR2X3 U2847 ( .A(n2643), .B(n3032), .Z(n1118) );
  HS65_LH_MX41X4 U2848 ( .D0(n2539), .S0(n1018), .D1(n2546), .S1(n2602), .D2(
        n2542), .S2(n2604), .D3(n2538), .S3(n2606), .Z(n3032) );
  HS65_LHS_XOR2X3 U2849 ( .A(n103), .B(n3033), .Z(n1117) );
  HS65_LH_MX41X4 U2850 ( .D0(n2539), .S0(n1017), .D1(n2546), .S1(n2604), .D2(
        n2542), .S2(n2606), .D3(n2538), .S3(n2608), .Z(n3033) );
  HS65_LHS_XOR2X3 U2851 ( .A(n103), .B(n3034), .Z(n1116) );
  HS65_LH_MX41X4 U2852 ( .D0(n2539), .S0(n1016), .D1(n2546), .S1(n2606), .D2(
        n2542), .S2(n2608), .D3(n2538), .S3(n2610), .Z(n3034) );
  HS65_LHS_XOR2X3 U2853 ( .A(n2643), .B(n3035), .Z(n1115) );
  HS65_LH_MX41X4 U2854 ( .D0(n2539), .S0(n1015), .D1(n2546), .S1(n2608), .D2(
        n2542), .S2(n2610), .D3(n2538), .S3(n2612), .Z(n3035) );
  HS65_LHS_XOR2X3 U2855 ( .A(n2643), .B(n3036), .Z(n1114) );
  HS65_LH_MX41X4 U2856 ( .D0(n2539), .S0(n1014), .D1(n2546), .S1(n2610), .D2(
        n2542), .S2(n2612), .D3(n2538), .S3(n2614), .Z(n3036) );
  HS65_LHS_XOR2X3 U2857 ( .A(n103), .B(n3037), .Z(n1113) );
  HS65_LH_MX41X4 U2858 ( .D0(n2539), .S0(n1013), .D1(n2546), .S1(n2612), .D2(
        n2543), .S2(n2614), .D3(n2538), .S3(n2616), .Z(n3037) );
  HS65_LHS_XOR2X3 U2859 ( .A(n103), .B(n3038), .Z(n1112) );
  HS65_LH_MX41X4 U2860 ( .D0(n2539), .S0(n1012), .D1(n2547), .S1(n2614), .D2(
        n2543), .S2(n2616), .D3(n2538), .S3(n2618), .Z(n3038) );
  HS65_LHS_XOR2X3 U2861 ( .A(n2643), .B(n3039), .Z(n1111) );
  HS65_LH_MX41X4 U2862 ( .D0(n2539), .S0(n1011), .D1(n2547), .S1(n2616), .D2(
        n2543), .S2(n2618), .D3(n2538), .S3(n2620), .Z(n3039) );
  HS65_LHS_XOR2X3 U2863 ( .A(n103), .B(n3040), .Z(n1110) );
  HS65_LH_MX41X4 U2864 ( .D0(n2539), .S0(n1010), .D1(n2547), .S1(n2618), .D2(
        n2543), .S2(n2620), .D3(n2538), .S3(n2622), .Z(n3040) );
  HS65_LHS_XOR2X3 U2865 ( .A(n103), .B(n3041), .Z(n1109) );
  HS65_LH_MX41X4 U2866 ( .D0(n3009), .S0(n1009), .D1(n2547), .S1(n2620), .D2(
        n2543), .S2(n2622), .D3(n2538), .S3(n2624), .Z(n3041) );
  HS65_LHS_XOR2X3 U2867 ( .A(n103), .B(n3042), .Z(n1108) );
  HS65_LH_MX41X4 U2868 ( .D0(n3009), .S0(n1008), .D1(n2547), .S1(n2622), .D2(
        n2541), .S2(n2624), .D3(n2538), .S3(n2626), .Z(n3042) );
  HS65_LH_AND2X4 U2869 ( .A(n3043), .B(n3044), .Z(n3008) );
  HS65_LHS_XOR2X3 U2870 ( .A(n103), .B(n3045), .Z(n1107) );
  HS65_LH_OAI12X2 U2871 ( .A(n2657), .B(n2540), .C(n3046), .Z(n3045) );
  HS65_LH_OAI22X1 U2872 ( .A(n2625), .B(n3047), .C(n2545), .D(n3047), .Z(n3046) );
  HS65_LH_AND2X4 U2873 ( .A(n2541), .B(n2626), .Z(n3047) );
  HS65_LH_NOR2X2 U2874 ( .A(n3043), .B(n3048), .Z(n3011) );
  HS65_LHS_XOR2X3 U2875 ( .A(n2644), .B(n3049), .Z(n1106) );
  HS65_LH_AOI22X1 U2876 ( .A(n3009), .B(n1006), .C(n2547), .D(n2627), .Z(n3049) );
  HS65_LH_NOR3AX2 U2877 ( .A(n3048), .B(n3044), .C(n3043), .Z(n3013) );
  HS65_LHS_XNOR2X3 U2878 ( .A(a[25]), .B(a[24]), .Z(n3048) );
  HS65_LH_NOR2AX3 U2879 ( .A(n3043), .B(n3044), .Z(n3009) );
  HS65_LHS_XNOR2X3 U2880 ( .A(n2643), .B(a[25]), .Z(n3044) );
  HS65_LHS_XOR2X3 U2881 ( .A(n2641), .B(a[24]), .Z(n3043) );
  HS65_LHS_XOR2X3 U2882 ( .A(n2645), .B(n3050), .Z(n1104) );
  HS65_LH_AO22X4 U2883 ( .A(n2565), .B(n2550), .C(n2564), .D(n3052), .Z(n3050)
         );
  HS65_LHS_XOR2X3 U2884 ( .A(n2645), .B(n3053), .Z(n1103) );
  HS65_LH_AO222X4 U2885 ( .A(n2567), .B(n2550), .C(n2563), .D(n2554), .E(n1038), .F(n3052), .Z(n3053) );
  HS65_LHS_XOR2X3 U2886 ( .A(n2645), .B(n3055), .Z(n1102) );
  HS65_LH_MX41X4 U2887 ( .D0(n3052), .S0(n1037), .D1(n2559), .S1(n2563), .D2(
        n2554), .S2(n2566), .D3(n2550), .S3(n2568), .Z(n3055) );
  HS65_LHS_XOR2X3 U2888 ( .A(n2645), .B(n3057), .Z(n1101) );
  HS65_LH_MX41X4 U2889 ( .D0(n2552), .S0(n1036), .D1(n2558), .S1(n2567), .D2(
        n2554), .S2(n2568), .D3(n2550), .S3(n2570), .Z(n3057) );
  HS65_LHS_XOR2X3 U2890 ( .A(n2645), .B(n3058), .Z(n1100) );
  HS65_LH_MX41X4 U2891 ( .D0(n3052), .S0(n1035), .D1(n2558), .S1(n2568), .D2(
        n2554), .S2(n2570), .D3(n2550), .S3(n2572), .Z(n3058) );
  HS65_LHS_XOR2X3 U2892 ( .A(n2645), .B(n3059), .Z(n1099) );
  HS65_LH_MX41X4 U2893 ( .D0(n2552), .S0(n1034), .D1(n2558), .S1(n2570), .D2(
        n2554), .S2(n2572), .D3(n2550), .S3(n2574), .Z(n3059) );
  HS65_LHS_XOR2X3 U2894 ( .A(n2645), .B(n3060), .Z(n1098) );
  HS65_LH_MX41X4 U2895 ( .D0(n3052), .S0(n1033), .D1(n2558), .S1(n2572), .D2(
        n2554), .S2(n2574), .D3(n2550), .S3(n2576), .Z(n3060) );
  HS65_LHS_XOR2X3 U2896 ( .A(n115), .B(n3061), .Z(n1097) );
  HS65_LH_MX41X4 U2897 ( .D0(n3052), .S0(n1032), .D1(n2558), .S1(n2574), .D2(
        n2554), .S2(n2576), .D3(n2550), .S3(n2578), .Z(n3061) );
  HS65_LHS_XOR2X3 U2898 ( .A(n2645), .B(n3062), .Z(n1096) );
  HS65_LH_MX41X4 U2899 ( .D0(n2552), .S0(n1031), .D1(n2558), .S1(n2576), .D2(
        n2554), .S2(n2578), .D3(n2550), .S3(n2580), .Z(n3062) );
  HS65_LHS_XOR2X3 U2900 ( .A(n2645), .B(n3063), .Z(n1095) );
  HS65_LH_MX41X4 U2901 ( .D0(n3052), .S0(n1030), .D1(n2558), .S1(n2578), .D2(
        n2555), .S2(n2580), .D3(n2550), .S3(n2582), .Z(n3063) );
  HS65_LHS_XOR2X3 U2902 ( .A(n2645), .B(n3064), .Z(n1094) );
  HS65_LH_MX41X4 U2903 ( .D0(n3052), .S0(n1029), .D1(n2558), .S1(n2580), .D2(
        n2554), .S2(n2582), .D3(n2550), .S3(n2584), .Z(n3064) );
  HS65_LHS_XOR2X3 U2904 ( .A(n2645), .B(n3065), .Z(n1093) );
  HS65_LH_MX41X4 U2905 ( .D0(n3052), .S0(n1028), .D1(n2558), .S1(n2582), .D2(
        n2554), .S2(n2584), .D3(n2550), .S3(n2586), .Z(n3065) );
  HS65_LHS_XOR2X3 U2906 ( .A(n115), .B(n3066), .Z(n1092) );
  HS65_LH_MX41X4 U2907 ( .D0(n3052), .S0(n1027), .D1(n2558), .S1(n2584), .D2(
        n2554), .S2(n2586), .D3(n2550), .S3(n2588), .Z(n3066) );
  HS65_LHS_XOR2X3 U2908 ( .A(n115), .B(n3067), .Z(n1091) );
  HS65_LH_MX41X4 U2909 ( .D0(n3052), .S0(n1026), .D1(n2558), .S1(n2586), .D2(
        n2555), .S2(n2588), .D3(n2550), .S3(n2590), .Z(n3067) );
  HS65_LHS_XOR2X3 U2910 ( .A(n115), .B(n3068), .Z(n1090) );
  HS65_LH_MX41X4 U2911 ( .D0(n3052), .S0(n1025), .D1(n2558), .S1(n2588), .D2(
        n2555), .S2(n2590), .D3(n2550), .S3(n2592), .Z(n3068) );
  HS65_LHS_XOR2X3 U2912 ( .A(n115), .B(n3069), .Z(n1089) );
  HS65_LH_MX41X4 U2913 ( .D0(n3052), .S0(n1024), .D1(n2559), .S1(n2590), .D2(
        n2555), .S2(n2592), .D3(n2550), .S3(n2594), .Z(n3069) );
  HS65_LHS_XOR2X3 U2914 ( .A(n2645), .B(n3070), .Z(n1088) );
  HS65_LH_MX41X4 U2915 ( .D0(n2552), .S0(n1023), .D1(n2559), .S1(n2592), .D2(
        n2555), .S2(n2594), .D3(n2550), .S3(n2596), .Z(n3070) );
  HS65_LHS_XOR2X3 U2916 ( .A(n2645), .B(n3071), .Z(n1087) );
  HS65_LH_MX41X4 U2917 ( .D0(n2552), .S0(n1022), .D1(n2559), .S1(n2594), .D2(
        n2555), .S2(n2596), .D3(n2551), .S3(n2598), .Z(n3071) );
  HS65_LHS_XOR2X3 U2918 ( .A(n115), .B(n3072), .Z(n1086) );
  HS65_LH_MX41X4 U2919 ( .D0(n2552), .S0(n1021), .D1(n2559), .S1(n2596), .D2(
        n2555), .S2(n2598), .D3(n2551), .S3(n2600), .Z(n3072) );
  HS65_LHS_XOR2X3 U2920 ( .A(n2645), .B(n3073), .Z(n1085) );
  HS65_LH_MX41X4 U2921 ( .D0(n2552), .S0(n1020), .D1(n2559), .S1(n2598), .D2(
        n2555), .S2(n2600), .D3(n2551), .S3(n2602), .Z(n3073) );
  HS65_LHS_XOR2X3 U2922 ( .A(n115), .B(n3074), .Z(n1084) );
  HS65_LH_MX41X4 U2923 ( .D0(n2552), .S0(n1019), .D1(n2559), .S1(n2600), .D2(
        n2555), .S2(n2602), .D3(n2551), .S3(n2604), .Z(n3074) );
  HS65_LHS_XOR2X3 U2924 ( .A(n2645), .B(n3075), .Z(n1083) );
  HS65_LH_MX41X4 U2925 ( .D0(n2552), .S0(n1018), .D1(n2559), .S1(n2602), .D2(
        n2555), .S2(n2604), .D3(n2551), .S3(n2606), .Z(n3075) );
  HS65_LHS_XOR2X3 U2926 ( .A(n115), .B(n3076), .Z(n1082) );
  HS65_LH_MX41X4 U2927 ( .D0(n2552), .S0(n1017), .D1(n2559), .S1(n2604), .D2(
        n2555), .S2(n2606), .D3(n2551), .S3(n2608), .Z(n3076) );
  HS65_LHS_XOR2X3 U2928 ( .A(n2645), .B(n3077), .Z(n1081) );
  HS65_LH_MX41X4 U2929 ( .D0(n2552), .S0(n1016), .D1(n2559), .S1(n2606), .D2(
        n2555), .S2(n2608), .D3(n2551), .S3(n2610), .Z(n3077) );
  HS65_LHS_XOR2X3 U2930 ( .A(n2645), .B(n3078), .Z(n1080) );
  HS65_LH_MX41X4 U2931 ( .D0(n2552), .S0(n1015), .D1(n2559), .S1(n2608), .D2(
        n2555), .S2(n2610), .D3(n2551), .S3(n2612), .Z(n3078) );
  HS65_LHS_XOR2X3 U2932 ( .A(n115), .B(n3079), .Z(n1079) );
  HS65_LH_MX41X4 U2933 ( .D0(n2552), .S0(n1014), .D1(n2559), .S1(n2610), .D2(
        n2555), .S2(n2612), .D3(n2551), .S3(n2614), .Z(n3079) );
  HS65_LHS_XOR2X3 U2934 ( .A(n115), .B(n3080), .Z(n1078) );
  HS65_LH_MX41X4 U2935 ( .D0(n2552), .S0(n1013), .D1(n2559), .S1(n2612), .D2(
        n2556), .S2(n2614), .D3(n2551), .S3(n2616), .Z(n3080) );
  HS65_LHS_XOR2X3 U2936 ( .A(n2645), .B(n3081), .Z(n1077) );
  HS65_LH_MX41X4 U2937 ( .D0(n2552), .S0(n1012), .D1(n2560), .S1(n2614), .D2(
        n2556), .S2(n2616), .D3(n2551), .S3(n2618), .Z(n3081) );
  HS65_LHS_XOR2X3 U2938 ( .A(n115), .B(n3082), .Z(n1076) );
  HS65_LH_MX41X4 U2939 ( .D0(n2552), .S0(n1011), .D1(n2560), .S1(n2616), .D2(
        n2556), .S2(n2618), .D3(n2551), .S3(n2620), .Z(n3082) );
  HS65_LHS_XOR2X3 U2940 ( .A(n115), .B(n3083), .Z(n1075) );
  HS65_LH_MX41X4 U2941 ( .D0(n2552), .S0(n1010), .D1(n2560), .S1(n2618), .D2(
        n2556), .S2(n2620), .D3(n2551), .S3(n2622), .Z(n3083) );
  HS65_LHS_XOR2X3 U2942 ( .A(n115), .B(n3084), .Z(n1074) );
  HS65_LH_MX41X4 U2943 ( .D0(n3052), .S0(n1009), .D1(n2560), .S1(n2620), .D2(
        n2556), .S2(n2622), .D3(n2551), .S3(n2624), .Z(n3084) );
  HS65_LHS_XOR2X3 U2944 ( .A(n115), .B(n3085), .Z(n1073) );
  HS65_LH_MX41X4 U2945 ( .D0(n3052), .S0(n1008), .D1(n2560), .S1(n2622), .D2(
        n2554), .S2(n2624), .D3(n2551), .S3(n2626), .Z(n3085) );
  HS65_LH_AND2X4 U2946 ( .A(n3086), .B(n3087), .Z(n3051) );
  HS65_LHS_XOR2X3 U2947 ( .A(n115), .B(n3088), .Z(n1072) );
  HS65_LH_OAI12X2 U2948 ( .A(n2657), .B(n2553), .C(n3089), .Z(n3088) );
  HS65_LH_OAI22X1 U2949 ( .A(n2625), .B(n3090), .C(n2558), .D(n3090), .Z(n3089) );
  HS65_LH_AND2X4 U2950 ( .A(n2554), .B(n2626), .Z(n3090) );
  HS65_LH_NOR2X2 U2951 ( .A(n3086), .B(n3091), .Z(n3054) );
  HS65_LHS_XOR2X3 U2952 ( .A(n2646), .B(n3092), .Z(n1071) );
  HS65_LH_AOI22X1 U2953 ( .A(n3052), .B(n1006), .C(n2560), .D(n2627), .Z(n3092) );
  HS65_LH_NOR3AX2 U2954 ( .A(n3091), .B(n3087), .C(n3086), .Z(n3056) );
  HS65_LHS_XNOR2X3 U2955 ( .A(a[28]), .B(a[27]), .Z(n3091) );
  HS65_LH_NOR2AX3 U2956 ( .A(n3086), .B(n3087), .Z(n3052) );
  HS65_LHS_XNOR2X3 U2957 ( .A(n115), .B(a[28]), .Z(n3087) );
  HS65_LHS_XOR2X3 U2958 ( .A(n2643), .B(a[27]), .Z(n3086) );
  HS65_LH_AO22X4 U2959 ( .A(n2428), .B(n2563), .C(n2419), .D(n2564), .Z(n1069)
         );
  HS65_LH_AO222X4 U2960 ( .A(n2428), .B(n2566), .C(n2432), .D(n2563), .E(n2419), .F(n1038), .Z(n1068) );
  HS65_LH_MX41X4 U2961 ( .D0(n1037), .S0(n2419), .D1(n2569), .S1(n2426), .D2(
        n2567), .S2(n2430), .D3(n2564), .S3(n2423), .Z(n1067) );
  HS65_LH_MX41X4 U2962 ( .D0(n1036), .S0(n2419), .D1(n2571), .S1(n2426), .D2(
        n2569), .S2(n2430), .D3(n2567), .S3(n2423), .Z(n1066) );
  HS65_LH_MX41X4 U2963 ( .D0(n1035), .S0(n2419), .D1(n2573), .S1(n2426), .D2(
        n2571), .S2(n2430), .D3(n2569), .S3(n2423), .Z(n1065) );
  HS65_LH_MX41X4 U2964 ( .D0(n1034), .S0(n2418), .D1(n2575), .S1(n2426), .D2(
        n2573), .S2(n2430), .D3(n2571), .S3(n2423), .Z(n1064) );
  HS65_LH_MX41X4 U2965 ( .D0(n1033), .S0(n2418), .D1(n2577), .S1(n2426), .D2(
        n2575), .S2(n2430), .D3(n2573), .S3(n2423), .Z(n1063) );
  HS65_LH_MX41X4 U2966 ( .D0(n1032), .S0(n2418), .D1(n2579), .S1(n2426), .D2(
        n2577), .S2(n2430), .D3(n2575), .S3(n2423), .Z(n1062) );
  HS65_LH_MX41X4 U2967 ( .D0(n1031), .S0(n2418), .D1(n2581), .S1(n2426), .D2(
        n2579), .S2(n2430), .D3(n2577), .S3(n2423), .Z(n1061) );
  HS65_LH_MX41X4 U2968 ( .D0(n1030), .S0(n2418), .D1(n2583), .S1(n2426), .D2(
        n2581), .S2(n2430), .D3(n2579), .S3(n2423), .Z(n1060) );
  HS65_LH_MX41X4 U2969 ( .D0(n1029), .S0(n2418), .D1(n2585), .S1(n2426), .D2(
        n2583), .S2(n2430), .D3(n2581), .S3(n2423), .Z(n1059) );
  HS65_LH_MX41X4 U2970 ( .D0(n1028), .S0(n2418), .D1(n2587), .S1(n2426), .D2(
        n2585), .S2(n2431), .D3(n2583), .S3(n2424), .Z(n1058) );
  HS65_LH_MX41X4 U2971 ( .D0(n1027), .S0(n2418), .D1(n2428), .S1(n2588), .D2(
        n2587), .S2(n2431), .D3(n2585), .S3(n2424), .Z(n1057) );
  HS65_LH_MX41X4 U2972 ( .D0(n1026), .S0(n2418), .D1(n2428), .S1(n2590), .D2(
        n2589), .S2(n2431), .D3(n2587), .S3(n2424), .Z(n1056) );
  HS65_LH_MX41X4 U2973 ( .D0(n1024), .S0(n2418), .D1(n2593), .S1(n2432), .D2(
        n2591), .S2(n2423), .D3(n2595), .S3(n2426), .Z(n1055) );
  HS65_LH_MX41X4 U2974 ( .D0(n1023), .S0(n2418), .D1(n2593), .S1(n2424), .D2(
        n2595), .S2(n2431), .D3(n2597), .S3(n2427), .Z(n1054) );
  HS65_LH_MX41X4 U2975 ( .D0(n1022), .S0(n2417), .D1(n2595), .S1(n2424), .D2(
        n2597), .S2(n2431), .D3(n2599), .S3(n2427), .Z(n1053) );
  HS65_LH_MX41X4 U2976 ( .D0(n1021), .S0(n2417), .D1(n2597), .S1(n2424), .D2(
        n2599), .S2(n2431), .D3(n2601), .S3(n2427), .Z(n1052) );
  HS65_LH_MX41X4 U2977 ( .D0(n1020), .S0(n2417), .D1(n2599), .S1(n2424), .D2(
        n2601), .S2(n2431), .D3(n2603), .S3(n2427), .Z(n1051) );
  HS65_LH_MX41X4 U2978 ( .D0(n1018), .S0(n2417), .D1(n2603), .S1(n2424), .D2(
        n2605), .S2(n2431), .D3(n2607), .S3(n2427), .Z(n1050) );
  HS65_LH_MX41X4 U2979 ( .D0(n1017), .S0(n2417), .D1(n2605), .S1(n2424), .D2(
        n2607), .S2(n2431), .D3(n2609), .S3(n2427), .Z(n1049) );
  HS65_LH_MX41X4 U2980 ( .D0(n1016), .S0(n2417), .D1(n2607), .S1(n2424), .D2(
        n2609), .S2(n2431), .D3(n2611), .S3(n2427), .Z(n1048) );
  HS65_LH_MX41X4 U2981 ( .D0(n1015), .S0(n2417), .D1(n2609), .S1(n2424), .D2(
        n2611), .S2(n2431), .D3(n2613), .S3(n2427), .Z(n1047) );
  HS65_LH_MX41X4 U2982 ( .D0(n1014), .S0(n2417), .D1(n2611), .S1(n2424), .D2(
        n2613), .S2(n2432), .D3(n2615), .S3(n2427), .Z(n1046) );
  HS65_LH_MX41X4 U2983 ( .D0(n1012), .S0(n2417), .D1(n2615), .S1(n2424), .D2(
        n2617), .S2(n2432), .D3(n2619), .S3(n2427), .Z(n1045) );
  HS65_LH_MX41X4 U2984 ( .D0(n1011), .S0(n2417), .D1(n2617), .S1(n2424), .D2(
        n2619), .S2(n2432), .D3(n2621), .S3(n2427), .Z(n1044) );
  HS65_LH_MX41X4 U2985 ( .D0(n1010), .S0(n2417), .D1(n2619), .S1(n2424), .D2(
        n2621), .S2(n2432), .D3(n2623), .S3(n2427), .Z(n1043) );
  HS65_LH_MX41X4 U2986 ( .D0(n1009), .S0(n2417), .D1(n2621), .S1(n2423), .D2(
        n2623), .S2(n2431), .D3(n2625), .S3(n2428), .Z(n1042) );
  HS65_LH_MX41X4 U2987 ( .D0(n1008), .S0(n2418), .D1(n2623), .S1(n2424), .D2(
        n2625), .S2(n2430), .D3(n2428), .S3(n2626), .Z(n1041) );
  HS65_LH_NOR2AX3 U2988 ( .A(n3093), .B(a[31]), .Z(n2660) );
  HS65_LH_NOR2AX3 U2989 ( .A(n3094), .B(n3093), .Z(n2661) );
  HS65_LH_NOR3AX2 U2990 ( .A(a[31]), .B(n3094), .C(n3093), .Z(n2659) );
  HS65_LHS_XOR2X3 U2991 ( .A(a[31]), .B(a[30]), .Z(n3094) );
  HS65_LH_NAND2X2 U2992 ( .A(a[31]), .B(n3093), .Z(n2662) );
  HS65_LHS_XOR2X3 U2993 ( .A(n2645), .B(a[30]), .Z(n3093) );
endmodule


module alu ( clk, rst_n, .alu_i({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , 
        \alu_i[SRC_B][31] , \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , 
        \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , 
        \alu_i[SRC_B][25] , \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , 
        \alu_i[SRC_B][22] , \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , 
        \alu_i[SRC_B][19] , \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , 
        \alu_i[SRC_B][16] , \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , 
        \alu_i[SRC_B][13] , \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , 
        \alu_i[SRC_B][10] , \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , 
        \alu_i[SRC_B][7] , \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , 
        \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , 
        \alu_i[SRC_B][1] , \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , 
        \alu_i[OP][2] , \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , 
        \alu_i[SHAMT][3] , \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , 
        \alu_i[SHAMT][0] }), .alu_o({\alu_o[BRANCH] , \alu_o[RESULT][31] , 
        \alu_o[RESULT][30] , \alu_o[RESULT][29] , \alu_o[RESULT][28] , 
        \alu_o[RESULT][27] , \alu_o[RESULT][26] , \alu_o[RESULT][25] , 
        \alu_o[RESULT][24] , \alu_o[RESULT][23] , \alu_o[RESULT][22] , 
        \alu_o[RESULT][21] , \alu_o[RESULT][20] , \alu_o[RESULT][19] , 
        \alu_o[RESULT][18] , \alu_o[RESULT][17] , \alu_o[RESULT][16] , 
        \alu_o[RESULT][15] , \alu_o[RESULT][14] , \alu_o[RESULT][13] , 
        \alu_o[RESULT][12] , \alu_o[RESULT][11] , \alu_o[RESULT][10] , 
        \alu_o[RESULT][9] , \alu_o[RESULT][8] , \alu_o[RESULT][7] , 
        \alu_o[RESULT][6] , \alu_o[RESULT][5] , \alu_o[RESULT][4] , 
        \alu_o[RESULT][3] , \alu_o[RESULT][2] , \alu_o[RESULT][1] , 
        \alu_o[RESULT][0] }) );
  input clk, rst_n, \alu_i[SRC_A][31] , \alu_i[SRC_A][30] , \alu_i[SRC_A][29] ,
         \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , \alu_i[SRC_A][26] ,
         \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , \alu_i[SRC_A][23] ,
         \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , \alu_i[SRC_A][20] ,
         \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , \alu_i[SRC_A][17] ,
         \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , \alu_i[SRC_A][14] ,
         \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , \alu_i[SRC_A][11] ,
         \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , \alu_i[SRC_A][8] ,
         \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , \alu_i[SRC_A][5] ,
         \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , \alu_i[SRC_A][2] ,
         \alu_i[SRC_A][1] , \alu_i[SRC_A][0] , \alu_i[SRC_B][31] ,
         \alu_i[SRC_B][30] , \alu_i[SRC_B][29] , \alu_i[SRC_B][28] ,
         \alu_i[SRC_B][27] , \alu_i[SRC_B][26] , \alu_i[SRC_B][25] ,
         \alu_i[SRC_B][24] , \alu_i[SRC_B][23] , \alu_i[SRC_B][22] ,
         \alu_i[SRC_B][21] , \alu_i[SRC_B][20] , \alu_i[SRC_B][19] ,
         \alu_i[SRC_B][18] , \alu_i[SRC_B][17] , \alu_i[SRC_B][16] ,
         \alu_i[SRC_B][15] , \alu_i[SRC_B][14] , \alu_i[SRC_B][13] ,
         \alu_i[SRC_B][12] , \alu_i[SRC_B][11] , \alu_i[SRC_B][10] ,
         \alu_i[SRC_B][9] , \alu_i[SRC_B][8] , \alu_i[SRC_B][7] ,
         \alu_i[SRC_B][6] , \alu_i[SRC_B][5] , \alu_i[SRC_B][4] ,
         \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , \alu_i[SRC_B][1] ,
         \alu_i[SRC_B][0] , \alu_i[OP][4] , \alu_i[OP][3] , \alu_i[OP][2] ,
         \alu_i[OP][1] , \alu_i[OP][0] , \alu_i[SHAMT][4] , \alu_i[SHAMT][3] ,
         \alu_i[SHAMT][2] , \alu_i[SHAMT][1] , \alu_i[SHAMT][0] ;
  output \alu_o[BRANCH] , \alu_o[RESULT][31] , \alu_o[RESULT][30] ,
         \alu_o[RESULT][29] , \alu_o[RESULT][28] , \alu_o[RESULT][27] ,
         \alu_o[RESULT][26] , \alu_o[RESULT][25] , \alu_o[RESULT][24] ,
         \alu_o[RESULT][23] , \alu_o[RESULT][22] , \alu_o[RESULT][21] ,
         \alu_o[RESULT][20] , \alu_o[RESULT][19] , \alu_o[RESULT][18] ,
         \alu_o[RESULT][17] , \alu_o[RESULT][16] , \alu_o[RESULT][15] ,
         \alu_o[RESULT][14] , \alu_o[RESULT][13] , \alu_o[RESULT][12] ,
         \alu_o[RESULT][11] , \alu_o[RESULT][10] , \alu_o[RESULT][9] ,
         \alu_o[RESULT][8] , \alu_o[RESULT][7] , \alu_o[RESULT][6] ,
         \alu_o[RESULT][5] , \alu_o[RESULT][4] , \alu_o[RESULT][3] ,
         \alu_o[RESULT][2] , \alu_o[RESULT][1] , \alu_o[RESULT][0] ;
  wire   \HI_LO_c[HI][31] , \HI_LO_c[HI][30] , \HI_LO_c[HI][29] ,
         \HI_LO_c[HI][28] , \HI_LO_c[HI][27] , \HI_LO_c[HI][26] ,
         \HI_LO_c[HI][25] , \HI_LO_c[HI][24] , \HI_LO_c[HI][23] ,
         \HI_LO_c[HI][22] , \HI_LO_c[HI][21] , \HI_LO_c[HI][20] ,
         \HI_LO_c[HI][19] , \HI_LO_c[HI][18] , \HI_LO_c[HI][17] ,
         \HI_LO_c[HI][16] , \HI_LO_c[HI][15] , \HI_LO_c[HI][14] ,
         \HI_LO_c[HI][13] , \HI_LO_c[HI][12] , \HI_LO_c[HI][11] ,
         \HI_LO_c[HI][10] , \HI_LO_c[HI][9] , \HI_LO_c[HI][8] ,
         \HI_LO_c[HI][7] , \HI_LO_c[HI][6] , \HI_LO_c[HI][5] ,
         \HI_LO_c[HI][4] , \HI_LO_c[HI][3] , \HI_LO_c[HI][2] ,
         \HI_LO_c[HI][1] , \HI_LO_c[HI][0] , \HI_LO_c[LO][31] ,
         \HI_LO_c[LO][30] , \HI_LO_c[LO][29] , \HI_LO_c[LO][28] ,
         \HI_LO_c[LO][27] , \HI_LO_c[LO][26] , \HI_LO_c[LO][25] ,
         \HI_LO_c[LO][24] , \HI_LO_c[LO][23] , \HI_LO_c[LO][22] ,
         \HI_LO_c[LO][21] , \HI_LO_c[LO][20] , \HI_LO_c[LO][19] ,
         \HI_LO_c[LO][18] , \HI_LO_c[LO][17] , \HI_LO_c[LO][16] ,
         \HI_LO_c[LO][15] , \HI_LO_c[LO][14] , \HI_LO_c[LO][13] ,
         \HI_LO_c[LO][12] , \HI_LO_c[LO][11] , \HI_LO_c[LO][10] ,
         \HI_LO_c[LO][9] , \HI_LO_c[LO][8] , \HI_LO_c[LO][7] ,
         \HI_LO_c[LO][6] , \HI_LO_c[LO][5] , \HI_LO_c[LO][4] ,
         \HI_LO_c[LO][3] , \HI_LO_c[LO][2] , \HI_LO_c[LO][1] ,
         \HI_LO_c[LO][0] , N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N648, N649,
         N714, N715, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n300, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594;

  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][31]  ( .D(n516), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][30]  ( .D(n515), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][29]  ( .D(n514), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][28]  ( .D(n513), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][27]  ( .D(n512), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][26]  ( .D(n511), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][25]  ( .D(n510), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][24]  ( .D(n509), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][23]  ( .D(n508), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][22]  ( .D(n507), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][21]  ( .D(n506), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][20]  ( .D(n505), .CP(clk), .RN(n538), .Q(
        \HI_LO_c[HI][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][19]  ( .D(n504), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][18]  ( .D(n503), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][17]  ( .D(n502), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][16]  ( .D(n501), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][15]  ( .D(n500), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][14]  ( .D(n499), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][13]  ( .D(n498), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][12]  ( .D(n497), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][11]  ( .D(n496), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][10]  ( .D(n495), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][9]  ( .D(n494), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][8]  ( .D(n493), .CP(clk), .RN(n539), .Q(
        \HI_LO_c[HI][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][7]  ( .D(n492), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][6]  ( .D(n491), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][5]  ( .D(n490), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][4]  ( .D(n489), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][3]  ( .D(n488), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][2]  ( .D(n487), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][1]  ( .D(n486), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[HI][0]  ( .D(n485), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[HI][0] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][31]  ( .D(n484), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[LO][31] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][30]  ( .D(n483), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[LO][30] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][29]  ( .D(n482), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[LO][29] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][28]  ( .D(n481), .CP(clk), .RN(n540), .Q(
        \HI_LO_c[LO][28] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][27]  ( .D(n480), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][27] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][26]  ( .D(n479), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][26] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][25]  ( .D(n478), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][25] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][24]  ( .D(n477), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][24] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][23]  ( .D(n476), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][23] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][22]  ( .D(n475), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][22] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][21]  ( .D(n474), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][21] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][20]  ( .D(n473), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][20] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][19]  ( .D(n472), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][19] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][18]  ( .D(n471), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][18] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][17]  ( .D(n470), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][17] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][16]  ( .D(n469), .CP(clk), .RN(n541), .Q(
        \HI_LO_c[LO][16] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][15]  ( .D(n468), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][15] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][14]  ( .D(n467), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][14] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][13]  ( .D(n466), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][13] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][12]  ( .D(n465), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][12] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][11]  ( .D(n464), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][11] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][10]  ( .D(n463), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][10] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][9]  ( .D(n462), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][9] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][8]  ( .D(n461), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][8] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][7]  ( .D(n460), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][7] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][6]  ( .D(n459), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][6] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][5]  ( .D(n458), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][5] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][4]  ( .D(n457), .CP(clk), .RN(n542), .Q(
        \HI_LO_c[LO][4] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][3]  ( .D(n456), .CP(clk), .RN(n543), .Q(
        \HI_LO_c[LO][3] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][2]  ( .D(n455), .CP(clk), .RN(n543), .Q(
        \HI_LO_c[LO][2] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][1]  ( .D(n454), .CP(clk), .RN(n543), .Q(
        \HI_LO_c[LO][1] ) );
  HS65_LH_DFPRQX9 \HI_LO_c_reg[LO][0]  ( .D(n453), .CP(clk), .RN(n543), .Q(
        \HI_LO_c[LO][0] ) );
  alu_DW_cmp_0 lt_136 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({
        \alu_i[SRC_B][31] , n524, n523, \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , 
        n520, n519, n518, n517, n300, n90, \alu_i[SRC_B][20] , n88, n87, n86, 
        n85, n84, n83, n82, n81, \alu_i[SRC_B][11] , n79, n78, n77, n76, n75, 
        n74, \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , n70, n69}), .TC(1'b1), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N648) );
  alu_DW01_sub_0 sub_68 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({
        \alu_i[SRC_B][31] , n524, n523, \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , 
        n520, n519, n518, n517, n300, n90, \alu_i[SRC_B][20] , n88, n87, n86, 
        n85, n84, n83, n82, n81, \alu_i[SRC_B][11] , n79, n78, n77, n76, n75, 
        n74, \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , n70, n69}), .CI(1'b0), .DIFF({N162, N161, N160, N159, N158, N157, N156, N155, N154, 
        N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, 
        N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131}) );
  alu_DW01_cmp6_0 r325 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({
        \alu_i[SRC_B][31] , n524, n523, \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , 
        n520, n519, n518, n517, n300, n90, \alu_i[SRC_B][20] , n88, n87, n86, 
        n85, n84, n83, n82, n81, \alu_i[SRC_B][11] , n79, n78, n77, n76, n75, 
        n74, \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , n70, n69}), .TC(1'b0), .LT(N649), .EQ(N714), .NE(N715) );
  alu_DW01_add_0 r321 ( .A({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .B({
        \alu_i[SRC_B][31] , n524, n523, \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , 
        n520, n519, n518, n517, n300, n90, \alu_i[SRC_B][20] , n88, n87, n86, 
        n85, n84, n83, n82, n81, \alu_i[SRC_B][11] , n79, n78, n77, n76, n75, 
        n74, \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , n70, n69}), .CI(1'b0), .SUM({N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99}) );
  alu_DW_mult_uns_0 mult_71 ( .a({\alu_i[SRC_A][31] , \alu_i[SRC_A][30] , 
        \alu_i[SRC_A][29] , \alu_i[SRC_A][28] , \alu_i[SRC_A][27] , 
        \alu_i[SRC_A][26] , \alu_i[SRC_A][25] , \alu_i[SRC_A][24] , 
        \alu_i[SRC_A][23] , \alu_i[SRC_A][22] , \alu_i[SRC_A][21] , 
        \alu_i[SRC_A][20] , \alu_i[SRC_A][19] , \alu_i[SRC_A][18] , 
        \alu_i[SRC_A][17] , \alu_i[SRC_A][16] , \alu_i[SRC_A][15] , 
        \alu_i[SRC_A][14] , \alu_i[SRC_A][13] , \alu_i[SRC_A][12] , 
        \alu_i[SRC_A][11] , \alu_i[SRC_A][10] , \alu_i[SRC_A][9] , 
        \alu_i[SRC_A][8] , \alu_i[SRC_A][7] , \alu_i[SRC_A][6] , 
        \alu_i[SRC_A][5] , \alu_i[SRC_A][4] , \alu_i[SRC_A][3] , 
        \alu_i[SRC_A][2] , \alu_i[SRC_A][1] , \alu_i[SRC_A][0] }), .b({
        \alu_i[SRC_B][31] , n524, n523, \alu_i[SRC_B][28] , \alu_i[SRC_B][27] , 
        n520, n519, n518, n517, n300, n90, \alu_i[SRC_B][20] , n88, n87, n86, 
        n85, n84, n83, n82, n81, \alu_i[SRC_B][11] , n79, n78, n77, n76, n75, 
        n74, \alu_i[SRC_B][4] , \alu_i[SRC_B][3] , \alu_i[SRC_B][2] , n70, n69}), .product({N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, 
        N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, 
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163}) );
  HS65_LH_NOR4ABX2 U3 ( .A(n92), .B(n93), .C(n94), .D(n95), .Z(n91) );
  HS65_LH_NOR2X6 U4 ( .A(n98), .B(\alu_i[SHAMT][4] ), .Z(n284) );
  HS65_LH_BFX9 U5 ( .A(\alu_i[SRC_B][9] ), .Z(n78) );
  HS65_LH_BFX9 U6 ( .A(\alu_i[SRC_B][6] ), .Z(n75) );
  HS65_LH_BFX9 U7 ( .A(\alu_i[SRC_B][14] ), .Z(n83) );
  HS65_LH_BFX9 U13 ( .A(\alu_i[SRC_B][10] ), .Z(n79) );
  HS65_LH_BFX9 U14 ( .A(\alu_i[SRC_B][8] ), .Z(n77) );
  HS65_LH_BFX9 U15 ( .A(\alu_i[SRC_B][7] ), .Z(n76) );
  HS65_LH_BFX9 U16 ( .A(\alu_i[SRC_B][15] ), .Z(n84) );
  HS65_LH_BFX9 U17 ( .A(\alu_i[SRC_B][5] ), .Z(n74) );
  HS65_LH_BFX9 U18 ( .A(\alu_i[SRC_B][13] ), .Z(n82) );
  HS65_LH_BFX9 U19 ( .A(\alu_i[SRC_B][12] ), .Z(n81) );
  HS65_LH_BFX9 U20 ( .A(\alu_i[SRC_B][25] ), .Z(n519) );
  HS65_LH_BFX9 U21 ( .A(\alu_i[SRC_B][16] ), .Z(n85) );
  HS65_LH_BFX9 U22 ( .A(\alu_i[SRC_B][26] ), .Z(n520) );
  HS65_LH_BFX9 U23 ( .A(\alu_i[SRC_B][17] ), .Z(n86) );
  HS65_LH_BFX9 U24 ( .A(\alu_i[SRC_B][1] ), .Z(n70) );
  HS65_LH_BFX9 U25 ( .A(\alu_i[SRC_B][18] ), .Z(n87) );
  HS65_LH_BFX9 U26 ( .A(\alu_i[SRC_B][21] ), .Z(n90) );
  HS65_LH_BFX9 U27 ( .A(\alu_i[SRC_B][29] ), .Z(n523) );
  HS65_LH_BFX9 U28 ( .A(\alu_i[SRC_B][22] ), .Z(n300) );
  HS65_LH_BFX9 U29 ( .A(\alu_i[SRC_B][24] ), .Z(n518) );
  HS65_LH_BFX9 U30 ( .A(\alu_i[SRC_B][30] ), .Z(n524) );
  HS65_LH_BFX9 U31 ( .A(\alu_i[SRC_B][19] ), .Z(n88) );
  HS65_LH_BFX9 U32 ( .A(\alu_i[SRC_B][23] ), .Z(n517) );
  HS65_LH_OR2X9 U33 ( .A(\alu_i[SHAMT][2] ), .B(\alu_i[SHAMT][3] ), .Z(n6) );
  HS65_LH_IVX9 U34 ( .A(n61), .Z(n60) );
  HS65_LH_IVX9 U35 ( .A(n62), .Z(n59) );
  HS65_LH_IVX9 U36 ( .A(n62), .Z(n58) );
  HS65_LH_IVX9 U37 ( .A(n62), .Z(n57) );
  HS65_LH_IVX9 U38 ( .A(n98), .Z(n581) );
  HS65_LH_IVX9 U39 ( .A(n176), .Z(n580) );
  HS65_LH_IVX9 U40 ( .A(n281), .Z(n582) );
  HS65_LH_IVX9 U41 ( .A(n56), .Z(n55) );
  HS65_LH_IVX9 U42 ( .A(n42), .Z(n41) );
  HS65_LH_BFX9 U43 ( .A(n68), .Z(n61) );
  HS65_LH_BFX9 U44 ( .A(n68), .Z(n62) );
  HS65_LH_BFX9 U45 ( .A(n586), .Z(n15) );
  HS65_LH_BFX9 U46 ( .A(n586), .Z(n14) );
  HS65_LH_BFX9 U47 ( .A(n585), .Z(n11) );
  HS65_LH_BFX9 U48 ( .A(n585), .Z(n12) );
  HS65_LH_BFX9 U49 ( .A(n67), .Z(n65) );
  HS65_LH_BFX9 U50 ( .A(n67), .Z(n64) );
  HS65_LH_BFX9 U51 ( .A(n68), .Z(n63) );
  HS65_LH_BFX9 U52 ( .A(n586), .Z(n16) );
  HS65_LH_BFX9 U53 ( .A(n585), .Z(n13) );
  HS65_LH_BFX9 U54 ( .A(n67), .Z(n66) );
  HS65_LH_IVX9 U55 ( .A(n101), .Z(n585) );
  HS65_LH_IVX9 U56 ( .A(n100), .Z(n586) );
  HS65_LH_NOR2X6 U57 ( .A(n96), .B(n189), .Z(n279) );
  HS65_LH_AOI222X2 U58 ( .A(n275), .B(n276), .C(n277), .D(n278), .E(n279), .F(
        n214), .Z(n274) );
  HS65_LH_NAND2X7 U59 ( .A(n442), .B(n435), .Z(n98) );
  HS65_LH_IVX9 U60 ( .A(n96), .Z(n584) );
  HS65_LH_NOR2X6 U61 ( .A(n189), .B(n98), .Z(n115) );
  HS65_LH_IVX9 U62 ( .A(n208), .Z(n579) );
  HS65_LH_IVX9 U63 ( .A(n186), .Z(n583) );
  HS65_LH_NAND2X7 U64 ( .A(n195), .B(n581), .Z(n176) );
  HS65_LH_NAND2X7 U65 ( .A(n584), .B(n195), .Z(n281) );
  HS65_LH_OAI211X5 U66 ( .A(n39), .B(n208), .C(n101), .D(n40), .Z(n207) );
  HS65_LH_NOR3X4 U67 ( .A(n48), .B(n45), .C(n106), .Z(n92) );
  HS65_LH_IVX9 U68 ( .A(n189), .Z(n591) );
  HS65_LH_IVX9 U69 ( .A(n237), .Z(n576) );
  HS65_LH_AND2X4 U70 ( .A(n275), .B(n17), .Z(n368) );
  HS65_LH_AND2X4 U71 ( .A(n117), .B(n17), .Z(n397) );
  HS65_LH_IVX9 U72 ( .A(n54), .Z(n56) );
  HS65_LH_IVX9 U73 ( .A(n40), .Z(n42) );
  HS65_LH_BFX9 U74 ( .A(n43), .Z(n44) );
  HS65_LH_BFX9 U75 ( .A(n91), .Z(n68) );
  HS65_LH_BFX9 U76 ( .A(n91), .Z(n67) );
  HS65_LH_BFX9 U77 ( .A(n50), .Z(n52) );
  HS65_LH_BFX9 U78 ( .A(n50), .Z(n51) );
  HS65_LH_IVX9 U79 ( .A(n39), .Z(n37) );
  HS65_LH_BFX9 U80 ( .A(n577), .Z(n10) );
  HS65_LH_BFX9 U81 ( .A(n30), .Z(n32) );
  HS65_LH_BFX9 U82 ( .A(n577), .Z(n9) );
  HS65_LH_BFX9 U83 ( .A(n43), .Z(n45) );
  HS65_LH_BFX9 U84 ( .A(n30), .Z(n33) );
  HS65_LH_BFX9 U85 ( .A(n31), .Z(n34) );
  HS65_LH_IVX9 U86 ( .A(n39), .Z(n38) );
  HS65_LH_BFX9 U87 ( .A(n19), .Z(n21) );
  HS65_LH_BFX9 U88 ( .A(n19), .Z(n23) );
  HS65_LH_BFX9 U89 ( .A(n19), .Z(n22) );
  HS65_LH_BFX9 U90 ( .A(n20), .Z(n24) );
  HS65_LH_IVX9 U91 ( .A(n317), .Z(n572) );
  HS65_LH_BFX9 U92 ( .A(n50), .Z(n53) );
  HS65_LH_IVX9 U93 ( .A(n144), .Z(n569) );
  HS65_LH_IVX9 U94 ( .A(n130), .Z(n571) );
  HS65_LH_IVX9 U95 ( .A(n212), .Z(n570) );
  HS65_LH_BFX9 U96 ( .A(n20), .Z(n25) );
  HS65_LH_BFX9 U97 ( .A(n31), .Z(n35) );
  HS65_LH_NAND4ABX3 U98 ( .A(n42), .B(n53), .C(n578), .D(n10), .Z(n94) );
  HS65_LH_NAND3X5 U99 ( .A(n96), .B(n55), .C(n98), .Z(n95) );
  HS65_LH_NOR4ABX2 U100 ( .A(n100), .B(n101), .C(n102), .D(n103), .Z(n93) );
  HS65_LH_IVX9 U101 ( .A(n180), .Z(n577) );
  HS65_LH_AOI222X2 U102 ( .A(n32), .B(n70), .C(n27), .D(n69), .E(n196), .F(
        \alu_i[SRC_B][2] ), .Z(n237) );
  HS65_LH_NOR2X6 U103 ( .A(n592), .B(n96), .Z(n275) );
  HS65_LH_NAND2X7 U104 ( .A(n436), .B(n442), .Z(n96) );
  HS65_LH_AOI222X2 U105 ( .A(n284), .B(n387), .C(n277), .D(n314), .E(n279), 
        .F(n317), .Z(n386) );
  HS65_LH_AOI222X2 U106 ( .A(n284), .B(n360), .C(n277), .D(n302), .E(n279), 
        .F(n306), .Z(n380) );
  HS65_LH_AOI222X2 U107 ( .A(n284), .B(n239), .C(n277), .D(n336), .E(n279), 
        .F(n292), .Z(n373) );
  HS65_LH_AOI222X2 U108 ( .A(n284), .B(n566), .C(n277), .D(n326), .E(n279), 
        .F(n278), .Z(n366) );
  HS65_LH_IVX9 U109 ( .A(n190), .Z(n566) );
  HS65_LH_AOI222X2 U110 ( .A(n284), .B(n174), .C(n277), .D(n316), .E(n279), 
        .F(n266), .Z(n349) );
  HS65_LH_AOI222X2 U111 ( .A(n275), .B(n165), .C(n279), .D(n254), .E(n284), 
        .F(n166), .Z(n343) );
  HS65_LH_AOI222X2 U112 ( .A(n275), .B(n153), .C(n279), .D(n229), .E(n284), 
        .F(n155), .Z(n333) );
  HS65_LH_AOI222X2 U113 ( .A(n275), .B(n141), .C(n279), .D(n212), .E(n284), 
        .F(n143), .Z(n323) );
  HS65_LH_AOI222X2 U114 ( .A(n275), .B(n129), .C(n279), .D(n268), .E(n284), 
        .F(n131), .Z(n312) );
  HS65_LH_AOI222X2 U115 ( .A(n275), .B(n112), .C(n279), .D(n256), .E(n284), 
        .F(n116), .Z(n298) );
  HS65_LH_AOI222X2 U116 ( .A(n275), .B(n290), .C(n279), .D(n231), .E(n284), 
        .F(n291), .Z(n289) );
  HS65_LH_AOI212X4 U117 ( .A(\alu_i[SRC_A][11] ), .B(n180), .C(n56), .D(n529), 
        .E(n42), .Z(n421) );
  HS65_LH_AOI212X4 U118 ( .A(\alu_i[SRC_A][20] ), .B(n180), .C(n56), .D(n532), 
        .E(n42), .Z(n350) );
  HS65_LH_NAND2X7 U119 ( .A(n301), .B(n592), .Z(n189) );
  HS65_LH_OAI212X5 U120 ( .A(n574), .B(n189), .C(n190), .D(n592), .E(n191), 
        .Z(n183) );
  HS65_LH_IVX9 U121 ( .A(n140), .Z(n574) );
  HS65_LH_AOI222X2 U122 ( .A(n192), .B(n145), .C(n193), .D(n194), .E(n195), 
        .F(n142), .Z(n191) );
  HS65_LH_MX41X7 U123 ( .D0(\alu_i[SRC_B][3] ), .S0(n37), .D1(
        \alu_i[SRC_B][4] ), .S1(n33), .D2(n74), .S2(n28), .D3(n75), .S3(n23), 
        .Z(n194) );
  HS65_LH_OAI212X5 U124 ( .A(n568), .B(n189), .C(n264), .D(n592), .E(n265), 
        .Z(n259) );
  HS65_LH_IVX9 U125 ( .A(n269), .Z(n568) );
  HS65_LH_AOI222X2 U126 ( .A(n192), .B(n266), .C(n193), .D(n267), .E(n195), 
        .F(n268), .Z(n265) );
  HS65_LH_MX41X7 U127 ( .D0(\alu_i[SRC_B][28] ), .S0(n36), .D1(
        \alu_i[SRC_B][27] ), .S1(n32), .D2(n520), .S2(n27), .D3(n519), .S3(n21), .Z(n267) );
  HS65_LH_OAI212X5 U128 ( .A(n236), .B(n71), .C(n237), .D(n186), .E(n238), .Z(
        n235) );
  HS65_LH_CBI4I1X5 U129 ( .A(n56), .B(n71), .C(n42), .D(\alu_i[SRC_A][2] ), 
        .Z(n238) );
  HS65_LH_AOI212X4 U130 ( .A(\alu_i[SRC_A][2] ), .B(n180), .C(n56), .D(n526), 
        .E(n42), .Z(n236) );
  HS65_LH_NOR2X6 U131 ( .A(n594), .B(n593), .Z(n374) );
  HS65_LH_OAI212X5 U132 ( .A(\alu_i[SRC_A][29] ), .B(n55), .C(n9), .D(n535), 
        .E(n41), .Z(n248) );
  HS65_LH_NOR2X6 U133 ( .A(n592), .B(n98), .Z(n117) );
  HS65_LH_OAI212X5 U134 ( .A(\alu_i[SRC_A][14] ), .B(n54), .C(n10), .D(n530), 
        .E(n123), .Z(n403) );
  HS65_LH_OAI212X5 U135 ( .A(\alu_i[SRC_A][17] ), .B(n54), .C(n10), .D(n531), 
        .E(n40), .Z(n381) );
  HS65_LH_OAI212X5 U136 ( .A(\alu_i[SRC_A][5] ), .B(n55), .C(n9), .D(n527), 
        .E(n41), .Z(n167) );
  HS65_LH_OAI212X5 U137 ( .A(\alu_i[SRC_A][8] ), .B(n55), .C(n9), .D(n528), 
        .E(n41), .Z(n134) );
  HS65_LH_OAI212X5 U138 ( .A(\alu_i[SRC_A][23] ), .B(n55), .C(n9), .D(n533), 
        .E(n41), .Z(n328) );
  HS65_LH_OAI212X5 U139 ( .A(\alu_i[SRC_A][26] ), .B(n55), .C(n9), .D(n534), 
        .E(n41), .Z(n293) );
  HS65_LH_AOI32X5 U140 ( .A(n178), .B(n593), .C(n275), .D(\alu_i[SRC_A][20] ), 
        .E(n352), .Z(n351) );
  HS65_LH_OAI21X3 U141 ( .A(\alu_i[SRC_B][20] ), .B(n54), .C(n40), .Z(n352) );
  HS65_LH_AND2X4 U142 ( .A(n192), .B(n584), .Z(n277) );
  HS65_LH_NOR2X6 U143 ( .A(n588), .B(n590), .Z(n435) );
  HS65_LH_AOI32X5 U144 ( .A(n283), .B(n593), .C(n117), .D(\alu_i[SRC_A][11] ), 
        .E(n423), .Z(n422) );
  HS65_LH_OAI21X3 U145 ( .A(\alu_i[SRC_B][11] ), .B(n54), .C(n123), .Z(n423)
         );
  HS65_LH_NAND2X7 U146 ( .A(n193), .B(n581), .Z(n208) );
  HS65_LH_MX41X7 U147 ( .D0(n81), .S0(n38), .D1(\alu_i[SRC_B][11] ), .S1(n34), 
        .D2(n79), .S2(n29), .D3(n21), .S3(n78), .Z(n317) );
  HS65_LH_AND2X4 U148 ( .A(n390), .B(n391), .Z(n106) );
  HS65_LH_MX41X7 U149 ( .D0(n77), .S0(n38), .D1(n76), .S1(n34), .D2(n75), .S2(
        n28), .D3(n74), .S3(n23), .Z(n316) );
  HS65_LH_MX41X7 U150 ( .D0(n84), .S0(n38), .D1(n85), .S1(n34), .D2(n86), .S2(
        n29), .D3(n87), .S3(n24), .Z(n145) );
  HS65_LH_MX41X7 U151 ( .D0(n85), .S0(n37), .D1(n84), .S1(n33), .D2(n83), .S2(
        n28), .D3(n82), .S3(n22), .Z(n266) );
  HS65_LH_MX41X7 U152 ( .D0(n84), .S0(n37), .D1(n83), .S1(n33), .D2(n82), .S2(
        n28), .D3(n81), .S3(n22), .Z(n278) );
  HS65_LH_NOR2AX3 U153 ( .A(n69), .B(n39), .Z(n315) );
  HS65_LH_MX41X7 U154 ( .D0(n196), .S0(n88), .D1(n32), .S1(\alu_i[SRC_B][20] ), 
        .D2(n90), .S2(n29), .D3(n300), .S3(n24), .Z(n144) );
  HS65_LH_MX41X7 U155 ( .D0(\alu_i[SRC_B][28] ), .S0(n38), .D1(n523), .S1(n34), 
        .D2(n524), .S2(n29), .D3(\alu_i[SRC_B][31] ), .S3(n25), .Z(n263) );
  HS65_LH_MX41X7 U156 ( .D0(\alu_i[SRC_B][3] ), .S0(n38), .D1(
        \alu_i[SRC_B][2] ), .S1(n34), .D2(n70), .S2(n29), .D3(n69), .S3(n24), 
        .Z(n188) );
  HS65_LH_NAND2X7 U157 ( .A(n193), .B(n584), .Z(n186) );
  HS65_LH_MX41X7 U158 ( .D0(n81), .S0(n38), .D1(n82), .S1(n34), .D2(n83), .S2(
        n29), .D3(n84), .S3(n25), .Z(n130) );
  HS65_LH_MX41X7 U159 ( .D0(n36), .S0(n88), .D1(n87), .S1(n33), .D2(n86), .S2(
        n28), .D3(n85), .S3(n22), .Z(n212) );
  HS65_LH_MX41X7 U160 ( .D0(n517), .S0(n38), .D1(n518), .S1(n34), .D2(n519), 
        .S2(n29), .D3(n520), .S3(n24), .Z(n325) );
  HS65_LH_MX41X7 U161 ( .D0(n83), .S0(n38), .D1(n84), .S1(n34), .D2(n85), .S2(
        n29), .D3(n86), .S3(n24), .Z(n157) );
  HS65_LH_MX41X7 U162 ( .D0(n82), .S0(n37), .D1(n83), .S1(n33), .D2(n84), .S2(
        n28), .D3(n85), .S3(n23), .Z(n114) );
  HS65_LH_MX41X7 U163 ( .D0(\alu_i[SRC_B][11] ), .S0(n38), .D1(n81), .S1(n34), 
        .D2(n82), .S2(n29), .D3(n83), .S3(n23), .Z(n142) );
  HS65_LH_MX41X7 U164 ( .D0(n74), .S0(n37), .D1(\alu_i[SRC_B][4] ), .S1(n33), 
        .D2(\alu_i[SRC_B][3] ), .S2(n28), .D3(\alu_i[SRC_B][2] ), .S3(n23), 
        .Z(n302) );
  HS65_LH_MX41X7 U165 ( .D0(n75), .S0(n38), .D1(n74), .S1(n34), .D2(
        \alu_i[SRC_B][4] ), .S2(n29), .D3(\alu_i[SRC_B][3] ), .S3(n24), .Z(
        n336) );
  HS65_LH_MX41X7 U166 ( .D0(n76), .S0(n38), .D1(n75), .S1(n34), .D2(n74), .S2(
        n29), .D3(\alu_i[SRC_B][4] ), .S3(n24), .Z(n326) );
  HS65_LH_MX41X7 U167 ( .D0(n196), .S0(n87), .D1(n86), .S1(n33), .D2(n85), 
        .S2(n28), .D3(n84), .S3(n22), .Z(n229) );
  HS65_LH_MX41X7 U168 ( .D0(n36), .S0(\alu_i[SRC_B][20] ), .D1(n32), .S1(n88), 
        .D2(n87), .S2(n28), .D3(n86), .S3(n22), .Z(n268) );
  HS65_LH_AND2X4 U169 ( .A(n445), .B(n587), .Z(n442) );
  HS65_LH_MX41X7 U170 ( .D0(n86), .S0(n37), .D1(n85), .S1(n33), .D2(n84), .S2(
        n28), .D3(n83), .S3(n22), .Z(n254) );
  HS65_LH_MX41X7 U171 ( .D0(n83), .S0(n37), .D1(n82), .S1(n33), .D2(n81), .S2(
        n28), .D3(\alu_i[SRC_B][11] ), .S3(n23), .Z(n292) );
  HS65_LH_MX41X7 U172 ( .D0(n82), .S0(n37), .D1(n81), .S1(n33), .D2(
        \alu_i[SRC_B][11] ), .S2(n28), .D3(n79), .S3(n23), .Z(n306) );
  HS65_LH_CBI4I6X5 U173 ( .A(n69), .B(n55), .C(n123), .D(n565), .Z(n440) );
  HS65_LH_CBI4I6X5 U174 ( .A(n70), .B(n55), .C(n40), .D(n564), .Z(n358) );
  HS65_LH_CBI4I6X5 U175 ( .A(n523), .B(n55), .C(n123), .D(n535), .Z(n249) );
  HS65_LH_CBI4I6X5 U176 ( .A(n524), .B(n55), .C(n40), .D(n545), .Z(n224) );
  HS65_LH_AO222X4 U177 ( .A(n34), .B(n524), .C(n27), .D(\alu_i[SRC_B][31] ), 
        .E(n36), .F(n523), .Z(n247) );
  HS65_LH_AND2X4 U178 ( .A(n448), .B(n594), .Z(n195) );
  HS65_LH_MX41X7 U179 ( .D0(n518), .S0(n38), .D1(n519), .S1(n34), .D2(n520), 
        .S2(n29), .D3(\alu_i[SRC_B][27] ), .S3(n25), .Z(n313) );
  HS65_LH_MX41X7 U180 ( .D0(n196), .S0(n78), .D1(n79), .S1(n33), .D2(
        \alu_i[SRC_B][11] ), .S2(n28), .D3(n81), .S3(n22), .Z(n111) );
  HS65_LH_MX41X7 U181 ( .D0(n79), .S0(n38), .D1(\alu_i[SRC_B][11] ), .S1(n34), 
        .D2(n81), .S2(n29), .D3(n82), .S3(n24), .Z(n154) );
  HS65_LH_MX41X7 U182 ( .D0(n519), .S0(n37), .D1(n520), .S1(n33), .D2(
        \alu_i[SRC_B][27] ), .S2(n28), .D3(\alu_i[SRC_B][28] ), .S3(n23), .Z(
        n299) );
  HS65_LH_MX41X7 U183 ( .D0(n520), .S0(n38), .D1(\alu_i[SRC_B][27] ), .S1(n34), 
        .D2(\alu_i[SRC_B][28] ), .S2(n29), .D3(n523), .S3(n24), .Z(n334) );
  HS65_LH_MX41X7 U184 ( .D0(n85), .S0(n196), .D1(n86), .S1(n34), .D2(n87), 
        .S2(n29), .D3(n88), .S3(n25), .Z(n133) );
  HS65_LH_MX41X7 U185 ( .D0(n36), .S0(\alu_i[SRC_B][20] ), .D1(n90), .S1(n34), 
        .D2(n300), .S2(n29), .D3(n517), .S3(n25), .Z(n132) );
  HS65_LH_MX41X7 U186 ( .D0(n300), .S0(n37), .D1(n90), .S1(n33), .D2(n27), 
        .S2(\alu_i[SRC_B][20] ), .D3(n88), .S3(n22), .Z(n231) );
  HS65_LH_MX41X7 U187 ( .D0(n300), .S0(n38), .D1(n517), .S1(n34), .D2(n518), 
        .S2(n29), .D3(n519), .S3(n24), .Z(n335) );
  HS65_LH_MX41X7 U188 ( .D0(n79), .S0(n38), .D1(n32), .S1(n78), .D2(n77), .S2(
        n29), .D3(n76), .S3(n24), .Z(n337) );
  HS65_LH_MX41X7 U189 ( .D0(n90), .S0(n37), .D1(n300), .S1(n33), .D2(n517), 
        .S2(n28), .D3(n518), .S3(n23), .Z(n119) );
  HS65_LH_MX41X7 U190 ( .D0(n90), .S0(n37), .D1(n32), .S1(\alu_i[SRC_B][20] ), 
        .D2(n88), .S2(n27), .D3(n87), .S3(n22), .Z(n256) );
  HS65_LH_NOR2X6 U191 ( .A(n525), .B(n39), .Z(n216) );
  HS65_LH_MX41X7 U192 ( .D0(n196), .S0(n78), .D1(n77), .S1(n33), .D2(n76), 
        .S2(n28), .D3(n75), .S3(n23), .Z(n305) );
  HS65_LH_MX41X7 U193 ( .D0(\alu_i[SRC_B][11] ), .S0(n38), .D1(n79), .S1(n34), 
        .D2(n27), .S2(n78), .D3(n77), .S3(n23), .Z(n327) );
  HS65_LH_MX41X7 U194 ( .D0(\alu_i[SRC_B][4] ), .S0(n38), .D1(
        \alu_i[SRC_B][3] ), .S1(n33), .D2(\alu_i[SRC_B][2] ), .S2(n28), .D3(
        n70), .S3(n23), .Z(n314) );
  HS65_LH_MX41X7 U195 ( .D0(n86), .S0(n37), .D1(n87), .S1(n33), .D2(n88), .S2(
        n28), .D3(\alu_i[SRC_B][20] ), .S3(n23), .Z(n120) );
  HS65_LH_MX41X7 U196 ( .D0(n36), .S0(n87), .D1(n32), .S1(n88), .D2(n27), .S2(
        \alu_i[SRC_B][20] ), .D3(n90), .S3(n24), .Z(n156) );
  HS65_LH_MX41X7 U197 ( .D0(n77), .S0(n38), .D1(n32), .S1(n78), .D2(n79), .S2(
        n29), .D3(\alu_i[SRC_B][11] ), .S3(n25), .Z(n128) );
  HS65_LH_MX41X7 U198 ( .D0(n517), .S0(n37), .D1(n300), .S1(n32), .D2(n90), 
        .S2(n27), .D3(\alu_i[SRC_B][20] ), .S3(n22), .Z(n214) );
  HS65_LH_NAND2X7 U199 ( .A(n434), .B(n438), .Z(n101) );
  HS65_LH_MX41X7 U200 ( .D0(n76), .S0(n37), .D1(n77), .S1(n32), .D2(n27), .S2(
        n78), .D3(n79), .S3(n21), .Z(n140) );
  HS65_LH_AND2X4 U201 ( .A(n192), .B(n581), .Z(n118) );
  HS65_LH_AO22X9 U202 ( .A(n196), .B(n70), .C(n32), .D(n69), .Z(n303) );
  HS65_LH_AO22X9 U203 ( .A(n36), .B(n524), .C(n32), .D(\alu_i[SRC_B][31] ), 
        .Z(n222) );
  HS65_LH_MX41X7 U204 ( .D0(\alu_i[SRC_B][27] ), .S0(n38), .D1(
        \alu_i[SRC_B][28] ), .S1(n34), .D2(n523), .S2(n29), .D3(n524), .S3(n24), .Z(n324) );
  HS65_LH_MX41X7 U205 ( .D0(\alu_i[SRC_B][4] ), .S0(n196), .D1(n74), .S1(n32), 
        .D2(n75), .S2(n27), .D3(n76), .S3(n21), .Z(n173) );
  HS65_LH_MX41X7 U206 ( .D0(n17), .S0(n133), .D1(n301), .S1(n132), .D2(n304), 
        .S2(n313), .D3(n374), .S3(n263), .Z(n387) );
  HS65_LH_MX41X7 U207 ( .D0(n17), .S0(n120), .D1(n7), .S1(n119), .D2(n304), 
        .S2(n299), .D3(n374), .S3(n247), .Z(n360) );
  HS65_LH_MX41X7 U208 ( .D0(n17), .S0(n156), .D1(n8), .S1(n335), .D2(n304), 
        .S2(n334), .D3(n374), .S3(n222), .Z(n239) );
  HS65_LH_MX41X7 U209 ( .D0(n74), .S0(n37), .D1(n75), .S1(n33), .D2(n76), .S2(
        n28), .D3(n77), .S3(n22), .Z(n164) );
  HS65_LH_MX41X7 U210 ( .D0(n75), .S0(n37), .D1(n76), .S1(n32), .D2(n77), .S2(
        n27), .D3(n21), .S3(n78), .Z(n152) );
  HS65_LH_AO222X4 U211 ( .A(n313), .B(n301), .C(n263), .D(n304), .E(n132), .F(
        n17), .Z(n174) );
  HS65_LH_AO222X4 U212 ( .A(n326), .B(n8), .C(n188), .D(n304), .E(n327), .F(
        n17), .Z(n276) );
  HS65_LH_AO222X4 U213 ( .A(n314), .B(n7), .C(n304), .D(n315), .E(n316), .F(
        n18), .Z(n129) );
  HS65_LH_AO222X4 U214 ( .A(n302), .B(n8), .C(n303), .D(n304), .E(n305), .F(
        n18), .Z(n112) );
  HS65_LH_AO222X4 U215 ( .A(n336), .B(n7), .C(n576), .D(n304), .E(n337), .F(
        n17), .Z(n290) );
  HS65_LH_MX41X7 U216 ( .D0(n518), .S0(n36), .D1(n517), .S1(n33), .D2(n300), 
        .S2(n27), .D3(n90), .S3(n21), .Z(n269) );
  HS65_LH_AO222X4 U217 ( .A(n324), .B(n301), .C(n304), .D(n216), .E(n325), .F(
        n18), .Z(n143) );
  HS65_LH_AO222X4 U218 ( .A(n299), .B(n7), .C(n247), .D(n304), .E(n119), .F(
        n17), .Z(n166) );
  HS65_LH_AO222X4 U219 ( .A(n334), .B(n8), .C(n222), .D(n304), .E(n335), .F(
        n18), .Z(n155) );
  HS65_LH_MX41X7 U220 ( .D0(n520), .S0(n196), .D1(n519), .S1(n32), .D2(n518), 
        .S2(n27), .D3(n517), .S3(n21), .Z(n226) );
  HS65_LH_MX41X7 U221 ( .D0(n519), .S0(n37), .D1(n518), .S1(n32), .D2(n517), 
        .S2(n27), .D3(n300), .S3(n22), .Z(n251) );
  HS65_LH_MX41X7 U222 ( .D0(\alu_i[SRC_B][27] ), .S0(n36), .D1(n520), .S1(n32), 
        .D2(n519), .S2(n27), .D3(n518), .S3(n21), .Z(n209) );
  HS65_LH_OAI21X3 U223 ( .A(n74), .B(n97), .C(n40), .Z(n168) );
  HS65_LH_OAI21X3 U224 ( .A(n75), .B(n54), .C(n40), .Z(n159) );
  HS65_LH_OAI21X3 U225 ( .A(n76), .B(n97), .C(n123), .Z(n147) );
  HS65_LH_OAI21X3 U226 ( .A(n77), .B(n54), .C(n40), .Z(n135) );
  HS65_LH_OAI21X3 U227 ( .A(n79), .B(n97), .C(n123), .Z(n429) );
  HS65_LH_OAI21X3 U228 ( .A(n81), .B(n54), .C(n40), .Z(n416) );
  HS65_LH_OAI21X3 U229 ( .A(n82), .B(n97), .C(n123), .Z(n410) );
  HS65_LH_OAI21X3 U230 ( .A(n83), .B(n54), .C(n40), .Z(n404) );
  HS65_LH_OAI21X3 U231 ( .A(n84), .B(n97), .C(n123), .Z(n398) );
  HS65_LH_OAI21X3 U232 ( .A(n85), .B(n54), .C(n123), .Z(n389) );
  HS65_LH_OAI21X3 U233 ( .A(n86), .B(n97), .C(n40), .Z(n382) );
  HS65_LH_OAI21X3 U234 ( .A(n88), .B(n54), .C(n123), .Z(n369) );
  HS65_LH_OAI21X3 U235 ( .A(n518), .B(n97), .C(n40), .Z(n319) );
  HS65_LH_OAI21X3 U236 ( .A(n519), .B(n54), .C(n123), .Z(n308) );
  HS65_LH_OAI21X3 U237 ( .A(n520), .B(n97), .C(n40), .Z(n294) );
  HS65_LH_OAI21X3 U238 ( .A(n90), .B(n97), .C(n123), .Z(n345) );
  HS65_LH_OAI21X3 U239 ( .A(n300), .B(n54), .C(n40), .Z(n339) );
  HS65_LH_OAI21X3 U240 ( .A(n517), .B(n97), .C(n123), .Z(n329) );
  HS65_LH_MX41X7 U241 ( .D0(n17), .S0(n306), .D1(n7), .S1(n305), .D2(n304), 
        .S2(n302), .D3(n374), .S3(n303), .Z(n252) );
  HS65_LH_MX41X7 U242 ( .D0(n17), .S0(n292), .D1(n8), .S1(n337), .D2(n304), 
        .S2(n336), .D3(n374), .S3(n576), .Z(n227) );
  HS65_LH_MX41X7 U243 ( .D0(n17), .S0(n278), .D1(n301), .S1(n327), .D2(n304), 
        .S2(n326), .D3(n374), .S3(n188), .Z(n210) );
  HS65_LH_NAND2X7 U244 ( .A(n434), .B(n435), .Z(n100) );
  HS65_LH_OAI21X3 U245 ( .A(n78), .B(n97), .C(n40), .Z(n122) );
  HS65_LH_OAI21X3 U246 ( .A(n87), .B(n97), .C(n40), .Z(n376) );
  HS65_LH_IVX9 U247 ( .A(n36), .Z(n39) );
  HS65_LH_IVX9 U248 ( .A(n6), .Z(n17) );
  HS65_LH_NAND3X5 U249 ( .A(n243), .B(n244), .C(n245), .Z(\alu_o[RESULT][29] )
         );
  HS65_LH_AOI22X6 U250 ( .A(N128), .B(n48), .C(n584), .D(n250), .Z(n243) );
  HS65_LH_AOI212X4 U251 ( .A(n13), .B(n524), .C(N160), .D(n53), .E(n246), .Z(
        n245) );
  HS65_LH_AOI212X4 U252 ( .A(n579), .B(n247), .C(n523), .D(n248), .E(n249), 
        .Z(n244) );
  HS65_LH_NAND3X5 U253 ( .A(n218), .B(n219), .C(n220), .Z(\alu_o[RESULT][30] )
         );
  HS65_LH_AOI22X6 U254 ( .A(N129), .B(n48), .C(n584), .D(n225), .Z(n218) );
  HS65_LH_AOI212X4 U255 ( .A(n13), .B(\alu_i[SRC_B][31] ), .C(N161), .D(n53), 
        .E(n221), .Z(n220) );
  HS65_LH_AOI212X4 U256 ( .A(n579), .B(n222), .C(n524), .D(n223), .E(n224), 
        .Z(n219) );
  HS65_LH_NAND3X5 U257 ( .A(n353), .B(n354), .C(n355), .Z(\alu_o[RESULT][1] )
         );
  HS65_LH_AOI22X6 U258 ( .A(N100), .B(n48), .C(n581), .D(n359), .Z(n353) );
  HS65_LH_AOI212X4 U259 ( .A(n12), .B(\alu_i[SRC_B][2] ), .C(N132), .D(n53), 
        .E(n356), .Z(n355) );
  HS65_LH_AOI212X4 U260 ( .A(n583), .B(n303), .C(n70), .D(n357), .E(n358), .Z(
        n354) );
  HS65_LH_BFX9 U261 ( .A(n97), .Z(n54) );
  HS65_LH_NAND2X7 U262 ( .A(n391), .B(n442), .Z(n97) );
  HS65_LH_BFX9 U263 ( .A(n123), .Z(n40) );
  HS65_LH_NAND2X7 U264 ( .A(n438), .B(n442), .Z(n123) );
  HS65_LH_AO22X9 U265 ( .A(n302), .B(n17), .C(n303), .D(n7), .Z(n165) );
  HS65_LH_AO22X9 U266 ( .A(n336), .B(n17), .C(n576), .D(n8), .Z(n153) );
  HS65_LH_AO22X9 U267 ( .A(n326), .B(n17), .C(n188), .D(n301), .Z(n141) );
  HS65_LH_AO22X9 U268 ( .A(n313), .B(n17), .C(n263), .D(n7), .Z(n131) );
  HS65_LH_AO22X9 U269 ( .A(n299), .B(n17), .C(n247), .D(n8), .Z(n116) );
  HS65_LH_AO22X9 U270 ( .A(n334), .B(n17), .C(n222), .D(n301), .Z(n291) );
  HS65_LH_BFX9 U271 ( .A(n199), .Z(n19) );
  HS65_LH_BFX9 U272 ( .A(n105), .Z(n43) );
  HS65_LH_NOR2AX3 U273 ( .A(n390), .B(n589), .Z(n105) );
  HS65_LH_BFX9 U274 ( .A(n99), .Z(n50) );
  HS65_LH_NOR2X6 U275 ( .A(n590), .B(n437), .Z(n99) );
  HS65_LH_BFX9 U276 ( .A(n46), .Z(n48) );
  HS65_LH_IVX9 U277 ( .A(n438), .Z(n589) );
  HS65_LH_BFX9 U278 ( .A(n46), .Z(n47) );
  HS65_LH_AND2X4 U279 ( .A(n434), .B(n391), .Z(n102) );
  HS65_LH_BFX9 U280 ( .A(n197), .Z(n30) );
  HS65_LH_BFX9 U281 ( .A(n197), .Z(n31) );
  HS65_LH_BFX9 U282 ( .A(n26), .Z(n27) );
  HS65_LH_IVX9 U283 ( .A(n264), .Z(n573) );
  HS65_LH_AND2X4 U284 ( .A(n434), .B(n436), .Z(n103) );
  HS65_LH_BFX9 U285 ( .A(n26), .Z(n29) );
  HS65_LH_BFX9 U286 ( .A(n26), .Z(n28) );
  HS65_LH_BFX9 U287 ( .A(n199), .Z(n20) );
  HS65_LH_IVX9 U288 ( .A(n6), .Z(n18) );
  HS65_LH_BFX9 U289 ( .A(n537), .Z(n542) );
  HS65_LH_BFX9 U290 ( .A(n537), .Z(n541) );
  HS65_LH_BFX9 U291 ( .A(n536), .Z(n540) );
  HS65_LH_BFX9 U292 ( .A(n536), .Z(n539) );
  HS65_LH_BFX9 U293 ( .A(n536), .Z(n538) );
  HS65_LH_BFX9 U294 ( .A(n46), .Z(n49) );
  HS65_LH_BFX9 U295 ( .A(n537), .Z(n543) );
  HS65_LH_AO22X9 U296 ( .A(N167), .B(n63), .C(\HI_LO_c[LO][4] ), .D(n57), .Z(
        n457) );
  HS65_LH_AO22X9 U297 ( .A(N168), .B(n63), .C(\HI_LO_c[LO][5] ), .D(n57), .Z(
        n458) );
  HS65_LH_AO22X9 U298 ( .A(N169), .B(n62), .C(\HI_LO_c[LO][6] ), .D(n57), .Z(
        n459) );
  HS65_LH_AO22X9 U299 ( .A(N170), .B(n61), .C(\HI_LO_c[LO][7] ), .D(n57), .Z(
        n460) );
  HS65_LH_AO22X9 U300 ( .A(N171), .B(n66), .C(\HI_LO_c[LO][8] ), .D(n59), .Z(
        n461) );
  HS65_LH_AO22X9 U301 ( .A(N172), .B(n66), .C(\HI_LO_c[LO][9] ), .D(n58), .Z(
        n462) );
  HS65_LH_AO22X9 U302 ( .A(N173), .B(n65), .C(\HI_LO_c[LO][10] ), .D(n57), .Z(
        n463) );
  HS65_LH_AO22X9 U303 ( .A(N174), .B(n65), .C(\HI_LO_c[LO][11] ), .D(n60), .Z(
        n464) );
  HS65_LH_AO22X9 U304 ( .A(N175), .B(n65), .C(\HI_LO_c[LO][12] ), .D(n60), .Z(
        n465) );
  HS65_LH_AO22X9 U305 ( .A(N176), .B(n65), .C(\HI_LO_c[LO][13] ), .D(n60), .Z(
        n466) );
  HS65_LH_AO22X9 U306 ( .A(N177), .B(n65), .C(\HI_LO_c[LO][14] ), .D(n60), .Z(
        n467) );
  HS65_LH_AO22X9 U307 ( .A(N178), .B(n65), .C(\HI_LO_c[LO][15] ), .D(n60), .Z(
        n468) );
  HS65_LH_AO22X9 U308 ( .A(N199), .B(n64), .C(\HI_LO_c[HI][4] ), .D(n59), .Z(
        n489) );
  HS65_LH_AO22X9 U309 ( .A(N200), .B(n64), .C(\HI_LO_c[HI][5] ), .D(n59), .Z(
        n490) );
  HS65_LH_AO22X9 U310 ( .A(N201), .B(n64), .C(\HI_LO_c[HI][6] ), .D(n59), .Z(
        n491) );
  HS65_LH_AO22X9 U311 ( .A(N202), .B(n64), .C(\HI_LO_c[HI][7] ), .D(n59), .Z(
        n492) );
  HS65_LH_AO22X9 U312 ( .A(N203), .B(n64), .C(\HI_LO_c[HI][8] ), .D(n59), .Z(
        n493) );
  HS65_LH_AO22X9 U313 ( .A(N204), .B(n64), .C(\HI_LO_c[HI][9] ), .D(n59), .Z(
        n494) );
  HS65_LH_AO22X9 U314 ( .A(N205), .B(n64), .C(\HI_LO_c[HI][10] ), .D(n59), .Z(
        n495) );
  HS65_LH_AO22X9 U315 ( .A(N206), .B(n64), .C(\HI_LO_c[HI][11] ), .D(n59), .Z(
        n496) );
  HS65_LH_AO22X9 U316 ( .A(N207), .B(n64), .C(\HI_LO_c[HI][12] ), .D(n59), .Z(
        n497) );
  HS65_LH_AO22X9 U317 ( .A(N208), .B(n64), .C(\HI_LO_c[HI][13] ), .D(n59), .Z(
        n498) );
  HS65_LH_AO22X9 U318 ( .A(N209), .B(n64), .C(\HI_LO_c[HI][14] ), .D(n59), .Z(
        n499) );
  HS65_LH_AO22X9 U319 ( .A(N210), .B(n64), .C(\HI_LO_c[HI][15] ), .D(n59), .Z(
        n500) );
  HS65_LH_AO22X9 U320 ( .A(N211), .B(n64), .C(\HI_LO_c[HI][16] ), .D(n58), .Z(
        n501) );
  HS65_LH_AO22X9 U321 ( .A(N212), .B(n64), .C(\HI_LO_c[HI][17] ), .D(n58), .Z(
        n502) );
  HS65_LH_AO22X9 U322 ( .A(N213), .B(n63), .C(\HI_LO_c[HI][18] ), .D(n58), .Z(
        n503) );
  HS65_LH_AO22X9 U323 ( .A(N214), .B(n63), .C(\HI_LO_c[HI][19] ), .D(n58), .Z(
        n504) );
  HS65_LH_AO22X9 U324 ( .A(N215), .B(n63), .C(\HI_LO_c[HI][20] ), .D(n58), .Z(
        n505) );
  HS65_LH_AO22X9 U325 ( .A(N216), .B(n63), .C(\HI_LO_c[HI][21] ), .D(n58), .Z(
        n506) );
  HS65_LH_AO22X9 U326 ( .A(N217), .B(n63), .C(\HI_LO_c[HI][22] ), .D(n58), .Z(
        n507) );
  HS65_LH_AO22X9 U327 ( .A(N218), .B(n63), .C(\HI_LO_c[HI][23] ), .D(n58), .Z(
        n508) );
  HS65_LH_AO22X9 U328 ( .A(N219), .B(n63), .C(\HI_LO_c[HI][24] ), .D(n58), .Z(
        n509) );
  HS65_LH_AO22X9 U329 ( .A(N220), .B(n63), .C(\HI_LO_c[HI][25] ), .D(n58), .Z(
        n510) );
  HS65_LH_AO22X9 U330 ( .A(N221), .B(n63), .C(\HI_LO_c[HI][26] ), .D(n58), .Z(
        n511) );
  HS65_LH_AO22X9 U331 ( .A(N222), .B(n63), .C(\HI_LO_c[HI][27] ), .D(n58), .Z(
        n512) );
  HS65_LH_AO22X9 U332 ( .A(N226), .B(n63), .C(\HI_LO_c[HI][31] ), .D(n57), .Z(
        n516) );
  HS65_LH_AO22X9 U333 ( .A(N163), .B(n63), .C(\HI_LO_c[LO][0] ), .D(n57), .Z(
        n453) );
  HS65_LH_AO22X9 U334 ( .A(N164), .B(n63), .C(\HI_LO_c[LO][1] ), .D(n57), .Z(
        n454) );
  HS65_LH_AO22X9 U335 ( .A(N165), .B(n63), .C(\HI_LO_c[LO][2] ), .D(n57), .Z(
        n455) );
  HS65_LH_AO22X9 U336 ( .A(N166), .B(n63), .C(\HI_LO_c[LO][3] ), .D(n57), .Z(
        n456) );
  HS65_LH_AO22X9 U337 ( .A(N194), .B(n64), .C(\HI_LO_c[LO][31] ), .D(n59), .Z(
        n484) );
  HS65_LH_AO22X9 U338 ( .A(N196), .B(n64), .C(\HI_LO_c[HI][1] ), .D(n58), .Z(
        n486) );
  HS65_LH_AO22X9 U339 ( .A(N197), .B(n64), .C(\HI_LO_c[HI][2] ), .D(n57), .Z(
        n487) );
  HS65_LH_AO22X9 U340 ( .A(N198), .B(n64), .C(\HI_LO_c[HI][3] ), .D(n60), .Z(
        n488) );
  HS65_LH_AO22X9 U341 ( .A(N223), .B(n63), .C(\HI_LO_c[HI][28] ), .D(n57), .Z(
        n513) );
  HS65_LH_AO22X9 U342 ( .A(N224), .B(n63), .C(\HI_LO_c[HI][29] ), .D(n57), .Z(
        n514) );
  HS65_LH_AO22X9 U343 ( .A(N225), .B(n63), .C(\HI_LO_c[HI][30] ), .D(n57), .Z(
        n515) );
  HS65_LH_AO22X9 U344 ( .A(N179), .B(n65), .C(\HI_LO_c[LO][16] ), .D(n60), .Z(
        n469) );
  HS65_LH_AO22X9 U345 ( .A(N180), .B(n65), .C(\HI_LO_c[LO][17] ), .D(n60), .Z(
        n470) );
  HS65_LH_AO22X9 U346 ( .A(N181), .B(n65), .C(\HI_LO_c[LO][18] ), .D(n60), .Z(
        n471) );
  HS65_LH_AO22X9 U347 ( .A(N182), .B(n65), .C(\HI_LO_c[LO][19] ), .D(n60), .Z(
        n472) );
  HS65_LH_AO22X9 U348 ( .A(N183), .B(n65), .C(\HI_LO_c[LO][20] ), .D(n60), .Z(
        n473) );
  HS65_LH_AO22X9 U349 ( .A(N184), .B(n65), .C(\HI_LO_c[LO][21] ), .D(n60), .Z(
        n474) );
  HS65_LH_AO22X9 U350 ( .A(N185), .B(n65), .C(\HI_LO_c[LO][22] ), .D(n60), .Z(
        n475) );
  HS65_LH_AO22X9 U351 ( .A(N186), .B(n65), .C(\HI_LO_c[LO][23] ), .D(n60), .Z(
        n476) );
  HS65_LH_AO22X9 U352 ( .A(N187), .B(n65), .C(\HI_LO_c[LO][24] ), .D(n59), .Z(
        n477) );
  HS65_LH_AO22X9 U353 ( .A(N188), .B(n65), .C(\HI_LO_c[LO][25] ), .D(n58), .Z(
        n478) );
  HS65_LH_AO22X9 U354 ( .A(N189), .B(n65), .C(\HI_LO_c[LO][26] ), .D(n57), .Z(
        n479) );
  HS65_LH_AO22X9 U355 ( .A(N190), .B(n65), .C(\HI_LO_c[LO][27] ), .D(n60), .Z(
        n480) );
  HS65_LH_AO22X9 U356 ( .A(N191), .B(n65), .C(\HI_LO_c[LO][28] ), .D(n59), .Z(
        n481) );
  HS65_LH_AO22X9 U357 ( .A(N192), .B(n65), .C(\HI_LO_c[LO][29] ), .D(n58), .Z(
        n482) );
  HS65_LH_AO22X9 U358 ( .A(N193), .B(n64), .C(\HI_LO_c[LO][30] ), .D(n57), .Z(
        n483) );
  HS65_LH_AO22X9 U359 ( .A(N195), .B(n64), .C(\HI_LO_c[HI][0] ), .D(n60), .Z(
        n485) );
  HS65_LH_NOR4ABX4 U360 ( .A(n578), .B(n435), .C(\alu_i[OP][3] ), .D(
        \alu_i[OP][2] ), .Z(n180) );
  HS65_LH_NOR3X4 U361 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][4] ), .C(n587), .Z(
        n434) );
  HS65_LH_AND2X4 U362 ( .A(\alu_i[SHAMT][1] ), .B(\alu_i[SHAMT][0] ), .Z(n199)
         );
  HS65_LH_AOI222X2 U363 ( .A(n317), .B(n17), .C(n316), .D(n7), .E(n178), .F(
        \alu_i[SHAMT][3] ), .Z(n264) );
  HS65_LH_AOI222X2 U364 ( .A(n144), .B(n17), .C(n325), .D(n8), .E(n283), .F(
        \alu_i[SHAMT][3] ), .Z(n190) );
  HS65_LH_NOR2X6 U365 ( .A(n594), .B(\alu_i[SHAMT][3] ), .Z(n7) );
  HS65_LH_NOR2X6 U366 ( .A(n594), .B(\alu_i[SHAMT][3] ), .Z(n8) );
  HS65_LH_AOI222X2 U367 ( .A(n44), .B(\HI_LO_c[LO][4] ), .C(n579), .D(n173), 
        .E(N103), .F(n47), .Z(n172) );
  HS65_LH_AOI222X2 U368 ( .A(n44), .B(\HI_LO_c[LO][5] ), .C(n579), .D(n164), 
        .E(N104), .F(n47), .Z(n163) );
  HS65_LH_AOI222X2 U369 ( .A(n44), .B(\HI_LO_c[LO][6] ), .C(n579), .D(n152), 
        .E(N105), .F(n47), .Z(n151) );
  HS65_LH_AOI222X2 U370 ( .A(n44), .B(\HI_LO_c[LO][7] ), .C(n579), .D(n140), 
        .E(N106), .F(n47), .Z(n139) );
  HS65_LH_AOI222X2 U371 ( .A(n44), .B(\HI_LO_c[LO][8] ), .C(n579), .D(n128), 
        .E(N107), .F(n47), .Z(n127) );
  HS65_LH_AOI222X2 U372 ( .A(n44), .B(\HI_LO_c[LO][9] ), .C(n579), .D(n111), 
        .E(N108), .F(n47), .Z(n110) );
  HS65_LH_AOI222X2 U373 ( .A(n44), .B(\HI_LO_c[LO][10] ), .C(n579), .D(n154), 
        .E(N109), .F(n47), .Z(n427) );
  HS65_LH_AOI222X2 U374 ( .A(n44), .B(\HI_LO_c[LO][11] ), .C(n579), .D(n142), 
        .E(N110), .F(n47), .Z(n420) );
  HS65_LH_AOI222X2 U375 ( .A(n44), .B(\HI_LO_c[LO][12] ), .C(n579), .D(n130), 
        .E(N111), .F(n47), .Z(n414) );
  HS65_LH_AOI222X2 U376 ( .A(n44), .B(\HI_LO_c[LO][13] ), .C(n579), .D(n114), 
        .E(N112), .F(n47), .Z(n408) );
  HS65_LH_AOI222X2 U377 ( .A(n44), .B(\HI_LO_c[LO][14] ), .C(n579), .D(n157), 
        .E(N113), .F(n47), .Z(n402) );
  HS65_LH_AOI222X2 U378 ( .A(n44), .B(\HI_LO_c[LO][15] ), .C(n579), .D(n145), 
        .E(N114), .F(n47), .Z(n395) );
  HS65_LH_NOR2AX3 U379 ( .A(\alu_i[SHAMT][0] ), .B(\alu_i[SHAMT][1] ), .Z(n197) );
  HS65_LH_AOI212X4 U380 ( .A(\alu_i[SRC_A][4] ), .B(n180), .C(n56), .D(n562), 
        .E(n42), .Z(n175) );
  HS65_LH_IVX9 U381 ( .A(\alu_i[SRC_A][4] ), .Z(n562) );
  HS65_LH_AOI212X4 U382 ( .A(\alu_i[SRC_A][27] ), .B(n180), .C(n56), .D(n547), 
        .E(n42), .Z(n280) );
  HS65_LH_IVX9 U383 ( .A(\alu_i[SRC_A][27] ), .Z(n547) );
  HS65_LH_NOR2X6 U384 ( .A(n96), .B(\alu_i[SHAMT][4] ), .Z(n113) );
  HS65_LH_NOR2X6 U385 ( .A(n594), .B(\alu_i[SHAMT][3] ), .Z(n301) );
  HS65_LH_IVX9 U386 ( .A(\alu_i[SHAMT][3] ), .Z(n593) );
  HS65_LH_NOR2X6 U387 ( .A(n593), .B(\alu_i[SHAMT][2] ), .Z(n304) );
  HS65_LH_OAI212X5 U388 ( .A(n185), .B(n72), .C(n575), .D(n186), .E(n187), .Z(
        n184) );
  HS65_LH_IVX9 U389 ( .A(n188), .Z(n575) );
  HS65_LH_CBI4I1X5 U390 ( .A(n56), .B(n72), .C(n42), .D(\alu_i[SRC_A][3] ), 
        .Z(n187) );
  HS65_LH_AOI212X4 U391 ( .A(\alu_i[SRC_A][3] ), .B(n180), .C(n56), .D(n563), 
        .E(n42), .Z(n185) );
  HS65_LH_OAI212X5 U392 ( .A(n261), .B(n522), .C(n567), .D(n208), .E(n262), 
        .Z(n260) );
  HS65_LH_IVX9 U393 ( .A(n263), .Z(n567) );
  HS65_LH_CBI4I1X5 U394 ( .A(n56), .B(n522), .C(n42), .D(\alu_i[SRC_A][28] ), 
        .Z(n262) );
  HS65_LH_AOI212X4 U395 ( .A(\alu_i[SRC_A][28] ), .B(n180), .C(n56), .D(n546), 
        .E(n42), .Z(n261) );
  HS65_LH_OAI212X5 U396 ( .A(\alu_i[SRC_A][0] ), .B(n55), .C(n9), .D(n565), 
        .E(n441), .Z(n439) );
  HS65_LH_AOI12X2 U397 ( .A(n583), .B(n196), .C(n42), .Z(n441) );
  HS65_LH_OAI212X5 U398 ( .A(\alu_i[SRC_A][30] ), .B(n55), .C(n9), .D(n545), 
        .E(n41), .Z(n223) );
  HS65_LH_OAI212X5 U399 ( .A(\alu_i[SRC_A][1] ), .B(n97), .C(n10), .D(n564), 
        .E(n41), .Z(n357) );
  HS65_LH_NOR2X6 U400 ( .A(n6), .B(\alu_i[SHAMT][4] ), .Z(n193) );
  HS65_LH_OAI212X5 U401 ( .A(\alu_i[SRC_A][12] ), .B(n54), .C(n10), .D(n557), 
        .E(n123), .Z(n415) );
  HS65_LH_IVX9 U402 ( .A(\alu_i[SRC_A][12] ), .Z(n557) );
  HS65_LH_OAI212X5 U403 ( .A(\alu_i[SRC_A][13] ), .B(n97), .C(n10), .D(n556), 
        .E(n40), .Z(n409) );
  HS65_LH_IVX9 U404 ( .A(\alu_i[SRC_A][13] ), .Z(n556) );
  HS65_LH_OAI212X5 U405 ( .A(\alu_i[SRC_A][15] ), .B(n54), .C(n10), .D(n555), 
        .E(n123), .Z(n396) );
  HS65_LH_IVX9 U406 ( .A(\alu_i[SRC_A][15] ), .Z(n555) );
  HS65_LH_OAI212X5 U407 ( .A(\alu_i[SRC_A][16] ), .B(n97), .C(n10), .D(n554), 
        .E(n41), .Z(n388) );
  HS65_LH_IVX9 U408 ( .A(\alu_i[SRC_A][16] ), .Z(n554) );
  HS65_LH_OAI212X5 U409 ( .A(\alu_i[SRC_A][18] ), .B(n54), .C(n10), .D(n553), 
        .E(n40), .Z(n375) );
  HS65_LH_IVX9 U410 ( .A(\alu_i[SRC_A][18] ), .Z(n553) );
  HS65_LH_OAI212X5 U411 ( .A(\alu_i[SRC_A][19] ), .B(n97), .C(n10), .D(n552), 
        .E(n123), .Z(n367) );
  HS65_LH_IVX9 U412 ( .A(\alu_i[SRC_A][19] ), .Z(n552) );
  HS65_LH_OAI212X5 U413 ( .A(\alu_i[SRC_A][6] ), .B(n55), .C(n9), .D(n561), 
        .E(n41), .Z(n158) );
  HS65_LH_IVX9 U414 ( .A(\alu_i[SRC_A][6] ), .Z(n561) );
  HS65_LH_OAI212X5 U415 ( .A(\alu_i[SRC_A][7] ), .B(n55), .C(n9), .D(n560), 
        .E(n41), .Z(n146) );
  HS65_LH_IVX9 U416 ( .A(\alu_i[SRC_A][7] ), .Z(n560) );
  HS65_LH_OAI212X5 U417 ( .A(\alu_i[SRC_A][9] ), .B(n55), .C(n559), .D(n10), 
        .E(n123), .Z(n121) );
  HS65_LH_IVX9 U418 ( .A(\alu_i[SRC_A][9] ), .Z(n559) );
  HS65_LH_OAI212X5 U419 ( .A(\alu_i[SRC_A][24] ), .B(n55), .C(n9), .D(n549), 
        .E(n41), .Z(n318) );
  HS65_LH_IVX9 U420 ( .A(\alu_i[SRC_A][24] ), .Z(n549) );
  HS65_LH_AOI32X5 U421 ( .A(n283), .B(n593), .C(n284), .D(\alu_i[SRC_A][27] ), 
        .E(n285), .Z(n282) );
  HS65_LH_OAI21X3 U422 ( .A(\alu_i[SRC_B][27] ), .B(n54), .C(n123), .Z(n285)
         );
  HS65_LH_OAI212X5 U423 ( .A(\alu_i[SRC_A][10] ), .B(n54), .C(n10), .D(n558), 
        .E(n41), .Z(n428) );
  HS65_LH_IVX9 U424 ( .A(\alu_i[SRC_A][10] ), .Z(n558) );
  HS65_LH_OAI212X5 U425 ( .A(\alu_i[SRC_A][21] ), .B(n97), .C(n10), .D(n551), 
        .E(n41), .Z(n344) );
  HS65_LH_IVX9 U426 ( .A(\alu_i[SRC_A][21] ), .Z(n551) );
  HS65_LH_OAI212X5 U427 ( .A(\alu_i[SRC_A][22] ), .B(n54), .C(n9), .D(n550), 
        .E(n41), .Z(n338) );
  HS65_LH_IVX9 U428 ( .A(\alu_i[SRC_A][22] ), .Z(n550) );
  HS65_LH_OAI212X5 U429 ( .A(\alu_i[SRC_A][25] ), .B(n97), .C(n9), .D(n548), 
        .E(n41), .Z(n307) );
  HS65_LH_IVX9 U430 ( .A(\alu_i[SRC_A][25] ), .Z(n548) );
  HS65_LH_AOI32X5 U431 ( .A(n178), .B(n593), .C(n113), .D(\alu_i[SRC_A][4] ), 
        .E(n179), .Z(n177) );
  HS65_LH_OAI21X3 U432 ( .A(\alu_i[SRC_B][4] ), .B(n97), .C(n40), .Z(n179) );
  HS65_LH_NOR2X6 U433 ( .A(n590), .B(\alu_i[OP][1] ), .Z(n391) );
  HS65_LH_IVX9 U434 ( .A(\alu_i[SHAMT][4] ), .Z(n592) );
  HS65_LH_IVX9 U435 ( .A(\alu_i[SHAMT][2] ), .Z(n594) );
  HS65_LH_NOR2X6 U436 ( .A(\alu_i[OP][1] ), .B(\alu_i[OP][0] ), .Z(n438) );
  HS65_LH_NOR2X6 U437 ( .A(n588), .B(\alu_i[OP][0] ), .Z(n436) );
  HS65_LH_NOR2X6 U438 ( .A(n593), .B(\alu_i[SHAMT][4] ), .Z(n448) );
  HS65_LH_NAND4ABX3 U439 ( .A(\alu_i[OP][4] ), .B(\alu_i[OP][2] ), .C(n588), 
        .D(n587), .Z(n437) );
  HS65_LH_AND2X4 U440 ( .A(n448), .B(\alu_i[SHAMT][2] ), .Z(n192) );
  HS65_LH_AO22X9 U441 ( .A(n594), .B(n314), .C(\alu_i[SHAMT][2] ), .D(n315), 
        .Z(n178) );
  HS65_LH_AO22X9 U442 ( .A(n594), .B(n324), .C(\alu_i[SHAMT][2] ), .D(n216), 
        .Z(n283) );
  HS65_LH_OAI21X3 U443 ( .A(n205), .B(n525), .C(n206), .Z(n204) );
  HS65_LH_CBI4I1X5 U444 ( .A(n56), .B(n525), .C(n42), .D(\alu_i[SRC_A][31] ), 
        .Z(n206) );
  HS65_LH_AOI212X4 U445 ( .A(n56), .B(n544), .C(\alu_i[SRC_A][31] ), .D(n180), 
        .E(n207), .Z(n205) );
  HS65_LH_IVX9 U446 ( .A(\alu_i[SRC_A][31] ), .Z(n544) );
  HS65_LH_AND2X4 U447 ( .A(n445), .B(\alu_i[OP][3] ), .Z(n390) );
  HS65_LH_NOR2AX3 U448 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][4] ), .Z(n445) );
  HS65_LH_NAND4ABX3 U449 ( .A(n383), .B(n384), .C(n385), .D(n386), .Z(
        \alu_o[RESULT][16] ) );
  HS65_LH_MX41X7 U450 ( .D0(n582), .S0(n316), .D1(n85), .S1(n388), .D2(n368), 
        .S2(n315), .D3(\alu_i[SRC_A][16] ), .S3(n389), .Z(n384) );
  HS65_LH_MX41X7 U451 ( .D0(n45), .S0(\HI_LO_c[LO][16] ), .D1(n106), .S1(n69), 
        .D2(N115), .S2(n49), .D3(n583), .S3(n266), .Z(n383) );
  HS65_LH_AOI222X2 U452 ( .A(N147), .B(n52), .C(n15), .D(\HI_LO_c[HI][16] ), 
        .E(n12), .F(n86), .Z(n385) );
  HS65_LH_NAND4ABX3 U453 ( .A(n377), .B(n378), .C(n379), .D(n380), .Z(
        \alu_o[RESULT][17] ) );
  HS65_LH_MX41X7 U454 ( .D0(n582), .S0(n305), .D1(n86), .S1(n381), .D2(n368), 
        .S2(n303), .D3(\alu_i[SRC_A][17] ), .S3(n382), .Z(n378) );
  HS65_LH_MX41X7 U455 ( .D0(n45), .S0(\HI_LO_c[LO][17] ), .D1(n106), .S1(n70), 
        .D2(N116), .S2(n49), .D3(n583), .S3(n254), .Z(n377) );
  HS65_LH_AOI222X2 U456 ( .A(N148), .B(n52), .C(n15), .D(\HI_LO_c[HI][17] ), 
        .E(n12), .F(n87), .Z(n379) );
  HS65_LH_NAND4ABX3 U457 ( .A(n370), .B(n371), .C(n372), .D(n373), .Z(
        \alu_o[RESULT][18] ) );
  HS65_LH_MX41X7 U458 ( .D0(n582), .S0(n337), .D1(n87), .S1(n375), .D2(n368), 
        .S2(n576), .D3(\alu_i[SRC_A][18] ), .S3(n376), .Z(n371) );
  HS65_LH_MX41X7 U459 ( .D0(n45), .S0(\HI_LO_c[LO][18] ), .D1(n106), .S1(
        \alu_i[SRC_B][2] ), .D2(N117), .S2(n49), .D3(n583), .S3(n229), .Z(n370) );
  HS65_LH_AOI222X2 U460 ( .A(N149), .B(n52), .C(n15), .D(\HI_LO_c[HI][18] ), 
        .E(n12), .F(n88), .Z(n372) );
  HS65_LH_NAND4ABX3 U461 ( .A(n363), .B(n364), .C(n365), .D(n366), .Z(
        \alu_o[RESULT][19] ) );
  HS65_LH_MX41X7 U462 ( .D0(n582), .S0(n327), .D1(n88), .S1(n367), .D2(n368), 
        .S2(n188), .D3(\alu_i[SRC_A][19] ), .S3(n369), .Z(n364) );
  HS65_LH_MX41X7 U463 ( .D0(n45), .S0(\HI_LO_c[LO][19] ), .D1(n106), .S1(
        \alu_i[SRC_B][3] ), .D2(N118), .S2(n48), .D3(n583), .S3(n212), .Z(n363) );
  HS65_LH_AOI222X2 U464 ( .A(N150), .B(n52), .C(n15), .D(\HI_LO_c[HI][19] ), 
        .E(n12), .F(\alu_i[SRC_B][20] ), .Z(n365) );
  HS65_LH_NAND4ABX3 U465 ( .A(n346), .B(n347), .C(n348), .D(n349), .Z(
        \alu_o[RESULT][20] ) );
  HS65_LH_MX41X7 U466 ( .D0(n45), .S0(\HI_LO_c[LO][20] ), .D1(n106), .S1(
        \alu_i[SRC_B][4] ), .D2(N119), .S2(n48), .D3(n583), .S3(n268), .Z(n346) );
  HS65_LH_OAI212X5 U467 ( .A(n350), .B(n89), .C(n572), .D(n281), .E(n351), .Z(
        n347) );
  HS65_LH_AOI222X2 U468 ( .A(N151), .B(n52), .C(n15), .D(\HI_LO_c[HI][20] ), 
        .E(n12), .F(n90), .Z(n348) );
  HS65_LH_NAND4ABX3 U469 ( .A(n271), .B(n272), .C(n273), .D(n274), .Z(
        \alu_o[RESULT][27] ) );
  HS65_LH_MX41X7 U470 ( .D0(n45), .S0(\HI_LO_c[LO][27] ), .D1(n106), .S1(
        \alu_i[SRC_B][11] ), .D2(N126), .S2(n48), .D3(n583), .S3(n209), .Z(
        n271) );
  HS65_LH_OAI212X5 U471 ( .A(n280), .B(n521), .C(n570), .D(n281), .E(n282), 
        .Z(n272) );
  HS65_LH_AOI222X2 U472 ( .A(N158), .B(n51), .C(n14), .D(\HI_LO_c[HI][27] ), 
        .E(n11), .F(\alu_i[SRC_B][28] ), .Z(n273) );
  HS65_LH_NAND4ABX3 U473 ( .A(n340), .B(n341), .C(n342), .D(n343), .Z(
        \alu_o[RESULT][21] ) );
  HS65_LH_MX41X7 U474 ( .D0(n277), .S0(n305), .D1(n582), .S1(n306), .D2(n90), 
        .S2(n344), .D3(\alu_i[SRC_A][21] ), .S3(n345), .Z(n341) );
  HS65_LH_MX41X7 U475 ( .D0(n45), .S0(\HI_LO_c[LO][21] ), .D1(n106), .S1(n74), 
        .D2(N120), .S2(n48), .D3(n583), .S3(n256), .Z(n340) );
  HS65_LH_AOI222X2 U476 ( .A(N152), .B(n52), .C(n14), .D(\HI_LO_c[HI][21] ), 
        .E(n11), .F(n300), .Z(n342) );
  HS65_LH_NAND4ABX3 U477 ( .A(n330), .B(n331), .C(n332), .D(n333), .Z(
        \alu_o[RESULT][22] ) );
  HS65_LH_MX41X7 U478 ( .D0(n277), .S0(n337), .D1(n582), .S1(n292), .D2(n300), 
        .S2(n338), .D3(\alu_i[SRC_A][22] ), .S3(n339), .Z(n331) );
  HS65_LH_MX41X7 U479 ( .D0(n45), .S0(\HI_LO_c[LO][22] ), .D1(n106), .S1(n75), 
        .D2(N121), .S2(n48), .D3(n583), .S3(n231), .Z(n330) );
  HS65_LH_AOI222X2 U480 ( .A(N153), .B(n51), .C(n14), .D(\HI_LO_c[HI][22] ), 
        .E(n11), .F(n517), .Z(n332) );
  HS65_LH_NAND4ABX3 U481 ( .A(n320), .B(n321), .C(n322), .D(n323), .Z(
        \alu_o[RESULT][23] ) );
  HS65_LH_MX41X7 U482 ( .D0(n277), .S0(n327), .D1(n582), .S1(n278), .D2(n517), 
        .S2(n328), .D3(\alu_i[SRC_A][23] ), .S3(n329), .Z(n321) );
  HS65_LH_MX41X7 U483 ( .D0(n45), .S0(\HI_LO_c[LO][23] ), .D1(n106), .S1(n76), 
        .D2(N122), .S2(n48), .D3(n583), .S3(n214), .Z(n320) );
  HS65_LH_AOI222X2 U484 ( .A(N154), .B(n51), .C(n14), .D(\HI_LO_c[HI][23] ), 
        .E(n11), .F(n518), .Z(n322) );
  HS65_LH_NAND4ABX3 U485 ( .A(n309), .B(n310), .C(n311), .D(n312), .Z(
        \alu_o[RESULT][24] ) );
  HS65_LH_MX41X7 U486 ( .D0(n277), .S0(n317), .D1(n582), .S1(n266), .D2(n518), 
        .S2(n318), .D3(\alu_i[SRC_A][24] ), .S3(n319), .Z(n310) );
  HS65_LH_MX41X7 U487 ( .D0(n45), .S0(\HI_LO_c[LO][24] ), .D1(n106), .S1(n77), 
        .D2(N123), .S2(n48), .D3(n583), .S3(n269), .Z(n309) );
  HS65_LH_AOI222X2 U488 ( .A(N155), .B(n51), .C(n14), .D(\HI_LO_c[HI][24] ), 
        .E(n11), .F(n519), .Z(n311) );
  HS65_LH_NAND4ABX3 U489 ( .A(n295), .B(n296), .C(n297), .D(n298), .Z(
        \alu_o[RESULT][25] ) );
  HS65_LH_MX41X7 U490 ( .D0(n277), .S0(n306), .D1(n582), .S1(n254), .D2(n519), 
        .S2(n307), .D3(\alu_i[SRC_A][25] ), .S3(n308), .Z(n296) );
  HS65_LH_MX41X7 U491 ( .D0(n45), .S0(\HI_LO_c[LO][25] ), .D1(n106), .S1(n78), 
        .D2(N124), .S2(n48), .D3(n583), .S3(n251), .Z(n295) );
  HS65_LH_AOI222X2 U492 ( .A(N156), .B(n51), .C(n14), .D(\HI_LO_c[HI][25] ), 
        .E(n11), .F(n520), .Z(n297) );
  HS65_LH_NAND4ABX3 U493 ( .A(n286), .B(n287), .C(n288), .D(n289), .Z(
        \alu_o[RESULT][26] ) );
  HS65_LH_MX41X7 U494 ( .D0(n277), .S0(n292), .D1(n582), .S1(n229), .D2(n520), 
        .S2(n293), .D3(\alu_i[SRC_A][26] ), .S3(n294), .Z(n287) );
  HS65_LH_MX41X7 U495 ( .D0(n45), .S0(\HI_LO_c[LO][26] ), .D1(n106), .S1(n79), 
        .D2(N125), .S2(n48), .D3(n583), .S3(n226), .Z(n286) );
  HS65_LH_AOI222X2 U496 ( .A(N157), .B(n51), .C(n14), .D(\HI_LO_c[HI][26] ), 
        .E(n11), .F(\alu_i[SRC_B][27] ), .Z(n288) );
  HS65_LH_NAND4ABX3 U497 ( .A(n169), .B(n170), .C(n171), .D(n172), .Z(
        \alu_o[RESULT][4] ) );
  HS65_LH_AO222X4 U498 ( .A(n128), .B(n115), .C(n133), .D(n118), .E(n174), .F(
        n117), .Z(n170) );
  HS65_LH_OAI212X5 U499 ( .A(n175), .B(n73), .C(n571), .D(n176), .E(n177), .Z(
        n169) );
  HS65_LH_AOI222X2 U500 ( .A(N135), .B(n51), .C(n14), .D(\HI_LO_c[HI][4] ), 
        .E(n11), .F(n74), .Z(n171) );
  HS65_LH_NAND4ABX3 U501 ( .A(n160), .B(n161), .C(n162), .D(n163), .Z(
        \alu_o[RESULT][5] ) );
  HS65_LH_MX41X7 U502 ( .D0(n118), .S0(n120), .D1(n580), .S1(n114), .D2(n74), 
        .S2(n167), .D3(\alu_i[SRC_A][5] ), .S3(n168), .Z(n160) );
  HS65_LH_AO222X4 U503 ( .A(n165), .B(n113), .C(n111), .D(n115), .E(n166), .F(
        n117), .Z(n161) );
  HS65_LH_AOI222X2 U504 ( .A(N136), .B(n51), .C(n15), .D(\HI_LO_c[HI][5] ), 
        .E(n11), .F(n75), .Z(n162) );
  HS65_LH_NAND4ABX3 U505 ( .A(n148), .B(n149), .C(n150), .D(n151), .Z(
        \alu_o[RESULT][6] ) );
  HS65_LH_MX41X7 U506 ( .D0(n118), .S0(n156), .D1(n580), .S1(n157), .D2(n75), 
        .S2(n158), .D3(\alu_i[SRC_A][6] ), .S3(n159), .Z(n148) );
  HS65_LH_AO222X4 U507 ( .A(n153), .B(n113), .C(n154), .D(n115), .E(n155), .F(
        n117), .Z(n149) );
  HS65_LH_AOI222X2 U508 ( .A(N137), .B(n51), .C(n14), .D(\HI_LO_c[HI][6] ), 
        .E(n11), .F(n76), .Z(n150) );
  HS65_LH_NAND4ABX3 U509 ( .A(n136), .B(n137), .C(n138), .D(n139), .Z(
        \alu_o[RESULT][7] ) );
  HS65_LH_MX41X7 U510 ( .D0(n118), .S0(n144), .D1(n580), .S1(n145), .D2(n76), 
        .S2(n146), .D3(\alu_i[SRC_A][7] ), .S3(n147), .Z(n136) );
  HS65_LH_AO222X4 U511 ( .A(n141), .B(n113), .C(n142), .D(n115), .E(n143), .F(
        n117), .Z(n137) );
  HS65_LH_AOI222X2 U512 ( .A(N138), .B(n51), .C(n14), .D(\HI_LO_c[HI][7] ), 
        .E(n11), .F(n77), .Z(n138) );
  HS65_LH_NAND4ABX3 U513 ( .A(n124), .B(n125), .C(n126), .D(n127), .Z(
        \alu_o[RESULT][8] ) );
  HS65_LH_MX41X7 U514 ( .D0(n118), .S0(n132), .D1(n580), .S1(n133), .D2(n77), 
        .S2(n134), .D3(\alu_i[SRC_A][8] ), .S3(n135), .Z(n124) );
  HS65_LH_AO222X4 U515 ( .A(n129), .B(n113), .C(n130), .D(n115), .E(n131), .F(
        n117), .Z(n125) );
  HS65_LH_AOI222X2 U516 ( .A(N139), .B(n51), .C(n14), .D(\HI_LO_c[HI][8] ), 
        .E(n11), .F(n78), .Z(n126) );
  HS65_LH_NAND4ABX3 U517 ( .A(n107), .B(n108), .C(n109), .D(n110), .Z(
        \alu_o[RESULT][9] ) );
  HS65_LH_MX41X7 U518 ( .D0(n118), .S0(n119), .D1(n580), .S1(n120), .D2(n78), 
        .S2(n121), .D3(\alu_i[SRC_A][9] ), .S3(n122), .Z(n107) );
  HS65_LH_AO222X4 U519 ( .A(n112), .B(n113), .C(n114), .D(n115), .E(n116), .F(
        n117), .Z(n108) );
  HS65_LH_AOI222X2 U520 ( .A(N140), .B(n51), .C(n14), .D(\HI_LO_c[HI][9] ), 
        .E(n11), .F(n79), .Z(n109) );
  HS65_LH_NAND4ABX3 U521 ( .A(n424), .B(n425), .C(n426), .D(n427), .Z(
        \alu_o[RESULT][10] ) );
  HS65_LH_MX41X7 U522 ( .D0(n118), .S0(n335), .D1(n580), .S1(n156), .D2(n79), 
        .S2(n428), .D3(\alu_i[SRC_A][10] ), .S3(n429), .Z(n424) );
  HS65_LH_AO222X4 U523 ( .A(n290), .B(n113), .C(n157), .D(n115), .E(n291), .F(
        n117), .Z(n425) );
  HS65_LH_AOI222X2 U524 ( .A(N141), .B(n52), .C(n15), .D(\HI_LO_c[HI][10] ), 
        .E(n12), .F(\alu_i[SRC_B][11] ), .Z(n426) );
  HS65_LH_NAND4ABX3 U525 ( .A(n417), .B(n418), .C(n419), .D(n420), .Z(
        \alu_o[RESULT][11] ) );
  HS65_LH_AO222X4 U526 ( .A(n145), .B(n115), .C(n325), .D(n118), .E(n276), .F(
        n113), .Z(n418) );
  HS65_LH_OAI212X5 U527 ( .A(n421), .B(n80), .C(n569), .D(n176), .E(n422), .Z(
        n417) );
  HS65_LH_AOI222X2 U528 ( .A(N142), .B(n52), .C(n15), .D(\HI_LO_c[HI][11] ), 
        .E(n12), .F(n81), .Z(n419) );
  HS65_LH_NAND4ABX3 U529 ( .A(n411), .B(n412), .C(n413), .D(n414), .Z(
        \alu_o[RESULT][12] ) );
  HS65_LH_MX41X7 U530 ( .D0(n580), .S0(n132), .D1(n81), .S1(n415), .D2(n397), 
        .S2(n263), .D3(\alu_i[SRC_A][12] ), .S3(n416), .Z(n411) );
  HS65_LH_AO222X4 U531 ( .A(n133), .B(n115), .C(n313), .D(n118), .E(n573), .F(
        n113), .Z(n412) );
  HS65_LH_AOI222X2 U532 ( .A(N143), .B(n52), .C(n15), .D(\HI_LO_c[HI][12] ), 
        .E(n12), .F(n82), .Z(n413) );
  HS65_LH_NAND4ABX3 U533 ( .A(n405), .B(n406), .C(n407), .D(n408), .Z(
        \alu_o[RESULT][13] ) );
  HS65_LH_MX41X7 U534 ( .D0(n580), .S0(n119), .D1(n82), .S1(n409), .D2(n397), 
        .S2(n247), .D3(\alu_i[SRC_A][13] ), .S3(n410), .Z(n405) );
  HS65_LH_AO222X4 U535 ( .A(n120), .B(n115), .C(n299), .D(n118), .E(n252), .F(
        n113), .Z(n406) );
  HS65_LH_AOI222X2 U536 ( .A(N144), .B(n52), .C(n15), .D(\HI_LO_c[HI][13] ), 
        .E(n12), .F(n83), .Z(n407) );
  HS65_LH_NAND4ABX3 U537 ( .A(n399), .B(n400), .C(n401), .D(n402), .Z(
        \alu_o[RESULT][14] ) );
  HS65_LH_MX41X7 U538 ( .D0(n580), .S0(n335), .D1(n83), .S1(n403), .D2(n397), 
        .S2(n222), .D3(\alu_i[SRC_A][14] ), .S3(n404), .Z(n399) );
  HS65_LH_AO222X4 U539 ( .A(n156), .B(n115), .C(n334), .D(n118), .E(n227), .F(
        n113), .Z(n400) );
  HS65_LH_AOI222X2 U540 ( .A(N145), .B(n52), .C(n15), .D(\HI_LO_c[HI][14] ), 
        .E(n12), .F(n84), .Z(n401) );
  HS65_LH_NAND4ABX3 U541 ( .A(n392), .B(n393), .C(n394), .D(n395), .Z(
        \alu_o[RESULT][15] ) );
  HS65_LH_MX41X7 U542 ( .D0(n580), .S0(n325), .D1(n84), .S1(n396), .D2(n397), 
        .S2(n216), .D3(\alu_i[SRC_A][15] ), .S3(n398), .Z(n392) );
  HS65_LH_AO222X4 U543 ( .A(n144), .B(n115), .C(n324), .D(n118), .E(n210), .F(
        n113), .Z(n393) );
  HS65_LH_AOI222X2 U544 ( .A(N146), .B(n52), .C(n15), .D(\HI_LO_c[HI][15] ), 
        .E(n12), .F(n85), .Z(n394) );
  HS65_LH_AO222X4 U545 ( .A(N649), .B(n103), .C(n16), .D(\HI_LO_c[HI][0] ), 
        .E(N648), .F(n102), .Z(n433) );
  HS65_LH_AO222X4 U546 ( .A(\HI_LO_c[LO][29] ), .B(n45), .C(n82), .D(n106), 
        .E(\HI_LO_c[HI][29] ), .F(n16), .Z(n246) );
  HS65_LH_AO222X4 U547 ( .A(\HI_LO_c[LO][30] ), .B(n105), .C(n83), .D(n106), 
        .E(\HI_LO_c[HI][30] ), .F(n16), .Z(n221) );
  HS65_LH_IVX9 U548 ( .A(\alu_i[OP][4] ), .Z(n578) );
  HS65_LH_AO212X4 U549 ( .A(n173), .B(n591), .C(n387), .D(\alu_i[SHAMT][4] ), 
        .E(n446), .Z(n444) );
  HS65_LH_AO222X4 U550 ( .A(n192), .B(n130), .C(n193), .D(n447), .E(n195), .F(
        n128), .Z(n446) );
  HS65_LH_AO212X4 U551 ( .A(n27), .B(\alu_i[SRC_B][2] ), .C(n35), .D(n70), .E(
        n449), .Z(n447) );
  HS65_LH_AO12X9 U552 ( .A(\alu_i[SRC_B][3] ), .B(n21), .C(n315), .Z(n449) );
  HS65_LH_AO212X4 U553 ( .A(n164), .B(n591), .C(n360), .D(\alu_i[SHAMT][4] ), 
        .E(n361), .Z(n359) );
  HS65_LH_AO222X4 U554 ( .A(n192), .B(n114), .C(n193), .D(n362), .E(n195), .F(
        n111), .Z(n361) );
  HS65_LH_MX41X7 U555 ( .D0(n70), .S0(n37), .D1(\alu_i[SRC_B][2] ), .S1(n33), 
        .D2(\alu_i[SRC_B][3] ), .S2(n28), .D3(\alu_i[SRC_B][4] ), .S3(n22), 
        .Z(n362) );
  HS65_LH_AO212X4 U556 ( .A(n251), .B(n591), .C(n252), .D(\alu_i[SHAMT][4] ), 
        .E(n253), .Z(n250) );
  HS65_LH_AO222X4 U557 ( .A(n192), .B(n254), .C(n193), .D(n255), .E(n195), .F(
        n256), .Z(n253) );
  HS65_LH_MX41X7 U558 ( .D0(n523), .S0(n196), .D1(\alu_i[SRC_B][28] ), .S1(n32), .D2(\alu_i[SRC_B][27] ), .S2(n27), .D3(n520), .S3(n21), .Z(n255) );
  HS65_LH_AO212X4 U559 ( .A(n226), .B(n591), .C(n227), .D(\alu_i[SHAMT][4] ), 
        .E(n228), .Z(n225) );
  HS65_LH_AO222X4 U560 ( .A(n192), .B(n229), .C(n193), .D(n230), .E(n195), .F(
        n231), .Z(n228) );
  HS65_LH_MX41X7 U561 ( .D0(n524), .S0(n37), .D1(n523), .S1(n32), .D2(
        \alu_i[SRC_B][28] ), .S2(n27), .D3(\alu_i[SRC_B][27] ), .S3(n21), .Z(
        n230) );
  HS65_LH_NAND3X5 U562 ( .A(n430), .B(n431), .C(n432), .Z(\alu_o[RESULT][0] )
         );
  HS65_LH_AOI22X6 U563 ( .A(n581), .B(n444), .C(n45), .D(\HI_LO_c[LO][0] ), 
        .Z(n430) );
  HS65_LH_AOI212X4 U564 ( .A(n13), .B(n70), .C(N131), .D(n53), .E(n433), .Z(
        n432) );
  HS65_LH_AOI212X4 U565 ( .A(N99), .B(n48), .C(n69), .D(n439), .E(n440), .Z(
        n431) );
  HS65_LH_BFX9 U566 ( .A(n196), .Z(n36) );
  HS65_LH_NOR2X6 U567 ( .A(\alu_i[SHAMT][0] ), .B(\alu_i[SHAMT][1] ), .Z(n196)
         );
  HS65_LH_AO212X4 U568 ( .A(n152), .B(n591), .C(n239), .D(\alu_i[SHAMT][4] ), 
        .E(n240), .Z(n234) );
  HS65_LH_AO222X4 U569 ( .A(n192), .B(n157), .C(n193), .D(n241), .E(n195), .F(
        n154), .Z(n240) );
  HS65_LH_MX41X7 U570 ( .D0(\alu_i[SRC_B][2] ), .S0(n36), .D1(
        \alu_i[SRC_B][3] ), .S1(n32), .D2(\alu_i[SRC_B][4] ), .S2(n27), .D3(
        n74), .S3(n21), .Z(n241) );
  HS65_LH_AO212X4 U571 ( .A(n209), .B(n591), .C(n210), .D(\alu_i[SHAMT][4] ), 
        .E(n211), .Z(n203) );
  HS65_LH_AO222X4 U572 ( .A(n192), .B(n212), .C(n193), .D(n213), .E(n195), .F(
        n214), .Z(n211) );
  HS65_LH_AO212X4 U573 ( .A(n27), .B(n523), .C(n35), .D(n524), .E(n215), .Z(
        n213) );
  HS65_LH_AO12X9 U574 ( .A(\alu_i[SRC_B][28] ), .B(n21), .C(n216), .Z(n215) );
  HS65_LH_BFX9 U575 ( .A(\alu_i[SRC_B][0] ), .Z(n69) );
  HS65_LH_IVX9 U576 ( .A(\alu_i[OP][1] ), .Z(n588) );
  HS65_LH_IVX9 U577 ( .A(\alu_i[OP][0] ), .Z(n590) );
  HS65_LH_IVX9 U578 ( .A(\alu_i[OP][3] ), .Z(n587) );
  HS65_LH_IVX9 U579 ( .A(\alu_i[SRC_B][31] ), .Z(n525) );
  HS65_LH_IVX9 U580 ( .A(\alu_i[SRC_B][2] ), .Z(n71) );
  HS65_LH_IVX9 U581 ( .A(\alu_i[SRC_B][3] ), .Z(n72) );
  HS65_LH_IVX9 U582 ( .A(\alu_i[SRC_B][28] ), .Z(n522) );
  HS65_LH_IVX9 U583 ( .A(\alu_i[SRC_A][29] ), .Z(n535) );
  HS65_LH_BFX9 U584 ( .A(n104), .Z(n46) );
  HS65_LH_OAI21X3 U585 ( .A(\alu_i[OP][0] ), .B(n437), .C(n443), .Z(n104) );
  HS65_LH_OAI21X3 U586 ( .A(n436), .B(n435), .C(n390), .Z(n443) );
  HS65_LH_BFX9 U587 ( .A(n198), .Z(n26) );
  HS65_LH_NOR2AX3 U588 ( .A(\alu_i[SHAMT][1] ), .B(\alu_i[SHAMT][0] ), .Z(n198) );
  HS65_LH_IVX9 U589 ( .A(\alu_i[SRC_B][4] ), .Z(n73) );
  HS65_LH_IVX9 U590 ( .A(\alu_i[SRC_B][11] ), .Z(n80) );
  HS65_LH_IVX9 U591 ( .A(\alu_i[SRC_B][20] ), .Z(n89) );
  HS65_LH_IVX9 U592 ( .A(\alu_i[SRC_B][27] ), .Z(n521) );
  HS65_LH_IVX9 U593 ( .A(\alu_i[SRC_A][5] ), .Z(n527) );
  HS65_LH_IVX9 U594 ( .A(\alu_i[SRC_A][8] ), .Z(n528) );
  HS65_LH_IVX9 U595 ( .A(\alu_i[SRC_A][14] ), .Z(n530) );
  HS65_LH_IVX9 U596 ( .A(\alu_i[SRC_A][17] ), .Z(n531) );
  HS65_LH_IVX9 U597 ( .A(\alu_i[SRC_A][23] ), .Z(n533) );
  HS65_LH_IVX9 U598 ( .A(\alu_i[SRC_A][26] ), .Z(n534) );
  HS65_LH_IVX9 U599 ( .A(\alu_i[SRC_A][2] ), .Z(n526) );
  HS65_LH_IVX9 U600 ( .A(\alu_i[SRC_A][11] ), .Z(n529) );
  HS65_LH_IVX9 U601 ( .A(\alu_i[SRC_A][20] ), .Z(n532) );
  HS65_LH_BFX9 U602 ( .A(rst_n), .Z(n537) );
  HS65_LH_BFX9 U603 ( .A(rst_n), .Z(n536) );
  HS65_LH_AO112X9 U604 ( .A(N714), .B(n450), .C(n451), .D(n452), .Z(
        \alu_o[BRANCH] ) );
  HS65_LH_AO222X4 U605 ( .A(n391), .B(n450), .C(n438), .D(n450), .E(n436), .F(
        n450), .Z(n452) );
  HS65_LH_NOR4ABX2 U606 ( .A(N715), .B(n587), .C(n578), .D(n589), .Z(n451) );
  HS65_LH_NOR3X4 U607 ( .A(\alu_i[OP][2] ), .B(\alu_i[OP][3] ), .C(n578), .Z(
        n450) );
  HS65_LH_NAND2X7 U608 ( .A(n257), .B(n258), .Z(\alu_o[RESULT][28] ) );
  HS65_LH_AOI212X4 U609 ( .A(n12), .B(n523), .C(N159), .D(n53), .E(n270), .Z(
        n257) );
  HS65_LH_AOI212X4 U610 ( .A(N127), .B(n48), .C(n584), .D(n259), .E(n260), .Z(
        n258) );
  HS65_LH_AO222X4 U611 ( .A(\HI_LO_c[LO][28] ), .B(n45), .C(n81), .D(n106), 
        .E(\HI_LO_c[HI][28] ), .F(n16), .Z(n270) );
  HS65_LH_NAND2X7 U612 ( .A(n201), .B(n202), .Z(\alu_o[RESULT][31] ) );
  HS65_LH_AOI212X4 U613 ( .A(n16), .B(\HI_LO_c[HI][31] ), .C(N162), .D(n53), 
        .E(n217), .Z(n201) );
  HS65_LH_AOI212X4 U614 ( .A(N130), .B(n48), .C(n584), .D(n203), .E(n204), .Z(
        n202) );
  HS65_LH_AO22X9 U615 ( .A(\HI_LO_c[LO][31] ), .B(n45), .C(n84), .D(n106), .Z(
        n217) );
  HS65_LH_NAND2X7 U616 ( .A(n232), .B(n233), .Z(\alu_o[RESULT][2] ) );
  HS65_LH_AOI212X4 U617 ( .A(n13), .B(\alu_i[SRC_B][3] ), .C(N133), .D(n53), 
        .E(n242), .Z(n232) );
  HS65_LH_AOI212X4 U618 ( .A(N101), .B(n48), .C(n581), .D(n234), .E(n235), .Z(
        n233) );
  HS65_LH_AO22X9 U619 ( .A(\HI_LO_c[HI][2] ), .B(n16), .C(\HI_LO_c[LO][2] ), 
        .D(n45), .Z(n242) );
  HS65_LH_NAND2X7 U620 ( .A(n181), .B(n182), .Z(\alu_o[RESULT][3] ) );
  HS65_LH_AOI212X4 U621 ( .A(n13), .B(\alu_i[SRC_B][4] ), .C(N134), .D(n53), 
        .E(n200), .Z(n181) );
  HS65_LH_AOI212X4 U622 ( .A(N102), .B(n48), .C(n581), .D(n183), .E(n184), .Z(
        n182) );
  HS65_LH_AO22X9 U623 ( .A(\HI_LO_c[HI][3] ), .B(n16), .C(\HI_LO_c[LO][3] ), 
        .D(n45), .Z(n200) );
  HS65_LH_AO22X9 U624 ( .A(\HI_LO_c[HI][1] ), .B(n16), .C(\HI_LO_c[LO][1] ), 
        .D(n45), .Z(n356) );
  HS65_LH_IVX9 U625 ( .A(\alu_i[SRC_A][0] ), .Z(n565) );
  HS65_LH_IVX9 U626 ( .A(\alu_i[SRC_A][1] ), .Z(n564) );
  HS65_LH_IVX9 U627 ( .A(\alu_i[SRC_A][30] ), .Z(n545) );
  HS65_LH_IVX9 U628 ( .A(\alu_i[SRC_A][3] ), .Z(n563) );
  HS65_LH_IVX9 U629 ( .A(\alu_i[SRC_A][28] ), .Z(n546) );
endmodule


module alu_top ( clk, rst_n, src_a, src_b, op, shamt, result, branch );
  input [31:0] src_a;
  input [31:0] src_b;
  input [4:0] op;
  input [4:0] shamt;
  output [31:0] result;
  input clk, rst_n;
  output branch;


  alu alu_inst ( .clk(clk), .rst_n(rst_n), .alu_i({src_a, src_b, op, shamt}), 
        .alu_o({branch, result}) );
endmodule

