
library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity regfile is

   port( clk, rst_n : in std_logic;  regfile_i : in std_logic_vector (49 downto
         0);  regfile_o : out std_logic_vector (63 downto 0));

end regfile;

architecture SYN_Behavioral of regfile is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI222X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPRQNX9
      port( D, CP, RN : in std_logic;  QN : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal registers_13_31_port, registers_13_30_port, registers_13_29_port, 
      registers_13_28_port, registers_13_27_port, registers_13_26_port, 
      registers_13_25_port, registers_13_24_port, registers_13_23_port, 
      registers_13_22_port, registers_13_21_port, registers_13_20_port, 
      registers_13_19_port, registers_13_18_port, registers_13_17_port, 
      registers_13_16_port, registers_13_15_port, registers_13_14_port, 
      registers_13_13_port, registers_13_12_port, registers_13_11_port, 
      registers_13_10_port, registers_13_9_port, registers_13_8_port, 
      registers_13_7_port, registers_13_6_port, registers_13_5_port, 
      registers_13_4_port, registers_13_3_port, registers_13_2_port, 
      registers_13_1_port, registers_13_0_port, registers_12_31_port, 
      registers_12_30_port, registers_12_29_port, registers_12_28_port, 
      registers_12_27_port, registers_12_26_port, registers_12_25_port, 
      registers_12_24_port, registers_12_23_port, registers_12_22_port, 
      registers_12_21_port, registers_12_20_port, registers_12_19_port, 
      registers_12_18_port, registers_12_17_port, registers_12_16_port, 
      registers_12_15_port, registers_12_14_port, registers_12_13_port, 
      registers_12_12_port, registers_12_11_port, registers_12_10_port, 
      registers_12_9_port, registers_12_8_port, registers_12_7_port, 
      registers_12_6_port, registers_12_5_port, registers_12_4_port, 
      registers_12_3_port, registers_12_2_port, registers_12_1_port, 
      registers_12_0_port, registers_11_31_port, registers_11_30_port, 
      registers_11_29_port, registers_11_28_port, registers_11_27_port, 
      registers_11_26_port, registers_11_25_port, registers_11_24_port, 
      registers_11_23_port, registers_11_22_port, registers_11_21_port, 
      registers_11_20_port, registers_11_19_port, registers_11_18_port, 
      registers_11_17_port, registers_11_16_port, registers_11_15_port, 
      registers_11_14_port, registers_11_13_port, registers_11_12_port, 
      registers_11_11_port, registers_11_10_port, registers_11_9_port, 
      registers_11_8_port, registers_11_7_port, registers_11_6_port, 
      registers_11_5_port, registers_11_4_port, registers_11_3_port, 
      registers_11_2_port, registers_11_1_port, registers_11_0_port, 
      registers_10_31_port, registers_10_30_port, registers_10_29_port, 
      registers_10_28_port, registers_10_27_port, registers_10_26_port, 
      registers_10_25_port, registers_10_24_port, registers_10_23_port, 
      registers_10_22_port, registers_10_21_port, registers_10_20_port, 
      registers_10_19_port, registers_10_18_port, registers_10_17_port, 
      registers_10_16_port, registers_10_15_port, registers_10_14_port, 
      registers_10_13_port, registers_10_12_port, registers_10_11_port, 
      registers_10_10_port, registers_10_9_port, registers_10_8_port, 
      registers_10_7_port, registers_10_6_port, registers_10_5_port, 
      registers_10_4_port, registers_10_3_port, registers_10_2_port, 
      registers_10_1_port, registers_10_0_port, registers_7_31_port, 
      registers_7_30_port, registers_7_29_port, registers_7_28_port, 
      registers_7_27_port, registers_7_26_port, registers_7_25_port, 
      registers_7_24_port, registers_7_23_port, registers_7_22_port, 
      registers_7_21_port, registers_7_20_port, registers_7_19_port, 
      registers_7_18_port, registers_7_17_port, registers_7_16_port, 
      registers_7_15_port, registers_7_14_port, registers_7_13_port, 
      registers_7_12_port, registers_7_11_port, registers_7_10_port, 
      registers_7_9_port, registers_7_8_port, registers_7_7_port, 
      registers_7_6_port, registers_7_5_port, registers_7_4_port, 
      registers_7_3_port, registers_7_2_port, registers_7_1_port, 
      registers_7_0_port, registers_6_31_port, registers_6_30_port, 
      registers_6_29_port, registers_6_28_port, registers_6_27_port, 
      registers_6_26_port, registers_6_25_port, registers_6_24_port, 
      registers_6_23_port, registers_6_22_port, registers_6_21_port, 
      registers_6_20_port, registers_6_19_port, registers_6_18_port, 
      registers_6_17_port, registers_6_16_port, registers_6_15_port, 
      registers_6_14_port, registers_6_13_port, registers_6_12_port, 
      registers_6_11_port, registers_6_10_port, registers_6_9_port, 
      registers_6_8_port, registers_6_7_port, registers_6_6_port, 
      registers_6_5_port, registers_6_4_port, registers_6_3_port, 
      registers_6_2_port, registers_6_1_port, registers_6_0_port, 
      registers_5_31_port, registers_5_30_port, registers_5_29_port, 
      registers_5_28_port, registers_5_27_port, registers_5_26_port, 
      registers_5_25_port, registers_5_24_port, registers_5_23_port, 
      registers_5_22_port, registers_5_21_port, registers_5_20_port, 
      registers_5_19_port, registers_5_18_port, registers_5_17_port, 
      registers_5_16_port, registers_5_15_port, registers_5_14_port, 
      registers_5_13_port, registers_5_12_port, registers_5_11_port, 
      registers_5_10_port, registers_5_9_port, registers_5_8_port, 
      registers_5_7_port, registers_5_6_port, registers_5_5_port, 
      registers_5_4_port, registers_5_3_port, registers_5_2_port, 
      registers_5_1_port, registers_5_0_port, registers_4_31_port, 
      registers_4_30_port, registers_4_29_port, registers_4_28_port, 
      registers_4_27_port, registers_4_26_port, registers_4_25_port, 
      registers_4_24_port, registers_4_23_port, registers_4_22_port, 
      registers_4_21_port, registers_4_20_port, registers_4_19_port, 
      registers_4_18_port, registers_4_17_port, registers_4_16_port, 
      registers_4_15_port, registers_4_14_port, registers_4_13_port, 
      registers_4_12_port, registers_4_11_port, registers_4_10_port, 
      registers_4_9_port, registers_4_8_port, registers_4_7_port, 
      registers_4_6_port, registers_4_5_port, registers_4_4_port, 
      registers_4_3_port, registers_4_2_port, registers_4_1_port, 
      registers_4_0_port, registers_3_31_port, registers_3_30_port, 
      registers_3_29_port, registers_3_28_port, registers_3_27_port, 
      registers_3_26_port, registers_3_25_port, registers_3_24_port, 
      registers_3_23_port, registers_3_22_port, registers_3_21_port, 
      registers_3_20_port, registers_3_19_port, registers_3_18_port, 
      registers_3_17_port, registers_3_16_port, registers_3_15_port, 
      registers_3_14_port, registers_3_13_port, registers_3_12_port, 
      registers_3_11_port, registers_3_10_port, registers_3_9_port, 
      registers_3_8_port, registers_3_7_port, registers_3_6_port, 
      registers_3_5_port, registers_3_4_port, registers_3_3_port, 
      registers_3_2_port, registers_3_1_port, registers_3_0_port, 
      registers_2_31_port, registers_2_30_port, registers_2_29_port, 
      registers_2_28_port, registers_2_27_port, registers_2_26_port, 
      registers_2_25_port, registers_2_24_port, registers_2_23_port, 
      registers_2_22_port, registers_2_21_port, registers_2_20_port, 
      registers_2_19_port, registers_2_18_port, registers_2_17_port, 
      registers_2_16_port, registers_2_15_port, registers_2_14_port, 
      registers_2_13_port, registers_2_12_port, registers_2_11_port, 
      registers_2_10_port, registers_2_9_port, registers_2_8_port, 
      registers_2_7_port, registers_2_6_port, registers_2_5_port, 
      registers_2_4_port, registers_2_3_port, registers_2_2_port, 
      registers_2_1_port, registers_2_0_port, registers_1_31_port, 
      registers_1_30_port, registers_1_29_port, registers_1_28_port, 
      registers_1_27_port, registers_1_26_port, registers_1_25_port, 
      registers_1_24_port, registers_1_23_port, registers_1_22_port, 
      registers_1_21_port, registers_1_20_port, registers_1_19_port, 
      registers_1_18_port, registers_1_17_port, registers_1_16_port, 
      registers_1_15_port, registers_1_14_port, registers_1_13_port, 
      registers_1_12_port, registers_1_11_port, registers_1_10_port, 
      registers_1_9_port, registers_1_8_port, registers_1_7_port, 
      registers_1_6_port, registers_1_5_port, registers_1_4_port, 
      registers_1_3_port, registers_1_2_port, registers_1_1_port, 
      registers_1_0_port, registers_31_31_port, registers_31_30_port, 
      registers_31_29_port, registers_31_28_port, registers_31_27_port, 
      registers_31_26_port, registers_31_25_port, registers_31_24_port, 
      registers_31_23_port, registers_31_22_port, registers_31_21_port, 
      registers_31_20_port, registers_31_19_port, registers_31_18_port, 
      registers_31_17_port, registers_31_16_port, registers_31_15_port, 
      registers_31_14_port, registers_31_13_port, registers_31_12_port, 
      registers_31_11_port, registers_31_10_port, registers_31_9_port, 
      registers_31_8_port, registers_31_7_port, registers_31_6_port, 
      registers_31_5_port, registers_31_4_port, registers_31_3_port, 
      registers_31_2_port, registers_31_1_port, registers_31_0_port, 
      registers_30_31_port, registers_30_30_port, registers_30_29_port, 
      registers_30_28_port, registers_30_27_port, registers_30_26_port, 
      registers_30_25_port, registers_30_24_port, registers_30_23_port, 
      registers_30_22_port, registers_30_21_port, registers_30_20_port, 
      registers_30_19_port, registers_30_18_port, registers_30_17_port, 
      registers_30_16_port, registers_30_15_port, registers_30_14_port, 
      registers_30_13_port, registers_30_12_port, registers_30_11_port, 
      registers_30_10_port, registers_30_9_port, registers_30_8_port, 
      registers_30_7_port, registers_30_6_port, registers_30_5_port, 
      registers_30_4_port, registers_30_3_port, registers_30_2_port, 
      registers_30_1_port, registers_30_0_port, registers_25_31_port, 
      registers_25_30_port, registers_25_29_port, registers_25_28_port, 
      registers_25_27_port, registers_25_26_port, registers_25_25_port, 
      registers_25_24_port, registers_25_23_port, registers_25_22_port, 
      registers_25_21_port, registers_25_20_port, registers_25_19_port, 
      registers_25_18_port, registers_25_17_port, registers_25_16_port, 
      registers_25_15_port, registers_25_14_port, registers_25_13_port, 
      registers_25_12_port, registers_25_11_port, registers_25_10_port, 
      registers_25_9_port, registers_25_8_port, registers_25_7_port, 
      registers_25_6_port, registers_25_5_port, registers_25_4_port, 
      registers_25_3_port, registers_25_2_port, registers_25_1_port, 
      registers_25_0_port, registers_24_31_port, registers_24_30_port, 
      registers_24_29_port, registers_24_28_port, registers_24_27_port, 
      registers_24_26_port, registers_24_25_port, registers_24_24_port, 
      registers_24_23_port, registers_24_22_port, registers_24_21_port, 
      registers_24_20_port, registers_24_19_port, registers_24_18_port, 
      registers_24_17_port, registers_24_16_port, registers_24_15_port, 
      registers_24_14_port, registers_24_13_port, registers_24_12_port, 
      registers_24_11_port, registers_24_10_port, registers_24_9_port, 
      registers_24_8_port, registers_24_7_port, registers_24_6_port, 
      registers_24_5_port, registers_24_4_port, registers_24_3_port, 
      registers_24_2_port, registers_24_1_port, registers_24_0_port, 
      registers_23_31_port, registers_23_30_port, registers_23_29_port, 
      registers_23_28_port, registers_23_27_port, registers_23_26_port, 
      registers_23_25_port, registers_23_24_port, registers_23_23_port, 
      registers_23_22_port, registers_23_21_port, registers_23_20_port, 
      registers_23_19_port, registers_23_18_port, registers_23_17_port, 
      registers_23_16_port, registers_23_15_port, registers_23_14_port, 
      registers_23_13_port, registers_23_12_port, registers_23_11_port, 
      registers_23_10_port, registers_23_9_port, registers_23_8_port, 
      registers_23_7_port, registers_23_6_port, registers_23_5_port, 
      registers_23_4_port, registers_23_3_port, registers_23_2_port, 
      registers_23_1_port, registers_23_0_port, registers_22_31_port, 
      registers_22_30_port, registers_22_29_port, registers_22_28_port, 
      registers_22_27_port, registers_22_26_port, registers_22_25_port, 
      registers_22_24_port, registers_22_23_port, registers_22_22_port, 
      registers_22_21_port, registers_22_20_port, registers_22_19_port, 
      registers_22_18_port, registers_22_17_port, registers_22_16_port, 
      registers_22_15_port, registers_22_14_port, registers_22_13_port, 
      registers_22_12_port, registers_22_11_port, registers_22_10_port, 
      registers_22_9_port, registers_22_8_port, registers_22_7_port, 
      registers_22_6_port, registers_22_5_port, registers_22_4_port, 
      registers_22_3_port, registers_22_2_port, registers_22_1_port, 
      registers_22_0_port, registers_21_31_port, registers_21_30_port, 
      registers_21_29_port, registers_21_28_port, registers_21_27_port, 
      registers_21_26_port, registers_21_25_port, registers_21_24_port, 
      registers_21_23_port, registers_21_22_port, registers_21_21_port, 
      registers_21_20_port, registers_21_19_port, registers_21_18_port, 
      registers_21_17_port, registers_21_16_port, registers_21_15_port, 
      registers_21_14_port, registers_21_13_port, registers_21_12_port, 
      registers_21_11_port, registers_21_10_port, registers_21_9_port, 
      registers_21_8_port, registers_21_7_port, registers_21_6_port, 
      registers_21_5_port, registers_21_4_port, registers_21_3_port, 
      registers_21_2_port, registers_21_1_port, registers_21_0_port, 
      registers_20_31_port, registers_20_30_port, registers_20_29_port, 
      registers_20_28_port, registers_20_27_port, registers_20_26_port, 
      registers_20_25_port, registers_20_24_port, registers_20_23_port, 
      registers_20_22_port, registers_20_21_port, registers_20_20_port, 
      registers_20_19_port, registers_20_18_port, registers_20_17_port, 
      registers_20_16_port, registers_20_15_port, registers_20_14_port, 
      registers_20_13_port, registers_20_12_port, registers_20_11_port, 
      registers_20_10_port, registers_20_9_port, registers_20_8_port, 
      registers_20_7_port, registers_20_6_port, registers_20_5_port, 
      registers_20_4_port, registers_20_3_port, registers_20_2_port, 
      registers_20_1_port, registers_20_0_port, registers_19_31_port, 
      registers_19_30_port, registers_19_29_port, registers_19_28_port, 
      registers_19_27_port, registers_19_26_port, registers_19_25_port, 
      registers_19_24_port, registers_19_23_port, registers_19_22_port, 
      registers_19_21_port, registers_19_20_port, registers_19_19_port, 
      registers_19_18_port, registers_19_17_port, registers_19_16_port, 
      registers_19_15_port, registers_19_14_port, registers_19_13_port, 
      registers_19_12_port, registers_19_11_port, registers_19_10_port, 
      registers_19_9_port, registers_19_8_port, registers_19_7_port, 
      registers_19_6_port, registers_19_5_port, registers_19_4_port, 
      registers_19_3_port, registers_19_2_port, registers_19_1_port, 
      registers_19_0_port, registers_18_31_port, registers_18_30_port, 
      registers_18_29_port, registers_18_28_port, registers_18_27_port, 
      registers_18_26_port, registers_18_25_port, registers_18_24_port, 
      registers_18_23_port, registers_18_22_port, registers_18_21_port, 
      registers_18_20_port, registers_18_19_port, registers_18_18_port, 
      registers_18_17_port, registers_18_16_port, registers_18_15_port, 
      registers_18_14_port, registers_18_13_port, registers_18_12_port, 
      registers_18_11_port, registers_18_10_port, registers_18_9_port, 
      registers_18_8_port, registers_18_7_port, registers_18_6_port, 
      registers_18_5_port, registers_18_4_port, registers_18_3_port, 
      registers_18_2_port, registers_18_1_port, registers_18_0_port, 
      registers_17_31_port, registers_17_30_port, registers_17_29_port, 
      registers_17_28_port, registers_17_27_port, registers_17_26_port, 
      registers_17_25_port, registers_17_24_port, registers_17_23_port, 
      registers_17_22_port, registers_17_21_port, registers_17_20_port, 
      registers_17_19_port, registers_17_18_port, registers_17_17_port, 
      registers_17_16_port, registers_17_15_port, registers_17_14_port, 
      registers_17_13_port, registers_17_12_port, registers_17_11_port, 
      registers_17_10_port, registers_17_9_port, registers_17_8_port, 
      registers_17_7_port, registers_17_6_port, registers_17_5_port, 
      registers_17_4_port, registers_17_3_port, registers_17_2_port, 
      registers_17_1_port, registers_17_0_port, registers_16_31_port, 
      registers_16_30_port, registers_16_29_port, registers_16_28_port, 
      registers_16_27_port, registers_16_26_port, registers_16_25_port, 
      registers_16_24_port, registers_16_23_port, registers_16_22_port, 
      registers_16_21_port, registers_16_20_port, registers_16_19_port, 
      registers_16_18_port, registers_16_17_port, registers_16_16_port, 
      registers_16_15_port, registers_16_14_port, registers_16_13_port, 
      registers_16_12_port, registers_16_11_port, registers_16_10_port, 
      registers_16_9_port, registers_16_8_port, registers_16_7_port, 
      registers_16_6_port, registers_16_5_port, registers_16_4_port, 
      registers_16_3_port, registers_16_2_port, registers_16_1_port, 
      registers_16_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n257, n258, n259, n260, n261, n262, n263, n264, n265
      , n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
      n770, n771, n772, n773, n774, n775, n776, n777, n778, n795, n811, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
      n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, 
      n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
      n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, 
      n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
      n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, 
      n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
      n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, 
      n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
      n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, 
      n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, 
      n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
      n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, 
      n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, 
      n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, 
      n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, 
      n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, 
      n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, 
      n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, 
      n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, 
      n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, 
      n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, 
      n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
      n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, 
      n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, 
      n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, 
      n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, 
      n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, 
      n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
      n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, 
      n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, 
      n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, 
      n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, 
      n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, 
      n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
      n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
      n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
      n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
      n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, 
      n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, 
      n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, 
      n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, 
      n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, 
      n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
      n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
      n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, 
      n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
      n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
      n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, 
      n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
      n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
      n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2824, n2825, n2827, 
      n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, 
      n2838, n2839, n2841, n2846, n2847, n2848, n2849, n2850, n2851, n2853, 
      n2855, n2856, n2857, n2859, n2860, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664 : std_logic;

begin
   
   registers_reg_31_31_inst : HS65_LH_DFPRQX9 port map( D => n2425, CP => clk, 
                           RN => n6539, Q => registers_31_31_port);
   registers_reg_31_30_inst : HS65_LH_DFPRQX9 port map( D => n2424, CP => clk, 
                           RN => n6569, Q => registers_31_30_port);
   registers_reg_31_29_inst : HS65_LH_DFPRQX9 port map( D => n2423, CP => clk, 
                           RN => n6571, Q => registers_31_29_port);
   registers_reg_31_28_inst : HS65_LH_DFPRQX9 port map( D => n2422, CP => clk, 
                           RN => n6570, Q => registers_31_28_port);
   registers_reg_31_27_inst : HS65_LH_DFPRQX9 port map( D => n2421, CP => clk, 
                           RN => n6570, Q => registers_31_27_port);
   registers_reg_31_26_inst : HS65_LH_DFPRQX9 port map( D => n2420, CP => clk, 
                           RN => n6569, Q => registers_31_26_port);
   registers_reg_31_25_inst : HS65_LH_DFPRQX9 port map( D => n2419, CP => clk, 
                           RN => n6572, Q => registers_31_25_port);
   registers_reg_31_24_inst : HS65_LH_DFPRQX9 port map( D => n2418, CP => clk, 
                           RN => n6572, Q => registers_31_24_port);
   registers_reg_31_23_inst : HS65_LH_DFPRQX9 port map( D => n2417, CP => clk, 
                           RN => n6572, Q => registers_31_23_port);
   registers_reg_31_22_inst : HS65_LH_DFPRQX9 port map( D => n2416, CP => clk, 
                           RN => n6572, Q => registers_31_22_port);
   registers_reg_31_21_inst : HS65_LH_DFPRQX9 port map( D => n2415, CP => clk, 
                           RN => n6568, Q => registers_31_21_port);
   registers_reg_31_20_inst : HS65_LH_DFPRQX9 port map( D => n2414, CP => clk, 
                           RN => n6568, Q => registers_31_20_port);
   registers_reg_31_19_inst : HS65_LH_DFPRQX9 port map( D => n2413, CP => clk, 
                           RN => n6568, Q => registers_31_19_port);
   registers_reg_31_18_inst : HS65_LH_DFPRQX9 port map( D => n2412, CP => clk, 
                           RN => n6568, Q => registers_31_18_port);
   registers_reg_31_17_inst : HS65_LH_DFPRQX9 port map( D => n2411, CP => clk, 
                           RN => n6568, Q => registers_31_17_port);
   registers_reg_31_16_inst : HS65_LH_DFPRQX9 port map( D => n2410, CP => clk, 
                           RN => n6568, Q => registers_31_16_port);
   registers_reg_31_15_inst : HS65_LH_DFPRQX9 port map( D => n2409, CP => clk, 
                           RN => n6568, Q => registers_31_15_port);
   registers_reg_31_14_inst : HS65_LH_DFPRQX9 port map( D => n2408, CP => clk, 
                           RN => n6568, Q => registers_31_14_port);
   registers_reg_31_13_inst : HS65_LH_DFPRQX9 port map( D => n2407, CP => clk, 
                           RN => n6578, Q => registers_31_13_port);
   registers_reg_31_12_inst : HS65_LH_DFPRQX9 port map( D => n2406, CP => clk, 
                           RN => n6578, Q => registers_31_12_port);
   registers_reg_31_11_inst : HS65_LH_DFPRQX9 port map( D => n2405, CP => clk, 
                           RN => n6578, Q => registers_31_11_port);
   registers_reg_31_10_inst : HS65_LH_DFPRQX9 port map( D => n2404, CP => clk, 
                           RN => n6578, Q => registers_31_10_port);
   registers_reg_31_9_inst : HS65_LH_DFPRQX9 port map( D => n2403, CP => clk, 
                           RN => n6580, Q => registers_31_9_port);
   registers_reg_31_8_inst : HS65_LH_DFPRQX9 port map( D => n2402, CP => clk, 
                           RN => n6580, Q => registers_31_8_port);
   registers_reg_31_7_inst : HS65_LH_DFPRQX9 port map( D => n2401, CP => clk, 
                           RN => n6580, Q => registers_31_7_port);
   registers_reg_31_6_inst : HS65_LH_DFPRQX9 port map( D => n2400, CP => clk, 
                           RN => n6580, Q => registers_31_6_port);
   registers_reg_31_5_inst : HS65_LH_DFPRQX9 port map( D => n2399, CP => clk, 
                           RN => n6580, Q => registers_31_5_port);
   registers_reg_31_4_inst : HS65_LH_DFPRQX9 port map( D => n2398, CP => clk, 
                           RN => n6580, Q => registers_31_4_port);
   registers_reg_31_3_inst : HS65_LH_DFPRQX9 port map( D => n2397, CP => clk, 
                           RN => n6580, Q => registers_31_3_port);
   registers_reg_31_2_inst : HS65_LH_DFPRQX9 port map( D => n2396, CP => clk, 
                           RN => n6580, Q => registers_31_2_port);
   registers_reg_31_1_inst : HS65_LH_DFPRQX9 port map( D => n2395, CP => clk, 
                           RN => n6578, Q => registers_31_1_port);
   registers_reg_31_0_inst : HS65_LH_DFPRQX9 port map( D => n2394, CP => clk, 
                           RN => n6578, Q => registers_31_0_port);
   registers_reg_30_31_inst : HS65_LH_DFPRQX9 port map( D => n2393, CP => clk, 
                           RN => n6583, Q => registers_30_31_port);
   registers_reg_30_30_inst : HS65_LH_DFPRQX9 port map( D => n2392, CP => clk, 
                           RN => n6583, Q => registers_30_30_port);
   registers_reg_30_29_inst : HS65_LH_DFPRQX9 port map( D => n2391, CP => clk, 
                           RN => n6583, Q => registers_30_29_port);
   registers_reg_30_28_inst : HS65_LH_DFPRQX9 port map( D => n2390, CP => clk, 
                           RN => n6583, Q => registers_30_28_port);
   registers_reg_30_27_inst : HS65_LH_DFPRQX9 port map( D => n2389, CP => clk, 
                           RN => n6584, Q => registers_30_27_port);
   registers_reg_30_26_inst : HS65_LH_DFPRQX9 port map( D => n2388, CP => clk, 
                           RN => n6584, Q => registers_30_26_port);
   registers_reg_30_25_inst : HS65_LH_DFPRQX9 port map( D => n2387, CP => clk, 
                           RN => n6584, Q => registers_30_25_port);
   registers_reg_30_24_inst : HS65_LH_DFPRQX9 port map( D => n2386, CP => clk, 
                           RN => n6584, Q => registers_30_24_port);
   registers_reg_30_23_inst : HS65_LH_DFPRQX9 port map( D => n2385, CP => clk, 
                           RN => n6579, Q => registers_30_23_port);
   registers_reg_30_22_inst : HS65_LH_DFPRQX9 port map( D => n2384, CP => clk, 
                           RN => n6579, Q => registers_30_22_port);
   registers_reg_30_21_inst : HS65_LH_DFPRQX9 port map( D => n2383, CP => clk, 
                           RN => n6585, Q => registers_30_21_port);
   registers_reg_30_20_inst : HS65_LH_DFPRQX9 port map( D => n2382, CP => clk, 
                           RN => n6583, Q => registers_30_20_port);
   registers_reg_30_19_inst : HS65_LH_DFPRQX9 port map( D => n2381, CP => clk, 
                           RN => n6583, Q => registers_30_19_port);
   registers_reg_30_18_inst : HS65_LH_DFPRQX9 port map( D => n2380, CP => clk, 
                           RN => n6583, Q => registers_30_18_port);
   registers_reg_30_17_inst : HS65_LH_DFPRQX9 port map( D => n2379, CP => clk, 
                           RN => n6582, Q => registers_30_17_port);
   registers_reg_30_16_inst : HS65_LH_DFPRQX9 port map( D => n2378, CP => clk, 
                           RN => n6582, Q => registers_30_16_port);
   registers_reg_30_15_inst : HS65_LH_DFPRQX9 port map( D => n2377, CP => clk, 
                           RN => n6582, Q => registers_30_15_port);
   registers_reg_30_14_inst : HS65_LH_DFPRQX9 port map( D => n2376, CP => clk, 
                           RN => n6582, Q => registers_30_14_port);
   registers_reg_30_13_inst : HS65_LH_DFPRQX9 port map( D => n2375, CP => clk, 
                           RN => n6582, Q => registers_30_13_port);
   registers_reg_30_12_inst : HS65_LH_DFPRQX9 port map( D => n2374, CP => clk, 
                           RN => n6582, Q => registers_30_12_port);
   registers_reg_30_11_inst : HS65_LH_DFPRQX9 port map( D => n2373, CP => clk, 
                           RN => n6582, Q => registers_30_11_port);
   registers_reg_30_10_inst : HS65_LH_DFPRQX9 port map( D => n2372, CP => clk, 
                           RN => n6582, Q => registers_30_10_port);
   registers_reg_30_9_inst : HS65_LH_DFPRQX9 port map( D => n2371, CP => clk, 
                           RN => n6583, Q => registers_30_9_port);
   registers_reg_30_8_inst : HS65_LH_DFPRQX9 port map( D => n2370, CP => clk, 
                           RN => n6583, Q => registers_30_8_port);
   registers_reg_30_7_inst : HS65_LH_DFPRQX9 port map( D => n2369, CP => clk, 
                           RN => n6585, Q => registers_30_7_port);
   registers_reg_30_6_inst : HS65_LH_DFPRQX9 port map( D => n2368, CP => clk, 
                           RN => n6585, Q => registers_30_6_port);
   registers_reg_30_5_inst : HS65_LH_DFPRQX9 port map( D => n2367, CP => clk, 
                           RN => n6585, Q => registers_30_5_port);
   registers_reg_30_4_inst : HS65_LH_DFPRQX9 port map( D => n2366, CP => clk, 
                           RN => n6585, Q => registers_30_4_port);
   registers_reg_30_3_inst : HS65_LH_DFPRQX9 port map( D => n2365, CP => clk, 
                           RN => n6585, Q => registers_30_3_port);
   registers_reg_30_2_inst : HS65_LH_DFPRQX9 port map( D => n2364, CP => clk, 
                           RN => n6585, Q => registers_30_2_port);
   registers_reg_30_1_inst : HS65_LH_DFPRQX9 port map( D => n2363, CP => clk, 
                           RN => n6585, Q => registers_30_1_port);
   registers_reg_30_0_inst : HS65_LH_DFPRQX9 port map( D => n2362, CP => clk, 
                           RN => n6585, Q => registers_30_0_port);
   registers_reg_25_31_inst : HS65_LH_DFPRQX9 port map( D => n2233, CP => clk, 
                           RN => n6586, Q => registers_25_31_port);
   registers_reg_25_30_inst : HS65_LH_DFPRQX9 port map( D => n2232, CP => clk, 
                           RN => n6586, Q => registers_25_30_port);
   registers_reg_25_29_inst : HS65_LH_DFPRQX9 port map( D => n2231, CP => clk, 
                           RN => n6589, Q => registers_25_29_port);
   registers_reg_25_28_inst : HS65_LH_DFPRQX9 port map( D => n2230, CP => clk, 
                           RN => n6589, Q => registers_25_28_port);
   registers_reg_25_27_inst : HS65_LH_DFPRQX9 port map( D => n2229, CP => clk, 
                           RN => n6589, Q => registers_25_27_port);
   registers_reg_25_26_inst : HS65_LH_DFPRQX9 port map( D => n2228, CP => clk, 
                           RN => n6589, Q => registers_25_26_port);
   registers_reg_25_25_inst : HS65_LH_DFPRQX9 port map( D => n2227, CP => clk, 
                           RN => n6586, Q => registers_25_25_port);
   registers_reg_25_24_inst : HS65_LH_DFPRQX9 port map( D => n2226, CP => clk, 
                           RN => n6586, Q => registers_25_24_port);
   registers_reg_25_23_inst : HS65_LH_DFPRQX9 port map( D => n2225, CP => clk, 
                           RN => n6585, Q => registers_25_23_port);
   registers_reg_25_22_inst : HS65_LH_DFPRQX9 port map( D => n2224, CP => clk, 
                           RN => n6585, Q => registers_25_22_port);
   registers_reg_25_21_inst : HS65_LH_DFPRQX9 port map( D => n2223, CP => clk, 
                           RN => n6585, Q => registers_25_21_port);
   registers_reg_25_20_inst : HS65_LH_DFPRQX9 port map( D => n2222, CP => clk, 
                           RN => n6583, Q => registers_25_20_port);
   registers_reg_25_19_inst : HS65_LH_DFPRQX9 port map( D => n2221, CP => clk, 
                           RN => n6583, Q => registers_25_19_port);
   registers_reg_25_18_inst : HS65_LH_DFPRQX9 port map( D => n2220, CP => clk, 
                           RN => n6583, Q => registers_25_18_port);
   registers_reg_25_17_inst : HS65_LH_DFPRQX9 port map( D => n2219, CP => clk, 
                           RN => n6588, Q => registers_25_17_port);
   registers_reg_25_16_inst : HS65_LH_DFPRQX9 port map( D => n2218, CP => clk, 
                           RN => n6588, Q => registers_25_16_port);
   registers_reg_25_15_inst : HS65_LH_DFPRQX9 port map( D => n2217, CP => clk, 
                           RN => n6588, Q => registers_25_15_port);
   registers_reg_25_14_inst : HS65_LH_DFPRQX9 port map( D => n2216, CP => clk, 
                           RN => n6586, Q => registers_25_14_port);
   registers_reg_25_13_inst : HS65_LH_DFPRQX9 port map( D => n2215, CP => clk, 
                           RN => n6584, Q => registers_25_13_port);
   registers_reg_25_12_inst : HS65_LH_DFPRQX9 port map( D => n2214, CP => clk, 
                           RN => n6584, Q => registers_25_12_port);
   registers_reg_25_11_inst : HS65_LH_DFPRQX9 port map( D => n2213, CP => clk, 
                           RN => n6584, Q => registers_25_11_port);
   registers_reg_25_10_inst : HS65_LH_DFPRQX9 port map( D => n2212, CP => clk, 
                           RN => n6584, Q => registers_25_10_port);
   registers_reg_25_9_inst : HS65_LH_DFPRQX9 port map( D => n2211, CP => clk, 
                           RN => n6584, Q => registers_25_9_port);
   registers_reg_25_8_inst : HS65_LH_DFPRQX9 port map( D => n2210, CP => clk, 
                           RN => n6584, Q => registers_25_8_port);
   registers_reg_25_7_inst : HS65_LH_DFPRQX9 port map( D => n2209, CP => clk, 
                           RN => n6584, Q => registers_25_7_port);
   registers_reg_25_6_inst : HS65_LH_DFPRQX9 port map( D => n2208, CP => clk, 
                           RN => n6584, Q => registers_25_6_port);
   registers_reg_25_5_inst : HS65_LH_DFPRQX9 port map( D => n2207, CP => clk, 
                           RN => n6586, Q => registers_25_5_port);
   registers_reg_25_4_inst : HS65_LH_DFPRQX9 port map( D => n2206, CP => clk, 
                           RN => n6586, Q => registers_25_4_port);
   registers_reg_25_3_inst : HS65_LH_DFPRQX9 port map( D => n2205, CP => clk, 
                           RN => n6586, Q => registers_25_3_port);
   registers_reg_25_2_inst : HS65_LH_DFPRQX9 port map( D => n2204, CP => clk, 
                           RN => n6586, Q => registers_25_2_port);
   registers_reg_25_1_inst : HS65_LH_DFPRQX9 port map( D => n2203, CP => clk, 
                           RN => n6586, Q => registers_25_1_port);
   registers_reg_25_0_inst : HS65_LH_DFPRQX9 port map( D => n2202, CP => clk, 
                           RN => n6586, Q => registers_25_0_port);
   registers_reg_24_31_inst : HS65_LH_DFPRQX9 port map( D => n2201, CP => clk, 
                           RN => n6591, Q => registers_24_31_port);
   registers_reg_24_30_inst : HS65_LH_DFPRQX9 port map( D => n2200, CP => clk, 
                           RN => n6591, Q => registers_24_30_port);
   registers_reg_24_29_inst : HS65_LH_DFPRQX9 port map( D => n2199, CP => clk, 
                           RN => n6591, Q => registers_24_29_port);
   registers_reg_24_28_inst : HS65_LH_DFPRQX9 port map( D => n2198, CP => clk, 
                           RN => n6591, Q => registers_24_28_port);
   registers_reg_24_27_inst : HS65_LH_DFPRQX9 port map( D => n2197, CP => clk, 
                           RN => n6590, Q => registers_24_27_port);
   registers_reg_24_26_inst : HS65_LH_DFPRQX9 port map( D => n2196, CP => clk, 
                           RN => n6592, Q => registers_24_26_port);
   registers_reg_24_25_inst : HS65_LH_DFPRQX9 port map( D => n2195, CP => clk, 
                           RN => n6592, Q => registers_24_25_port);
   registers_reg_24_24_inst : HS65_LH_DFPRQX9 port map( D => n2194, CP => clk, 
                           RN => n6592, Q => registers_24_24_port);
   registers_reg_24_23_inst : HS65_LH_DFPRQX9 port map( D => n2193, CP => clk, 
                           RN => n6590, Q => registers_24_23_port);
   registers_reg_24_22_inst : HS65_LH_DFPRQX9 port map( D => n2192, CP => clk, 
                           RN => n6590, Q => registers_24_22_port);
   registers_reg_24_21_inst : HS65_LH_DFPRQX9 port map( D => n2191, CP => clk, 
                           RN => n6590, Q => registers_24_21_port);
   registers_reg_24_20_inst : HS65_LH_DFPRQX9 port map( D => n2190, CP => clk, 
                           RN => n6590, Q => registers_24_20_port);
   registers_reg_24_19_inst : HS65_LH_DFPRQX9 port map( D => n2189, CP => clk, 
                           RN => n6588, Q => registers_24_19_port);
   registers_reg_24_18_inst : HS65_LH_DFPRQX9 port map( D => n2188, CP => clk, 
                           RN => n6588, Q => registers_24_18_port);
   registers_reg_24_17_inst : HS65_LH_DFPRQX9 port map( D => n2187, CP => clk, 
                           RN => n6588, Q => registers_24_17_port);
   registers_reg_24_16_inst : HS65_LH_DFPRQX9 port map( D => n2186, CP => clk, 
                           RN => n6588, Q => registers_24_16_port);
   registers_reg_24_15_inst : HS65_LH_DFPRQX9 port map( D => n2185, CP => clk, 
                           RN => n6588, Q => registers_24_15_port);
   registers_reg_24_14_inst : HS65_LH_DFPRQX9 port map( D => n2184, CP => clk, 
                           RN => n6590, Q => registers_24_14_port);
   registers_reg_24_13_inst : HS65_LH_DFPRQX9 port map( D => n2183, CP => clk, 
                           RN => n6590, Q => registers_24_13_port);
   registers_reg_24_12_inst : HS65_LH_DFPRQX9 port map( D => n2182, CP => clk, 
                           RN => n6590, Q => registers_24_12_port);
   registers_reg_24_11_inst : HS65_LH_DFPRQX9 port map( D => n2181, CP => clk, 
                           RN => n6590, Q => registers_24_11_port);
   registers_reg_24_10_inst : HS65_LH_DFPRQX9 port map( D => n2180, CP => clk, 
                           RN => n6589, Q => registers_24_10_port);
   registers_reg_24_9_inst : HS65_LH_DFPRQX9 port map( D => n2179, CP => clk, 
                           RN => n6589, Q => registers_24_9_port);
   registers_reg_24_8_inst : HS65_LH_DFPRQX9 port map( D => n2178, CP => clk, 
                           RN => n6589, Q => registers_24_8_port);
   registers_reg_24_7_inst : HS65_LH_DFPRQX9 port map( D => n2177, CP => clk, 
                           RN => n6589, Q => registers_24_7_port);
   registers_reg_24_6_inst : HS65_LH_DFPRQX9 port map( D => n2176, CP => clk, 
                           RN => n6589, Q => registers_24_6_port);
   registers_reg_24_5_inst : HS65_LH_DFPRQX9 port map( D => n2175, CP => clk, 
                           RN => n6589, Q => registers_24_5_port);
   registers_reg_24_4_inst : HS65_LH_DFPRQX9 port map( D => n2174, CP => clk, 
                           RN => n6589, Q => registers_24_4_port);
   registers_reg_24_3_inst : HS65_LH_DFPRQX9 port map( D => n2173, CP => clk, 
                           RN => n6589, Q => registers_24_3_port);
   registers_reg_24_2_inst : HS65_LH_DFPRQX9 port map( D => n2172, CP => clk, 
                           RN => n6590, Q => registers_24_2_port);
   registers_reg_24_1_inst : HS65_LH_DFPRQX9 port map( D => n2171, CP => clk, 
                           RN => n6590, Q => registers_24_1_port);
   registers_reg_24_0_inst : HS65_LH_DFPRQX9 port map( D => n2170, CP => clk, 
                           RN => n6590, Q => registers_24_0_port);
   registers_reg_23_31_inst : HS65_LH_DFPRQX9 port map( D => n2169, CP => clk, 
                           RN => n6593, Q => registers_23_31_port);
   registers_reg_23_30_inst : HS65_LH_DFPRQX9 port map( D => n2168, CP => clk, 
                           RN => n6593, Q => registers_23_30_port);
   registers_reg_23_29_inst : HS65_LH_DFPRQX9 port map( D => n2167, CP => clk, 
                           RN => n6593, Q => registers_23_29_port);
   registers_reg_23_28_inst : HS65_LH_DFPRQX9 port map( D => n2166, CP => clk, 
                           RN => n6593, Q => registers_23_28_port);
   registers_reg_23_27_inst : HS65_LH_DFPRQX9 port map( D => n2165, CP => clk, 
                           RN => n6594, Q => registers_23_27_port);
   registers_reg_23_26_inst : HS65_LH_DFPRQX9 port map( D => n2164, CP => clk, 
                           RN => n6594, Q => registers_23_26_port);
   registers_reg_23_25_inst : HS65_LH_DFPRQX9 port map( D => n2163, CP => clk, 
                           RN => n6594, Q => registers_23_25_port);
   registers_reg_23_24_inst : HS65_LH_DFPRQX9 port map( D => n2162, CP => clk, 
                           RN => n6594, Q => registers_23_24_port);
   registers_reg_23_23_inst : HS65_LH_DFPRQX9 port map( D => n2161, CP => clk, 
                           RN => n6592, Q => registers_23_23_port);
   registers_reg_23_22_inst : HS65_LH_DFPRQX9 port map( D => n2160, CP => clk, 
                           RN => n6595, Q => registers_23_22_port);
   registers_reg_23_21_inst : HS65_LH_DFPRQX9 port map( D => n2159, CP => clk, 
                           RN => n6595, Q => registers_23_21_port);
   registers_reg_23_20_inst : HS65_LH_DFPRQX9 port map( D => n2158, CP => clk, 
                           RN => n6593, Q => registers_23_20_port);
   registers_reg_23_19_inst : HS65_LH_DFPRQX9 port map( D => n2157, CP => clk, 
                           RN => n6593, Q => registers_23_19_port);
   registers_reg_23_18_inst : HS65_LH_DFPRQX9 port map( D => n2156, CP => clk, 
                           RN => n6592, Q => registers_23_18_port);
   registers_reg_23_17_inst : HS65_LH_DFPRQX9 port map( D => n2155, CP => clk, 
                           RN => n6592, Q => registers_23_17_port);
   registers_reg_23_16_inst : HS65_LH_DFPRQX9 port map( D => n2154, CP => clk, 
                           RN => n6592, Q => registers_23_16_port);
   registers_reg_23_15_inst : HS65_LH_DFPRQX9 port map( D => n2153, CP => clk, 
                           RN => n6592, Q => registers_23_15_port);
   registers_reg_23_14_inst : HS65_LH_DFPRQX9 port map( D => n2152, CP => clk, 
                           RN => n6592, Q => registers_23_14_port);
   registers_reg_23_13_inst : HS65_LH_DFPRQX9 port map( D => n2151, CP => clk, 
                           RN => n6592, Q => registers_23_13_port);
   registers_reg_23_12_inst : HS65_LH_DFPRQX9 port map( D => n2150, CP => clk, 
                           RN => n6592, Q => registers_23_12_port);
   registers_reg_23_11_inst : HS65_LH_DFPRQX9 port map( D => n2149, CP => clk, 
                           RN => n6592, Q => registers_23_11_port);
   registers_reg_23_10_inst : HS65_LH_DFPRQX9 port map( D => n2148, CP => clk, 
                           RN => n6593, Q => registers_23_10_port);
   registers_reg_23_9_inst : HS65_LH_DFPRQX9 port map( D => n2147, CP => clk, 
                           RN => n6593, Q => registers_23_9_port);
   registers_reg_23_8_inst : HS65_LH_DFPRQX9 port map( D => n2146, CP => clk, 
                           RN => n6593, Q => registers_23_8_port);
   registers_reg_23_7_inst : HS65_LH_DFPRQX9 port map( D => n2145, CP => clk, 
                           RN => n6591, Q => registers_23_7_port);
   registers_reg_23_6_inst : HS65_LH_DFPRQX9 port map( D => n2144, CP => clk, 
                           RN => n6591, Q => registers_23_6_port);
   registers_reg_23_5_inst : HS65_LH_DFPRQX9 port map( D => n2143, CP => clk, 
                           RN => n6591, Q => registers_23_5_port);
   registers_reg_23_4_inst : HS65_LH_DFPRQX9 port map( D => n2142, CP => clk, 
                           RN => n6591, Q => registers_23_4_port);
   registers_reg_23_3_inst : HS65_LH_DFPRQX9 port map( D => n2141, CP => clk, 
                           RN => n6591, Q => registers_23_3_port);
   registers_reg_23_2_inst : HS65_LH_DFPRQX9 port map( D => n2140, CP => clk, 
                           RN => n6591, Q => registers_23_2_port);
   registers_reg_23_1_inst : HS65_LH_DFPRQX9 port map( D => n2139, CP => clk, 
                           RN => n6591, Q => registers_23_1_port);
   registers_reg_23_0_inst : HS65_LH_DFPRQX9 port map( D => n2138, CP => clk, 
                           RN => n6591, Q => registers_23_0_port);
   registers_reg_22_31_inst : HS65_LH_DFPRQX9 port map( D => n2137, CP => clk, 
                           RN => n6596, Q => registers_22_31_port);
   registers_reg_22_30_inst : HS65_LH_DFPRQX9 port map( D => n2136, CP => clk, 
                           RN => n6597, Q => registers_22_30_port);
   registers_reg_22_29_inst : HS65_LH_DFPRQX9 port map( D => n2135, CP => clk, 
                           RN => n6597, Q => registers_22_29_port);
   registers_reg_22_28_inst : HS65_LH_DFPRQX9 port map( D => n2134, CP => clk, 
                           RN => n6597, Q => registers_22_28_port);
   registers_reg_22_27_inst : HS65_LH_DFPRQX9 port map( D => n2133, CP => clk, 
                           RN => n6597, Q => registers_22_27_port);
   registers_reg_22_26_inst : HS65_LH_DFPRQX9 port map( D => n2132, CP => clk, 
                           RN => n6596, Q => registers_22_26_port);
   registers_reg_22_25_inst : HS65_LH_DFPRQX9 port map( D => n2131, CP => clk, 
                           RN => n6596, Q => registers_22_25_port);
   registers_reg_22_24_inst : HS65_LH_DFPRQX9 port map( D => n2130, CP => clk, 
                           RN => n6596, Q => registers_22_24_port);
   registers_reg_22_23_inst : HS65_LH_DFPRQX9 port map( D => n2129, CP => clk, 
                           RN => n6595, Q => registers_22_23_port);
   registers_reg_22_22_inst : HS65_LH_DFPRQX9 port map( D => n2128, CP => clk, 
                           RN => n6595, Q => registers_22_22_port);
   registers_reg_22_21_inst : HS65_LH_DFPRQX9 port map( D => n2127, CP => clk, 
                           RN => n6593, Q => registers_22_21_port);
   registers_reg_22_20_inst : HS65_LH_DFPRQX9 port map( D => n2126, CP => clk, 
                           RN => n6593, Q => registers_22_20_port);
   registers_reg_22_19_inst : HS65_LH_DFPRQX9 port map( D => n2125, CP => clk, 
                           RN => n6593, Q => registers_22_19_port);
   registers_reg_22_18_inst : HS65_LH_DFPRQX9 port map( D => n2124, CP => clk, 
                           RN => n6597, Q => registers_22_18_port);
   registers_reg_22_17_inst : HS65_LH_DFPRQX9 port map( D => n2123, CP => clk, 
                           RN => n6597, Q => registers_22_17_port);
   registers_reg_22_16_inst : HS65_LH_DFPRQX9 port map( D => n2122, CP => clk, 
                           RN => n6597, Q => registers_22_16_port);
   registers_reg_22_15_inst : HS65_LH_DFPRQX9 port map( D => n2121, CP => clk, 
                           RN => n6594, Q => registers_22_15_port);
   registers_reg_22_14_inst : HS65_LH_DFPRQX9 port map( D => n2120, CP => clk, 
                           RN => n6594, Q => registers_22_14_port);
   registers_reg_22_13_inst : HS65_LH_DFPRQX9 port map( D => n2119, CP => clk, 
                           RN => n6594, Q => registers_22_13_port);
   registers_reg_22_12_inst : HS65_LH_DFPRQX9 port map( D => n2118, CP => clk, 
                           RN => n6594, Q => registers_22_12_port);
   registers_reg_22_11_inst : HS65_LH_DFPRQX9 port map( D => n2117, CP => clk, 
                           RN => n6594, Q => registers_22_11_port);
   registers_reg_22_10_inst : HS65_LH_DFPRQX9 port map( D => n2116, CP => clk, 
                           RN => n6594, Q => registers_22_10_port);
   registers_reg_22_9_inst : HS65_LH_DFPRQX9 port map( D => n2115, CP => clk, 
                           RN => n6594, Q => registers_22_9_port);
   registers_reg_22_8_inst : HS65_LH_DFPRQX9 port map( D => n2114, CP => clk, 
                           RN => n6594, Q => registers_22_8_port);
   registers_reg_22_7_inst : HS65_LH_DFPRQX9 port map( D => n2113, CP => clk, 
                           RN => n6586, Q => registers_22_7_port);
   registers_reg_22_6_inst : HS65_LH_DFPRQX9 port map( D => n2112, CP => clk, 
                           RN => n6538, Q => registers_22_6_port);
   registers_reg_22_5_inst : HS65_LH_DFPRQX9 port map( D => n2111, CP => clk, 
                           RN => n6538, Q => registers_22_5_port);
   registers_reg_22_4_inst : HS65_LH_DFPRQX9 port map( D => n2110, CP => clk, 
                           RN => n6538, Q => registers_22_4_port);
   registers_reg_22_3_inst : HS65_LH_DFPRQX9 port map( D => n2109, CP => clk, 
                           RN => n6538, Q => registers_22_3_port);
   registers_reg_22_2_inst : HS65_LH_DFPRQX9 port map( D => n2108, CP => clk, 
                           RN => n6538, Q => registers_22_2_port);
   registers_reg_22_1_inst : HS65_LH_DFPRQX9 port map( D => n2107, CP => clk, 
                           RN => n6538, Q => registers_22_1_port);
   registers_reg_22_0_inst : HS65_LH_DFPRQX9 port map( D => n2106, CP => clk, 
                           RN => n6538, Q => registers_22_0_port);
   registers_reg_21_31_inst : HS65_LH_DFPRQX9 port map( D => n2105, CP => clk, 
                           RN => n6541, Q => registers_21_31_port);
   registers_reg_21_30_inst : HS65_LH_DFPRQX9 port map( D => n2104, CP => clk, 
                           RN => n6542, Q => registers_21_30_port);
   registers_reg_21_29_inst : HS65_LH_DFPRQX9 port map( D => n2103, CP => clk, 
                           RN => n6541, Q => registers_21_29_port);
   registers_reg_21_28_inst : HS65_LH_DFPRQX9 port map( D => n2102, CP => clk, 
                           RN => n6542, Q => registers_21_28_port);
   registers_reg_21_27_inst : HS65_LH_DFPRQX9 port map( D => n2101, CP => clk, 
                           RN => n6541, Q => registers_21_27_port);
   registers_reg_21_26_inst : HS65_LH_DFPRQX9 port map( D => n2100, CP => clk, 
                           RN => n6540, Q => registers_21_26_port);
   registers_reg_21_25_inst : HS65_LH_DFPRQX9 port map( D => n2099, CP => clk, 
                           RN => n6540, Q => registers_21_25_port);
   registers_reg_21_24_inst : HS65_LH_DFPRQX9 port map( D => n2098, CP => clk, 
                           RN => n6539, Q => registers_21_24_port);
   registers_reg_21_23_inst : HS65_LH_DFPRQX9 port map( D => n2097, CP => clk, 
                           RN => n6539, Q => registers_21_23_port);
   registers_reg_21_22_inst : HS65_LH_DFPRQX9 port map( D => n2096, CP => clk, 
                           RN => n6573, Q => registers_21_22_port);
   registers_reg_21_21_inst : HS65_LH_DFPRQX9 port map( D => n2095, CP => clk, 
                           RN => n6573, Q => registers_21_21_port);
   registers_reg_21_20_inst : HS65_LH_DFPRQX9 port map( D => n2094, CP => clk, 
                           RN => n6572, Q => registers_21_20_port);
   registers_reg_21_19_inst : HS65_LH_DFPRQX9 port map( D => n2093, CP => clk, 
                           RN => n6572, Q => registers_21_19_port);
   registers_reg_21_18_inst : HS65_LH_DFPRQX9 port map( D => n2092, CP => clk, 
                           RN => n6569, Q => registers_21_18_port);
   registers_reg_21_17_inst : HS65_LH_DFPRQX9 port map( D => n2091, CP => clk, 
                           RN => n6569, Q => registers_21_17_port);
   registers_reg_21_16_inst : HS65_LH_DFPRQX9 port map( D => n2090, CP => clk, 
                           RN => n6569, Q => registers_21_16_port);
   registers_reg_21_15_inst : HS65_LH_DFPRQX9 port map( D => n2089, CP => clk, 
                           RN => n6569, Q => registers_21_15_port);
   registers_reg_21_14_inst : HS65_LH_DFPRQX9 port map( D => n2088, CP => clk, 
                           RN => n6569, Q => registers_21_14_port);
   registers_reg_21_13_inst : HS65_LH_DFPRQX9 port map( D => n2087, CP => clk, 
                           RN => n6569, Q => registers_21_13_port);
   registers_reg_21_12_inst : HS65_LH_DFPRQX9 port map( D => n2086, CP => clk, 
                           RN => n6569, Q => registers_21_12_port);
   registers_reg_21_11_inst : HS65_LH_DFPRQX9 port map( D => n2085, CP => clk, 
                           RN => n6569, Q => registers_21_11_port);
   registers_reg_21_10_inst : HS65_LH_DFPRQX9 port map( D => n2084, CP => clk, 
                           RN => n6572, Q => registers_21_10_port);
   registers_reg_21_9_inst : HS65_LH_DFPRQX9 port map( D => n2083, CP => clk, 
                           RN => n6572, Q => registers_21_9_port);
   registers_reg_21_8_inst : HS65_LH_DFPRQX9 port map( D => n2082, CP => clk, 
                           RN => n6572, Q => registers_21_8_port);
   registers_reg_21_7_inst : HS65_LH_DFPRQX9 port map( D => n2081, CP => clk, 
                           RN => n6570, Q => registers_21_7_port);
   registers_reg_21_6_inst : HS65_LH_DFPRQX9 port map( D => n2080, CP => clk, 
                           RN => n6570, Q => registers_21_6_port);
   registers_reg_21_5_inst : HS65_LH_DFPRQX9 port map( D => n2079, CP => clk, 
                           RN => n6570, Q => registers_21_5_port);
   registers_reg_21_4_inst : HS65_LH_DFPRQX9 port map( D => n2078, CP => clk, 
                           RN => n6570, Q => registers_21_4_port);
   registers_reg_21_3_inst : HS65_LH_DFPRQX9 port map( D => n2077, CP => clk, 
                           RN => n6570, Q => registers_21_3_port);
   registers_reg_21_2_inst : HS65_LH_DFPRQX9 port map( D => n2076, CP => clk, 
                           RN => n6570, Q => registers_21_2_port);
   registers_reg_21_1_inst : HS65_LH_DFPRQX9 port map( D => n2075, CP => clk, 
                           RN => n6570, Q => registers_21_1_port);
   registers_reg_21_0_inst : HS65_LH_DFPRQX9 port map( D => n2074, CP => clk, 
                           RN => n6570, Q => registers_21_0_port);
   registers_reg_20_31_inst : HS65_LH_DFPRQX9 port map( D => n2073, CP => clk, 
                           RN => n6574, Q => registers_20_31_port);
   registers_reg_20_30_inst : HS65_LH_DFPRQX9 port map( D => n2072, CP => clk, 
                           RN => n6571, Q => registers_20_30_port);
   registers_reg_20_29_inst : HS65_LH_DFPRQX9 port map( D => n2071, CP => clk, 
                           RN => n6571, Q => registers_20_29_port);
   registers_reg_20_28_inst : HS65_LH_DFPRQX9 port map( D => n2070, CP => clk, 
                           RN => n6571, Q => registers_20_28_port);
   registers_reg_20_27_inst : HS65_LH_DFPRQX9 port map( D => n2069, CP => clk, 
                           RN => n6570, Q => registers_20_27_port);
   registers_reg_20_26_inst : HS65_LH_DFPRQX9 port map( D => n2068, CP => clk, 
                           RN => n6570, Q => registers_20_26_port);
   registers_reg_20_25_inst : HS65_LH_DFPRQX9 port map( D => n2067, CP => clk, 
                           RN => n6569, Q => registers_20_25_port);
   registers_reg_20_24_inst : HS65_LH_DFPRQX9 port map( D => n2066, CP => clk, 
                           RN => n6569, Q => registers_20_24_port);
   registers_reg_20_23_inst : HS65_LH_DFPRQX9 port map( D => n2065, CP => clk, 
                           RN => n6574, Q => registers_20_23_port);
   registers_reg_20_22_inst : HS65_LH_DFPRQX9 port map( D => n2064, CP => clk, 
                           RN => n6574, Q => registers_20_22_port);
   registers_reg_20_21_inst : HS65_LH_DFPRQX9 port map( D => n2063, CP => clk, 
                           RN => n6573, Q => registers_20_21_port);
   registers_reg_20_20_inst : HS65_LH_DFPRQX9 port map( D => n2062, CP => clk, 
                           RN => n6574, Q => registers_20_20_port);
   registers_reg_20_19_inst : HS65_LH_DFPRQX9 port map( D => n2061, CP => clk, 
                           RN => n6574, Q => registers_20_19_port);
   registers_reg_20_18_inst : HS65_LH_DFPRQX9 port map( D => n2060, CP => clk, 
                           RN => n6573, Q => registers_20_18_port);
   registers_reg_20_17_inst : HS65_LH_DFPRQX9 port map( D => n2059, CP => clk, 
                           RN => n6573, Q => registers_20_17_port);
   registers_reg_20_16_inst : HS65_LH_DFPRQX9 port map( D => n2058, CP => clk, 
                           RN => n6573, Q => registers_20_16_port);
   registers_reg_20_15_inst : HS65_LH_DFPRQX9 port map( D => n2057, CP => clk, 
                           RN => n6573, Q => registers_20_15_port);
   registers_reg_20_14_inst : HS65_LH_DFPRQX9 port map( D => n2056, CP => clk, 
                           RN => n6573, Q => registers_20_14_port);
   registers_reg_20_13_inst : HS65_LH_DFPRQX9 port map( D => n2055, CP => clk, 
                           RN => n6573, Q => registers_20_13_port);
   registers_reg_20_12_inst : HS65_LH_DFPRQX9 port map( D => n2054, CP => clk, 
                           RN => n6573, Q => registers_20_12_port);
   registers_reg_20_11_inst : HS65_LH_DFPRQX9 port map( D => n2053, CP => clk, 
                           RN => n6573, Q => registers_20_11_port);
   registers_reg_20_10_inst : HS65_LH_DFPRQX9 port map( D => n2052, CP => clk, 
                           RN => n6574, Q => registers_20_10_port);
   registers_reg_20_9_inst : HS65_LH_DFPRQX9 port map( D => n2051, CP => clk, 
                           RN => n6574, Q => registers_20_9_port);
   registers_reg_20_8_inst : HS65_LH_DFPRQX9 port map( D => n2050, CP => clk, 
                           RN => n6574, Q => registers_20_8_port);
   registers_reg_20_7_inst : HS65_LH_DFPRQX9 port map( D => n2049, CP => clk, 
                           RN => n6576, Q => registers_20_7_port);
   registers_reg_20_6_inst : HS65_LH_DFPRQX9 port map( D => n2048, CP => clk, 
                           RN => n6576, Q => registers_20_6_port);
   registers_reg_20_5_inst : HS65_LH_DFPRQX9 port map( D => n2047, CP => clk, 
                           RN => n6576, Q => registers_20_5_port);
   registers_reg_20_4_inst : HS65_LH_DFPRQX9 port map( D => n2046, CP => clk, 
                           RN => n6576, Q => registers_20_4_port);
   registers_reg_20_3_inst : HS65_LH_DFPRQX9 port map( D => n2045, CP => clk, 
                           RN => n6576, Q => registers_20_3_port);
   registers_reg_20_2_inst : HS65_LH_DFPRQX9 port map( D => n2044, CP => clk, 
                           RN => n6576, Q => registers_20_2_port);
   registers_reg_20_1_inst : HS65_LH_DFPRQX9 port map( D => n2043, CP => clk, 
                           RN => n6576, Q => registers_20_1_port);
   registers_reg_20_0_inst : HS65_LH_DFPRQX9 port map( D => n2042, CP => clk, 
                           RN => n6576, Q => registers_20_0_port);
   registers_reg_19_31_inst : HS65_LH_DFPRQX9 port map( D => n2041, CP => clk, 
                           RN => n6588, Q => registers_19_31_port);
   registers_reg_19_30_inst : HS65_LH_DFPRQX9 port map( D => n2040, CP => clk, 
                           RN => n6588, Q => registers_19_30_port);
   registers_reg_19_29_inst : HS65_LH_DFPRQX9 port map( D => n2039, CP => clk, 
                           RN => n6588, Q => registers_19_29_port);
   registers_reg_19_28_inst : HS65_LH_DFPRQX9 port map( D => n2038, CP => clk, 
                           RN => n6588, Q => registers_19_28_port);
   registers_reg_19_27_inst : HS65_LH_DFPRQX9 port map( D => n2037, CP => clk, 
                           RN => n6578, Q => registers_19_27_port);
   registers_reg_19_26_inst : HS65_LH_DFPRQX9 port map( D => n2036, CP => clk, 
                           RN => n6577, Q => registers_19_26_port);
   registers_reg_19_25_inst : HS65_LH_DFPRQX9 port map( D => n2035, CP => clk, 
                           RN => n6577, Q => registers_19_25_port);
   registers_reg_19_24_inst : HS65_LH_DFPRQX9 port map( D => n2034, CP => clk, 
                           RN => n6577, Q => registers_19_24_port);
   registers_reg_19_23_inst : HS65_LH_DFPRQX9 port map( D => n2033, CP => clk, 
                           RN => n6577, Q => registers_19_23_port);
   registers_reg_19_22_inst : HS65_LH_DFPRQX9 port map( D => n2032, CP => clk, 
                           RN => n6577, Q => registers_19_22_port);
   registers_reg_19_21_inst : HS65_LH_DFPRQX9 port map( D => n2031, CP => clk, 
                           RN => n6577, Q => registers_19_21_port);
   registers_reg_19_20_inst : HS65_LH_DFPRQX9 port map( D => n2030, CP => clk, 
                           RN => n6577, Q => registers_19_20_port);
   registers_reg_19_19_inst : HS65_LH_DFPRQX9 port map( D => n2029, CP => clk, 
                           RN => n6587, Q => registers_19_19_port);
   registers_reg_19_18_inst : HS65_LH_DFPRQX9 port map( D => n2028, CP => clk, 
                           RN => n6587, Q => registers_19_18_port);
   registers_reg_19_17_inst : HS65_LH_DFPRQX9 port map( D => n2027, CP => clk, 
                           RN => n6587, Q => registers_19_17_port);
   registers_reg_19_16_inst : HS65_LH_DFPRQX9 port map( D => n2026, CP => clk, 
                           RN => n6587, Q => registers_19_16_port);
   registers_reg_19_15_inst : HS65_LH_DFPRQX9 port map( D => n2025, CP => clk, 
                           RN => n6587, Q => registers_19_15_port);
   registers_reg_19_14_inst : HS65_LH_DFPRQX9 port map( D => n2024, CP => clk, 
                           RN => n6587, Q => registers_19_14_port);
   registers_reg_19_13_inst : HS65_LH_DFPRQX9 port map( D => n2023, CP => clk, 
                           RN => n6587, Q => registers_19_13_port);
   registers_reg_19_12_inst : HS65_LH_DFPRQX9 port map( D => n2022, CP => clk, 
                           RN => n6587, Q => registers_19_12_port);
   registers_reg_19_11_inst : HS65_LH_DFPRQX9 port map( D => n2021, CP => clk, 
                           RN => n6587, Q => registers_19_11_port);
   registers_reg_19_10_inst : HS65_LH_DFPRQX9 port map( D => n2020, CP => clk, 
                           RN => n6587, Q => registers_19_10_port);
   registers_reg_19_9_inst : HS65_LH_DFPRQX9 port map( D => n2019, CP => clk, 
                           RN => n6587, Q => registers_19_9_port);
   registers_reg_19_8_inst : HS65_LH_DFPRQX9 port map( D => n2018, CP => clk, 
                           RN => n6587, Q => registers_19_8_port);
   registers_reg_19_7_inst : HS65_LH_DFPRQX9 port map( D => n2017, CP => clk, 
                           RN => n6571, Q => registers_19_7_port);
   registers_reg_19_6_inst : HS65_LH_DFPRQX9 port map( D => n2016, CP => clk, 
                           RN => n6571, Q => registers_19_6_port);
   registers_reg_19_5_inst : HS65_LH_DFPRQX9 port map( D => n2015, CP => clk, 
                           RN => n6571, Q => registers_19_5_port);
   registers_reg_19_4_inst : HS65_LH_DFPRQX9 port map( D => n2014, CP => clk, 
                           RN => n6571, Q => registers_19_4_port);
   registers_reg_19_3_inst : HS65_LH_DFPRQX9 port map( D => n2013, CP => clk, 
                           RN => n6571, Q => registers_19_3_port);
   registers_reg_19_2_inst : HS65_LH_DFPRQX9 port map( D => n2012, CP => clk, 
                           RN => n6571, Q => registers_19_2_port);
   registers_reg_19_1_inst : HS65_LH_DFPRQX9 port map( D => n2011, CP => clk, 
                           RN => n6571, Q => registers_19_1_port);
   registers_reg_19_0_inst : HS65_LH_DFPRQX9 port map( D => n2010, CP => clk, 
                           RN => n6571, Q => registers_19_0_port);
   registers_reg_18_31_inst : HS65_LH_DFPRQX9 port map( D => n2009, CP => clk, 
                           RN => n6577, Q => registers_18_31_port);
   registers_reg_18_30_inst : HS65_LH_DFPRQX9 port map( D => n2008, CP => clk, 
                           RN => n6577, Q => registers_18_30_port);
   registers_reg_18_29_inst : HS65_LH_DFPRQX9 port map( D => n2007, CP => clk, 
                           RN => n6577, Q => registers_18_29_port);
   registers_reg_18_28_inst : HS65_LH_DFPRQX9 port map( D => n2006, CP => clk, 
                           RN => n6578, Q => registers_18_28_port);
   registers_reg_18_27_inst : HS65_LH_DFPRQX9 port map( D => n2005, CP => clk, 
                           RN => n6578, Q => registers_18_27_port);
   registers_reg_18_26_inst : HS65_LH_DFPRQX9 port map( D => n2004, CP => clk, 
                           RN => n6578, Q => registers_18_26_port);
   registers_reg_18_25_inst : HS65_LH_DFPRQX9 port map( D => n2003, CP => clk, 
                           RN => n6577, Q => registers_18_25_port);
   registers_reg_18_24_inst : HS65_LH_DFPRQX9 port map( D => n2002, CP => clk, 
                           RN => n6577, Q => registers_18_24_port);
   registers_reg_18_23_inst : HS65_LH_DFPRQX9 port map( D => n2001, CP => clk, 
                           RN => n6574, Q => registers_18_23_port);
   registers_reg_18_22_inst : HS65_LH_DFPRQX9 port map( D => n2000, CP => clk, 
                           RN => n6574, Q => registers_18_22_port);
   registers_reg_18_21_inst : HS65_LH_DFPRQX9 port map( D => n1999, CP => clk, 
                           RN => n6574, Q => registers_18_21_port);
   registers_reg_18_20_inst : HS65_LH_DFPRQX9 port map( D => n1998, CP => clk, 
                           RN => n6573, Q => registers_18_20_port);
   registers_reg_18_19_inst : HS65_LH_DFPRQX9 port map( D => n1997, CP => clk, 
                           RN => n6572, Q => registers_18_19_port);
   registers_reg_18_18_inst : HS65_LH_DFPRQX9 port map( D => n1996, CP => clk, 
                           RN => n6572, Q => registers_18_18_port);
   registers_reg_18_17_inst : HS65_LH_DFPRQX9 port map( D => n1995, CP => clk, 
                           RN => n6572, Q => registers_18_17_port);
   registers_reg_18_16_inst : HS65_LH_DFPRQX9 port map( D => n1994, CP => clk, 
                           RN => n6574, Q => registers_18_16_port);
   registers_reg_18_15_inst : HS65_LH_DFPRQX9 port map( D => n1993, CP => clk, 
                           RN => n6548, Q => registers_18_15_port);
   registers_reg_18_14_inst : HS65_LH_DFPRQX9 port map( D => n1992, CP => clk, 
                           RN => n6550, Q => registers_18_14_port);
   registers_reg_18_13_inst : HS65_LH_DFPRQX9 port map( D => n1991, CP => clk, 
                           RN => n6540, Q => registers_18_13_port);
   registers_reg_18_12_inst : HS65_LH_DFPRQX9 port map( D => n1990, CP => clk, 
                           RN => n6540, Q => registers_18_12_port);
   registers_reg_18_11_inst : HS65_LH_DFPRQX9 port map( D => n1989, CP => clk, 
                           RN => n6540, Q => registers_18_11_port);
   registers_reg_18_10_inst : HS65_LH_DFPRQX9 port map( D => n1988, CP => clk, 
                           RN => n6542, Q => registers_18_10_port);
   registers_reg_18_9_inst : HS65_LH_DFPRQX9 port map( D => n1987, CP => clk, 
                           RN => n6542, Q => registers_18_9_port);
   registers_reg_18_8_inst : HS65_LH_DFPRQX9 port map( D => n1986, CP => clk, 
                           RN => n6542, Q => registers_18_8_port);
   registers_reg_18_7_inst : HS65_LH_DFPRQX9 port map( D => n1985, CP => clk, 
                           RN => n6542, Q => registers_18_7_port);
   registers_reg_18_6_inst : HS65_LH_DFPRQX9 port map( D => n1984, CP => clk, 
                           RN => n6542, Q => registers_18_6_port);
   registers_reg_18_5_inst : HS65_LH_DFPRQX9 port map( D => n1983, CP => clk, 
                           RN => n6542, Q => registers_18_5_port);
   registers_reg_18_4_inst : HS65_LH_DFPRQX9 port map( D => n1982, CP => clk, 
                           RN => n6542, Q => registers_18_4_port);
   registers_reg_18_3_inst : HS65_LH_DFPRQX9 port map( D => n1981, CP => clk, 
                           RN => n6542, Q => registers_18_3_port);
   registers_reg_18_2_inst : HS65_LH_DFPRQX9 port map( D => n1980, CP => clk, 
                           RN => n6552, Q => registers_18_2_port);
   registers_reg_18_1_inst : HS65_LH_DFPRQX9 port map( D => n1979, CP => clk, 
                           RN => n6552, Q => registers_18_1_port);
   registers_reg_18_0_inst : HS65_LH_DFPRQX9 port map( D => n1978, CP => clk, 
                           RN => n6552, Q => registers_18_0_port);
   registers_reg_17_31_inst : HS65_LH_DFPRQX9 port map( D => n1977, CP => clk, 
                           RN => n6555, Q => registers_17_31_port);
   registers_reg_17_30_inst : HS65_LH_DFPRQX9 port map( D => n1976, CP => clk, 
                           RN => n6555, Q => registers_17_30_port);
   registers_reg_17_29_inst : HS65_LH_DFPRQX9 port map( D => n1975, CP => clk, 
                           RN => n6555, Q => registers_17_29_port);
   registers_reg_17_28_inst : HS65_LH_DFPRQX9 port map( D => n1974, CP => clk, 
                           RN => n6555, Q => registers_17_28_port);
   registers_reg_17_27_inst : HS65_LH_DFPRQX9 port map( D => n1973, CP => clk, 
                           RN => n6557, Q => registers_17_27_port);
   registers_reg_17_26_inst : HS65_LH_DFPRQX9 port map( D => n1972, CP => clk, 
                           RN => n6557, Q => registers_17_26_port);
   registers_reg_17_25_inst : HS65_LH_DFPRQX9 port map( D => n1971, CP => clk, 
                           RN => n6557, Q => registers_17_25_port);
   registers_reg_17_24_inst : HS65_LH_DFPRQX9 port map( D => n1970, CP => clk, 
                           RN => n6552, Q => registers_17_24_port);
   registers_reg_17_23_inst : HS65_LH_DFPRQX9 port map( D => n1969, CP => clk, 
                           RN => n6552, Q => registers_17_23_port);
   registers_reg_17_22_inst : HS65_LH_DFPRQX9 port map( D => n1968, CP => clk, 
                           RN => n6556, Q => registers_17_22_port);
   registers_reg_17_21_inst : HS65_LH_DFPRQX9 port map( D => n1967, CP => clk, 
                           RN => n6556, Q => registers_17_21_port);
   registers_reg_17_20_inst : HS65_LH_DFPRQX9 port map( D => n1966, CP => clk, 
                           RN => n6556, Q => registers_17_20_port);
   registers_reg_17_19_inst : HS65_LH_DFPRQX9 port map( D => n1965, CP => clk, 
                           RN => n6556, Q => registers_17_19_port);
   registers_reg_17_18_inst : HS65_LH_DFPRQX9 port map( D => n1964, CP => clk, 
                           RN => n6556, Q => registers_17_18_port);
   registers_reg_17_17_inst : HS65_LH_DFPRQX9 port map( D => n1963, CP => clk, 
                           RN => n6556, Q => registers_17_17_port);
   registers_reg_17_16_inst : HS65_LH_DFPRQX9 port map( D => n1962, CP => clk, 
                           RN => n6556, Q => registers_17_16_port);
   registers_reg_17_15_inst : HS65_LH_DFPRQX9 port map( D => n1961, CP => clk, 
                           RN => n6556, Q => registers_17_15_port);
   registers_reg_17_14_inst : HS65_LH_DFPRQX9 port map( D => n1960, CP => clk, 
                           RN => n6556, Q => registers_17_14_port);
   registers_reg_17_13_inst : HS65_LH_DFPRQX9 port map( D => n1959, CP => clk, 
                           RN => n6556, Q => registers_17_13_port);
   registers_reg_17_12_inst : HS65_LH_DFPRQX9 port map( D => n1958, CP => clk, 
                           RN => n6556, Q => registers_17_12_port);
   registers_reg_17_11_inst : HS65_LH_DFPRQX9 port map( D => n1957, CP => clk, 
                           RN => n6556, Q => registers_17_11_port);
   registers_reg_17_10_inst : HS65_LH_DFPRQX9 port map( D => n1956, CP => clk, 
                           RN => n6552, Q => registers_17_10_port);
   registers_reg_17_9_inst : HS65_LH_DFPRQX9 port map( D => n1955, CP => clk, 
                           RN => n6552, Q => registers_17_9_port);
   registers_reg_17_8_inst : HS65_LH_DFPRQX9 port map( D => n1954, CP => clk, 
                           RN => n6552, Q => registers_17_8_port);
   registers_reg_17_7_inst : HS65_LH_DFPRQX9 port map( D => n1953, CP => clk, 
                           RN => n6555, Q => registers_17_7_port);
   registers_reg_17_6_inst : HS65_LH_DFPRQX9 port map( D => n1952, CP => clk, 
                           RN => n6555, Q => registers_17_6_port);
   registers_reg_17_5_inst : HS65_LH_DFPRQX9 port map( D => n1951, CP => clk, 
                           RN => n6555, Q => registers_17_5_port);
   registers_reg_17_4_inst : HS65_LH_DFPRQX9 port map( D => n1950, CP => clk, 
                           RN => n6555, Q => registers_17_4_port);
   registers_reg_17_3_inst : HS65_LH_DFPRQX9 port map( D => n1949, CP => clk, 
                           RN => n6555, Q => registers_17_3_port);
   registers_reg_17_2_inst : HS65_LH_DFPRQX9 port map( D => n1948, CP => clk, 
                           RN => n6555, Q => registers_17_2_port);
   registers_reg_17_1_inst : HS65_LH_DFPRQX9 port map( D => n1947, CP => clk, 
                           RN => n6555, Q => registers_17_1_port);
   registers_reg_17_0_inst : HS65_LH_DFPRQX9 port map( D => n1946, CP => clk, 
                           RN => n6555, Q => registers_17_0_port);
   registers_reg_16_31_inst : HS65_LH_DFPRQX9 port map( D => n1945, CP => clk, 
                           RN => n6557, Q => registers_16_31_port);
   registers_reg_16_30_inst : HS65_LH_DFPRQX9 port map( D => n1944, CP => clk, 
                           RN => n6558, Q => registers_16_30_port);
   registers_reg_16_29_inst : HS65_LH_DFPRQX9 port map( D => n1943, CP => clk, 
                           RN => n6558, Q => registers_16_29_port);
   registers_reg_16_28_inst : HS65_LH_DFPRQX9 port map( D => n1942, CP => clk, 
                           RN => n6558, Q => registers_16_28_port);
   registers_reg_16_27_inst : HS65_LH_DFPRQX9 port map( D => n1941, CP => clk, 
                           RN => n6558, Q => registers_16_27_port);
   registers_reg_16_26_inst : HS65_LH_DFPRQX9 port map( D => n1940, CP => clk, 
                           RN => n6553, Q => registers_16_26_port);
   registers_reg_16_25_inst : HS65_LH_DFPRQX9 port map( D => n1939, CP => clk, 
                           RN => n6553, Q => registers_16_25_port);
   registers_reg_16_24_inst : HS65_LH_DFPRQX9 port map( D => n1938, CP => clk, 
                           RN => n6550, Q => registers_16_24_port);
   registers_reg_16_23_inst : HS65_LH_DFPRQX9 port map( D => n1937, CP => clk, 
                           RN => n6550, Q => registers_16_23_port);
   registers_reg_16_22_inst : HS65_LH_DFPRQX9 port map( D => n1936, CP => clk, 
                           RN => n6550, Q => registers_16_22_port);
   registers_reg_16_21_inst : HS65_LH_DFPRQX9 port map( D => n1935, CP => clk, 
                           RN => n6550, Q => registers_16_21_port);
   registers_reg_16_20_inst : HS65_LH_DFPRQX9 port map( D => n1934, CP => clk, 
                           RN => n6550, Q => registers_16_20_port);
   registers_reg_16_19_inst : HS65_LH_DFPRQX9 port map( D => n1933, CP => clk, 
                           RN => n6557, Q => registers_16_19_port);
   registers_reg_16_18_inst : HS65_LH_DFPRQX9 port map( D => n1932, CP => clk, 
                           RN => n6557, Q => registers_16_18_port);
   registers_reg_16_17_inst : HS65_LH_DFPRQX9 port map( D => n1931, CP => clk, 
                           RN => n6557, Q => registers_16_17_port);
   registers_reg_16_16_inst : HS65_LH_DFPRQX9 port map( D => n1930, CP => clk, 
                           RN => n6557, Q => registers_16_16_port);
   registers_reg_16_15_inst : HS65_LH_DFPRQX9 port map( D => n1929, CP => clk, 
                           RN => n6553, Q => registers_16_15_port);
   registers_reg_16_14_inst : HS65_LH_DFPRQX9 port map( D => n1928, CP => clk, 
                           RN => n6553, Q => registers_16_14_port);
   registers_reg_16_13_inst : HS65_LH_DFPRQX9 port map( D => n1927, CP => clk, 
                           RN => n6553, Q => registers_16_13_port);
   registers_reg_16_12_inst : HS65_LH_DFPRQX9 port map( D => n1926, CP => clk, 
                           RN => n6553, Q => registers_16_12_port);
   registers_reg_16_11_inst : HS65_LH_DFPRQX9 port map( D => n1925, CP => clk, 
                           RN => n6553, Q => registers_16_11_port);
   registers_reg_16_10_inst : HS65_LH_DFPRQX9 port map( D => n1924, CP => clk, 
                           RN => n6553, Q => registers_16_10_port);
   registers_reg_16_9_inst : HS65_LH_DFPRQX9 port map( D => n1923, CP => clk, 
                           RN => n6553, Q => registers_16_9_port);
   registers_reg_16_8_inst : HS65_LH_DFPRQX9 port map( D => n1922, CP => clk, 
                           RN => n6553, Q => registers_16_8_port);
   registers_reg_16_7_inst : HS65_LH_DFPRQX9 port map( D => n1921, CP => clk, 
                           RN => n6554, Q => registers_16_7_port);
   registers_reg_16_6_inst : HS65_LH_DFPRQX9 port map( D => n1920, CP => clk, 
                           RN => n6554, Q => registers_16_6_port);
   registers_reg_16_5_inst : HS65_LH_DFPRQX9 port map( D => n1919, CP => clk, 
                           RN => n6554, Q => registers_16_5_port);
   registers_reg_16_4_inst : HS65_LH_DFPRQX9 port map( D => n1918, CP => clk, 
                           RN => n6554, Q => registers_16_4_port);
   registers_reg_16_3_inst : HS65_LH_DFPRQX9 port map( D => n1917, CP => clk, 
                           RN => n6554, Q => registers_16_3_port);
   registers_reg_16_2_inst : HS65_LH_DFPRQX9 port map( D => n1916, CP => clk, 
                           RN => n6554, Q => registers_16_2_port);
   registers_reg_16_1_inst : HS65_LH_DFPRQX9 port map( D => n1915, CP => clk, 
                           RN => n6554, Q => registers_16_1_port);
   registers_reg_16_0_inst : HS65_LH_DFPRQX9 port map( D => n1914, CP => clk, 
                           RN => n6554, Q => registers_16_0_port);
   registers_reg_13_31_inst : HS65_LH_DFPRQX9 port map( D => n1849, CP => clk, 
                           RN => n6559, Q => registers_13_31_port);
   registers_reg_13_30_inst : HS65_LH_DFPRQX9 port map( D => n1848, CP => clk, 
                           RN => n6559, Q => registers_13_30_port);
   registers_reg_13_29_inst : HS65_LH_DFPRQX9 port map( D => n1847, CP => clk, 
                           RN => n6559, Q => registers_13_29_port);
   registers_reg_13_28_inst : HS65_LH_DFPRQX9 port map( D => n1846, CP => clk, 
                           RN => n6559, Q => registers_13_28_port);
   registers_reg_13_27_inst : HS65_LH_DFPRQX9 port map( D => n1845, CP => clk, 
                           RN => n6561, Q => registers_13_27_port);
   registers_reg_13_26_inst : HS65_LH_DFPRQX9 port map( D => n1844, CP => clk, 
                           RN => n6561, Q => registers_13_26_port);
   registers_reg_13_25_inst : HS65_LH_DFPRQX9 port map( D => n1843, CP => clk, 
                           RN => n6561, Q => registers_13_25_port);
   registers_reg_13_24_inst : HS65_LH_DFPRQX9 port map( D => n1842, CP => clk, 
                           RN => n6561, Q => registers_13_24_port);
   registers_reg_13_23_inst : HS65_LH_DFPRQX9 port map( D => n1841, CP => clk, 
                           RN => n6560, Q => registers_13_23_port);
   registers_reg_13_22_inst : HS65_LH_DFPRQX9 port map( D => n1840, CP => clk, 
                           RN => n6560, Q => registers_13_22_port);
   registers_reg_13_21_inst : HS65_LH_DFPRQX9 port map( D => n1839, CP => clk, 
                           RN => n6560, Q => registers_13_21_port);
   registers_reg_13_20_inst : HS65_LH_DFPRQX9 port map( D => n1838, CP => clk, 
                           RN => n6560, Q => registers_13_20_port);
   registers_reg_13_19_inst : HS65_LH_DFPRQX9 port map( D => n1837, CP => clk, 
                           RN => n6557, Q => registers_13_19_port);
   registers_reg_13_18_inst : HS65_LH_DFPRQX9 port map( D => n1836, CP => clk, 
                           RN => n6557, Q => registers_13_18_port);
   registers_reg_13_17_inst : HS65_LH_DFPRQX9 port map( D => n1835, CP => clk, 
                           RN => n6557, Q => registers_13_17_port);
   registers_reg_13_16_inst : HS65_LH_DFPRQX9 port map( D => n1834, CP => clk, 
                           RN => n6557, Q => registers_13_16_port);
   registers_reg_13_15_inst : HS65_LH_DFPRQX9 port map( D => n1833, CP => clk, 
                           RN => n6562, Q => registers_13_15_port);
   registers_reg_13_14_inst : HS65_LH_DFPRQX9 port map( D => n1832, CP => clk, 
                           RN => n6558, Q => registers_13_14_port);
   registers_reg_13_13_inst : HS65_LH_DFPRQX9 port map( D => n1831, CP => clk, 
                           RN => n6558, Q => registers_13_13_port);
   registers_reg_13_12_inst : HS65_LH_DFPRQX9 port map( D => n1830, CP => clk, 
                           RN => n6558, Q => registers_13_12_port);
   registers_reg_13_11_inst : HS65_LH_DFPRQX9 port map( D => n1829, CP => clk, 
                           RN => n6561, Q => registers_13_11_port);
   registers_reg_13_10_inst : HS65_LH_DFPRQX9 port map( D => n1828, CP => clk, 
                           RN => n6561, Q => registers_13_10_port);
   registers_reg_13_9_inst : HS65_LH_DFPRQX9 port map( D => n1827, CP => clk, 
                           RN => n6561, Q => registers_13_9_port);
   registers_reg_13_8_inst : HS65_LH_DFPRQX9 port map( D => n1826, CP => clk, 
                           RN => n6561, Q => registers_13_8_port);
   registers_reg_13_7_inst : HS65_LH_DFPRQX9 port map( D => n1825, CP => clk, 
                           RN => n6561, Q => registers_13_7_port);
   registers_reg_13_6_inst : HS65_LH_DFPRQX9 port map( D => n1824, CP => clk, 
                           RN => n6561, Q => registers_13_6_port);
   registers_reg_13_5_inst : HS65_LH_DFPRQX9 port map( D => n1823, CP => clk, 
                           RN => n6561, Q => registers_13_5_port);
   registers_reg_13_4_inst : HS65_LH_DFPRQX9 port map( D => n1822, CP => clk, 
                           RN => n6561, Q => registers_13_4_port);
   registers_reg_13_3_inst : HS65_LH_DFPRQX9 port map( D => n1821, CP => clk, 
                           RN => n6541, Q => registers_13_3_port);
   registers_reg_13_2_inst : HS65_LH_DFPRQX9 port map( D => n1820, CP => clk, 
                           RN => n6539, Q => registers_13_2_port);
   registers_reg_13_1_inst : HS65_LH_DFPRQX9 port map( D => n1819, CP => clk, 
                           RN => n6539, Q => registers_13_1_port);
   registers_reg_13_0_inst : HS65_LH_DFPRQX9 port map( D => n1818, CP => clk, 
                           RN => n6539, Q => registers_13_0_port);
   registers_reg_12_31_inst : HS65_LH_DFPRQX9 port map( D => n1817, CP => clk, 
                           RN => n6539, Q => registers_12_31_port);
   registers_reg_12_30_inst : HS65_LH_DFPRQX9 port map( D => n1816, CP => clk, 
                           RN => n6539, Q => registers_12_30_port);
   registers_reg_12_29_inst : HS65_LH_DFPRQX9 port map( D => n1815, CP => clk, 
                           RN => n6539, Q => registers_12_29_port);
   registers_reg_12_28_inst : HS65_LH_DFPRQX9 port map( D => n1814, CP => clk, 
                           RN => n6542, Q => registers_12_28_port);
   registers_reg_12_27_inst : HS65_LH_DFPRQX9 port map( D => n1813, CP => clk, 
                           RN => n6542, Q => registers_12_27_port);
   registers_reg_12_26_inst : HS65_LH_DFPRQX9 port map( D => n1812, CP => clk, 
                           RN => n6541, Q => registers_12_26_port);
   registers_reg_12_25_inst : HS65_LH_DFPRQX9 port map( D => n1811, CP => clk, 
                           RN => n6540, Q => registers_12_25_port);
   registers_reg_12_24_inst : HS65_LH_DFPRQX9 port map( D => n1810, CP => clk, 
                           RN => n6540, Q => registers_12_24_port);
   registers_reg_12_23_inst : HS65_LH_DFPRQX9 port map( D => n1809, CP => clk, 
                           RN => n6539, Q => registers_12_23_port);
   registers_reg_12_22_inst : HS65_LH_DFPRQX9 port map( D => n1808, CP => clk, 
                           RN => n6539, Q => registers_12_22_port);
   registers_reg_12_21_inst : HS65_LH_DFPRQX9 port map( D => n1807, CP => clk, 
                           RN => n6539, Q => registers_12_21_port);
   registers_reg_12_20_inst : HS65_LH_DFPRQX9 port map( D => n1806, CP => clk, 
                           RN => n6538, Q => registers_12_20_port);
   registers_reg_12_19_inst : HS65_LH_DFPRQX9 port map( D => n1805, CP => clk, 
                           RN => n6544, Q => registers_12_19_port);
   registers_reg_12_18_inst : HS65_LH_DFPRQX9 port map( D => n1804, CP => clk, 
                           RN => n6544, Q => registers_12_18_port);
   registers_reg_12_17_inst : HS65_LH_DFPRQX9 port map( D => n1803, CP => clk, 
                           RN => n6544, Q => registers_12_17_port);
   registers_reg_12_16_inst : HS65_LH_DFPRQX9 port map( D => n1802, CP => clk, 
                           RN => n6544, Q => registers_12_16_port);
   registers_reg_12_15_inst : HS65_LH_DFPRQX9 port map( D => n1801, CP => clk, 
                           RN => n6544, Q => registers_12_15_port);
   registers_reg_12_14_inst : HS65_LH_DFPRQX9 port map( D => n1800, CP => clk, 
                           RN => n6544, Q => registers_12_14_port);
   registers_reg_12_13_inst : HS65_LH_DFPRQX9 port map( D => n1799, CP => clk, 
                           RN => n6544, Q => registers_12_13_port);
   registers_reg_12_12_inst : HS65_LH_DFPRQX9 port map( D => n1798, CP => clk, 
                           RN => n6544, Q => registers_12_12_port);
   registers_reg_12_11_inst : HS65_LH_DFPRQX9 port map( D => n1797, CP => clk, 
                           RN => n6545, Q => registers_12_11_port);
   registers_reg_12_10_inst : HS65_LH_DFPRQX9 port map( D => n1796, CP => clk, 
                           RN => n6545, Q => registers_12_10_port);
   registers_reg_12_9_inst : HS65_LH_DFPRQX9 port map( D => n1795, CP => clk, 
                           RN => n6545, Q => registers_12_9_port);
   registers_reg_12_8_inst : HS65_LH_DFPRQX9 port map( D => n1794, CP => clk, 
                           RN => n6545, Q => registers_12_8_port);
   registers_reg_12_7_inst : HS65_LH_DFPRQX9 port map( D => n1793, CP => clk, 
                           RN => n6546, Q => registers_12_7_port);
   registers_reg_12_6_inst : HS65_LH_DFPRQX9 port map( D => n1792, CP => clk, 
                           RN => n6546, Q => registers_12_6_port);
   registers_reg_12_5_inst : HS65_LH_DFPRQX9 port map( D => n1791, CP => clk, 
                           RN => n6546, Q => registers_12_5_port);
   registers_reg_12_4_inst : HS65_LH_DFPRQX9 port map( D => n1790, CP => clk, 
                           RN => n6546, Q => registers_12_4_port);
   registers_reg_12_3_inst : HS65_LH_DFPRQX9 port map( D => n1789, CP => clk, 
                           RN => n6546, Q => registers_12_3_port);
   registers_reg_12_2_inst : HS65_LH_DFPRQX9 port map( D => n1788, CP => clk, 
                           RN => n6546, Q => registers_12_2_port);
   registers_reg_12_1_inst : HS65_LH_DFPRQX9 port map( D => n1787, CP => clk, 
                           RN => n6546, Q => registers_12_1_port);
   registers_reg_12_0_inst : HS65_LH_DFPRQX9 port map( D => n1786, CP => clk, 
                           RN => n6546, Q => registers_12_0_port);
   registers_reg_11_31_inst : HS65_LH_DFPRQX9 port map( D => n1785, CP => clk, 
                           RN => n6550, Q => registers_11_31_port);
   registers_reg_11_30_inst : HS65_LH_DFPRQX9 port map( D => n1784, CP => clk, 
                           RN => n6550, Q => registers_11_30_port);
   registers_reg_11_29_inst : HS65_LH_DFPRQX9 port map( D => n1783, CP => clk, 
                           RN => n6550, Q => registers_11_29_port);
   registers_reg_11_28_inst : HS65_LH_DFPRQX9 port map( D => n1782, CP => clk, 
                           RN => n6550, Q => registers_11_28_port);
   registers_reg_11_27_inst : HS65_LH_DFPRQX9 port map( D => n1781, CP => clk, 
                           RN => n6549, Q => registers_11_27_port);
   registers_reg_11_26_inst : HS65_LH_DFPRQX9 port map( D => n1780, CP => clk, 
                           RN => n6549, Q => registers_11_26_port);
   registers_reg_11_25_inst : HS65_LH_DFPRQX9 port map( D => n1779, CP => clk, 
                           RN => n6549, Q => registers_11_25_port);
   registers_reg_11_24_inst : HS65_LH_DFPRQX9 port map( D => n1778, CP => clk, 
                           RN => n6549, Q => registers_11_24_port);
   registers_reg_11_23_inst : HS65_LH_DFPRQX9 port map( D => n1777, CP => clk, 
                           RN => n6545, Q => registers_11_23_port);
   registers_reg_11_22_inst : HS65_LH_DFPRQX9 port map( D => n1776, CP => clk, 
                           RN => n6545, Q => registers_11_22_port);
   registers_reg_11_21_inst : HS65_LH_DFPRQX9 port map( D => n1775, CP => clk, 
                           RN => n6545, Q => registers_11_21_port);
   registers_reg_11_20_inst : HS65_LH_DFPRQX9 port map( D => n1774, CP => clk, 
                           RN => n6545, Q => registers_11_20_port);
   registers_reg_11_19_inst : HS65_LH_DFPRQX9 port map( D => n1773, CP => clk, 
                           RN => n6552, Q => registers_11_19_port);
   registers_reg_11_18_inst : HS65_LH_DFPRQX9 port map( D => n1772, CP => clk, 
                           RN => n6548, Q => registers_11_18_port);
   registers_reg_11_17_inst : HS65_LH_DFPRQX9 port map( D => n1771, CP => clk, 
                           RN => n6548, Q => registers_11_17_port);
   registers_reg_11_16_inst : HS65_LH_DFPRQX9 port map( D => n1770, CP => clk, 
                           RN => n6548, Q => registers_11_16_port);
   registers_reg_11_15_inst : HS65_LH_DFPRQX9 port map( D => n1769, CP => clk, 
                           RN => n6541, Q => registers_11_15_port);
   registers_reg_11_14_inst : HS65_LH_DFPRQX9 port map( D => n1768, CP => clk, 
                           RN => n6541, Q => registers_11_14_port);
   registers_reg_11_13_inst : HS65_LH_DFPRQX9 port map( D => n1767, CP => clk, 
                           RN => n6541, Q => registers_11_13_port);
   registers_reg_11_12_inst : HS65_LH_DFPRQX9 port map( D => n1766, CP => clk, 
                           RN => n6541, Q => registers_11_12_port);
   registers_reg_11_11_inst : HS65_LH_DFPRQX9 port map( D => n1765, CP => clk, 
                           RN => n6541, Q => registers_11_11_port);
   registers_reg_11_10_inst : HS65_LH_DFPRQX9 port map( D => n1764, CP => clk, 
                           RN => n6541, Q => registers_11_10_port);
   registers_reg_11_9_inst : HS65_LH_DFPRQX9 port map( D => n1763, CP => clk, 
                           RN => n6541, Q => registers_11_9_port);
   registers_reg_11_8_inst : HS65_LH_DFPRQX9 port map( D => n1762, CP => clk, 
                           RN => n6550, Q => registers_11_8_port);
   registers_reg_11_7_inst : HS65_LH_DFPRQX9 port map( D => n1761, CP => clk, 
                           RN => n6551, Q => registers_11_7_port);
   registers_reg_11_6_inst : HS65_LH_DFPRQX9 port map( D => n1760, CP => clk, 
                           RN => n6551, Q => registers_11_6_port);
   registers_reg_11_5_inst : HS65_LH_DFPRQX9 port map( D => n1759, CP => clk, 
                           RN => n6551, Q => registers_11_5_port);
   registers_reg_11_4_inst : HS65_LH_DFPRQX9 port map( D => n1758, CP => clk, 
                           RN => n6551, Q => registers_11_4_port);
   registers_reg_11_3_inst : HS65_LH_DFPRQX9 port map( D => n1757, CP => clk, 
                           RN => n6551, Q => registers_11_3_port);
   registers_reg_11_2_inst : HS65_LH_DFPRQX9 port map( D => n1756, CP => clk, 
                           RN => n6551, Q => registers_11_2_port);
   registers_reg_11_1_inst : HS65_LH_DFPRQX9 port map( D => n1755, CP => clk, 
                           RN => n6551, Q => registers_11_1_port);
   registers_reg_11_0_inst : HS65_LH_DFPRQX9 port map( D => n1754, CP => clk, 
                           RN => n6551, Q => registers_11_0_port);
   registers_reg_10_31_inst : HS65_LH_DFPRQX9 port map( D => n1753, CP => clk, 
                           RN => n6551, Q => registers_10_31_port);
   registers_reg_10_30_inst : HS65_LH_DFPRQX9 port map( D => n1752, CP => clk, 
                           RN => n6551, Q => registers_10_30_port);
   registers_reg_10_29_inst : HS65_LH_DFPRQX9 port map( D => n1751, CP => clk, 
                           RN => n6551, Q => registers_10_29_port);
   registers_reg_10_28_inst : HS65_LH_DFPRQX9 port map( D => n1750, CP => clk, 
                           RN => n6563, Q => registers_10_28_port);
   registers_reg_10_27_inst : HS65_LH_DFPRQX9 port map( D => n1749, CP => clk, 
                           RN => n6563, Q => registers_10_27_port);
   registers_reg_10_26_inst : HS65_LH_DFPRQX9 port map( D => n1748, CP => clk, 
                           RN => n6563, Q => registers_10_26_port);
   registers_reg_10_25_inst : HS65_LH_DFPRQX9 port map( D => n1747, CP => clk, 
                           RN => n6563, Q => registers_10_25_port);
   registers_reg_10_24_inst : HS65_LH_DFPRQX9 port map( D => n1746, CP => clk, 
                           RN => n6549, Q => registers_10_24_port);
   registers_reg_10_23_inst : HS65_LH_DFPRQX9 port map( D => n1745, CP => clk, 
                           RN => n6549, Q => registers_10_23_port);
   registers_reg_10_22_inst : HS65_LH_DFPRQX9 port map( D => n1744, CP => clk, 
                           RN => n6549, Q => registers_10_22_port);
   registers_reg_10_21_inst : HS65_LH_DFPRQX9 port map( D => n1743, CP => clk, 
                           RN => n6549, Q => registers_10_21_port);
   registers_reg_10_20_inst : HS65_LH_DFPRQX9 port map( D => n1742, CP => clk, 
                           RN => n6549, Q => registers_10_20_port);
   registers_reg_10_19_inst : HS65_LH_DFPRQX9 port map( D => n1741, CP => clk, 
                           RN => n6549, Q => registers_10_19_port);
   registers_reg_10_18_inst : HS65_LH_DFPRQX9 port map( D => n1740, CP => clk, 
                           RN => n6549, Q => registers_10_18_port);
   registers_reg_10_17_inst : HS65_LH_DFPRQX9 port map( D => n1739, CP => clk, 
                           RN => n6549, Q => registers_10_17_port);
   registers_reg_10_16_inst : HS65_LH_DFPRQX9 port map( D => n1738, CP => clk, 
                           RN => n6564, Q => registers_10_16_port);
   registers_reg_10_15_inst : HS65_LH_DFPRQX9 port map( D => n1737, CP => clk, 
                           RN => n6564, Q => registers_10_15_port);
   registers_reg_10_14_inst : HS65_LH_DFPRQX9 port map( D => n1736, CP => clk, 
                           RN => n6564, Q => registers_10_14_port);
   registers_reg_10_13_inst : HS65_LH_DFPRQX9 port map( D => n1735, CP => clk, 
                           RN => n6564, Q => registers_10_13_port);
   registers_reg_10_12_inst : HS65_LH_DFPRQX9 port map( D => n1734, CP => clk, 
                           RN => n6559, Q => registers_10_12_port);
   registers_reg_10_11_inst : HS65_LH_DFPRQX9 port map( D => n1733, CP => clk, 
                           RN => n6559, Q => registers_10_11_port);
   registers_reg_10_10_inst : HS65_LH_DFPRQX9 port map( D => n1732, CP => clk, 
                           RN => n6559, Q => registers_10_10_port);
   registers_reg_10_9_inst : HS65_LH_DFPRQX9 port map( D => n1731, CP => clk, 
                           RN => n6559, Q => registers_10_9_port);
   registers_reg_10_8_inst : HS65_LH_DFPRQX9 port map( D => n1730, CP => clk, 
                           RN => n6559, Q => registers_10_8_port);
   registers_reg_10_7_inst : HS65_LH_DFPRQX9 port map( D => n1729, CP => clk, 
                           RN => n6559, Q => registers_10_7_port);
   registers_reg_10_6_inst : HS65_LH_DFPRQX9 port map( D => n1728, CP => clk, 
                           RN => n6559, Q => registers_10_6_port);
   registers_reg_10_5_inst : HS65_LH_DFPRQX9 port map( D => n1727, CP => clk, 
                           RN => n6559, Q => registers_10_5_port);
   registers_reg_10_4_inst : HS65_LH_DFPRQX9 port map( D => n1726, CP => clk, 
                           RN => n6540, Q => registers_10_4_port);
   registers_reg_10_3_inst : HS65_LH_DFPRQX9 port map( D => n1725, CP => clk, 
                           RN => n6540, Q => registers_10_3_port);
   registers_reg_10_2_inst : HS65_LH_DFPRQX9 port map( D => n1724, CP => clk, 
                           RN => n6540, Q => registers_10_2_port);
   registers_reg_10_1_inst : HS65_LH_DFPRQX9 port map( D => n1723, CP => clk, 
                           RN => n6540, Q => registers_10_1_port);
   registers_reg_10_0_inst : HS65_LH_DFPRQX9 port map( D => n1722, CP => clk, 
                           RN => n6540, Q => registers_10_0_port);
   registers_reg_7_31_inst : HS65_LH_DFPRQX9 port map( D => n1657, CP => clk, 
                           RN => n6545, Q => registers_7_31_port);
   registers_reg_7_30_inst : HS65_LH_DFPRQX9 port map( D => n1656, CP => clk, 
                           RN => n6545, Q => registers_7_30_port);
   registers_reg_7_29_inst : HS65_LH_DFPRQX9 port map( D => n1655, CP => clk, 
                           RN => n6545, Q => registers_7_29_port);
   registers_reg_7_28_inst : HS65_LH_DFPRQX9 port map( D => n1654, CP => clk, 
                           RN => n6545, Q => registers_7_28_port);
   registers_reg_7_27_inst : HS65_LH_DFPRQX9 port map( D => n1653, CP => clk, 
                           RN => n6546, Q => registers_7_27_port);
   registers_reg_7_26_inst : HS65_LH_DFPRQX9 port map( D => n1652, CP => clk, 
                           RN => n6546, Q => registers_7_26_port);
   registers_reg_7_25_inst : HS65_LH_DFPRQX9 port map( D => n1651, CP => clk, 
                           RN => n6546, Q => registers_7_25_port);
   registers_reg_7_24_inst : HS65_LH_DFPRQX9 port map( D => n1650, CP => clk, 
                           RN => n6546, Q => registers_7_24_port);
   registers_reg_7_23_inst : HS65_LH_DFPRQX9 port map( D => n1649, CP => clk, 
                           RN => n6537, Q => registers_7_23_port);
   registers_reg_7_22_inst : HS65_LH_DFPRQX9 port map( D => n1648, CP => clk, 
                           RN => n6565, Q => registers_7_22_port);
   registers_reg_7_21_inst : HS65_LH_DFPRQX9 port map( D => n1647, CP => clk, 
                           RN => n6565, Q => registers_7_21_port);
   registers_reg_7_20_inst : HS65_LH_DFPRQX9 port map( D => n1646, CP => clk, 
                           RN => n6565, Q => registers_7_20_port);
   registers_reg_7_19_inst : HS65_LH_DFPRQX9 port map( D => n1645, CP => clk, 
                           RN => n6565, Q => registers_7_19_port);
   registers_reg_7_18_inst : HS65_LH_DFPRQX9 port map( D => n1644, CP => clk, 
                           RN => n6562, Q => registers_7_18_port);
   registers_reg_7_17_inst : HS65_LH_DFPRQX9 port map( D => n1643, CP => clk, 
                           RN => n6562, Q => registers_7_17_port);
   registers_reg_7_16_inst : HS65_LH_DFPRQX9 port map( D => n1642, CP => clk, 
                           RN => n6562, Q => registers_7_16_port);
   registers_reg_7_15_inst : HS65_LH_DFPRQX9 port map( D => n1641, CP => clk, 
                           RN => n6558, Q => registers_7_15_port);
   registers_reg_7_14_inst : HS65_LH_DFPRQX9 port map( D => n1640, CP => clk, 
                           RN => n6558, Q => registers_7_14_port);
   registers_reg_7_13_inst : HS65_LH_DFPRQX9 port map( D => n1639, CP => clk, 
                           RN => n6558, Q => registers_7_13_port);
   registers_reg_7_12_inst : HS65_LH_DFPRQX9 port map( D => n1638, CP => clk, 
                           RN => n6558, Q => registers_7_12_port);
   registers_reg_7_11_inst : HS65_LH_DFPRQX9 port map( D => n1637, CP => clk, 
                           RN => n6564, Q => registers_7_11_port);
   registers_reg_7_10_inst : HS65_LH_DFPRQX9 port map( D => n1636, CP => clk, 
                           RN => n6564, Q => registers_7_10_port);
   registers_reg_7_9_inst : HS65_LH_DFPRQX9 port map( D => n1635, CP => clk, RN
                           => n6564, Q => registers_7_9_port);
   registers_reg_7_8_inst : HS65_LH_DFPRQX9 port map( D => n1634, CP => clk, RN
                           => n6564, Q => registers_7_8_port);
   registers_reg_7_7_inst : HS65_LH_DFPRQX9 port map( D => n1633, CP => clk, RN
                           => n6562, Q => registers_7_7_port);
   registers_reg_7_6_inst : HS65_LH_DFPRQX9 port map( D => n1632, CP => clk, RN
                           => n6562, Q => registers_7_6_port);
   registers_reg_7_5_inst : HS65_LH_DFPRQX9 port map( D => n1631, CP => clk, RN
                           => n6562, Q => registers_7_5_port);
   registers_reg_7_4_inst : HS65_LH_DFPRQX9 port map( D => n1630, CP => clk, RN
                           => n6562, Q => registers_7_4_port);
   registers_reg_7_3_inst : HS65_LH_DFPRQX9 port map( D => n1629, CP => clk, RN
                           => n6562, Q => registers_7_3_port);
   registers_reg_7_2_inst : HS65_LH_DFPRQX9 port map( D => n1628, CP => clk, RN
                           => n6562, Q => registers_7_2_port);
   registers_reg_7_1_inst : HS65_LH_DFPRQX9 port map( D => n1627, CP => clk, RN
                           => n6562, Q => registers_7_1_port);
   registers_reg_7_0_inst : HS65_LH_DFPRQX9 port map( D => n1626, CP => clk, RN
                           => n6562, Q => registers_7_0_port);
   registers_reg_6_31_inst : HS65_LH_DFPRQX9 port map( D => n1625, CP => clk, 
                           RN => n6567, Q => registers_6_31_port);
   registers_reg_6_30_inst : HS65_LH_DFPRQX9 port map( D => n1624, CP => clk, 
                           RN => n6567, Q => registers_6_30_port);
   registers_reg_6_29_inst : HS65_LH_DFPRQX9 port map( D => n1623, CP => clk, 
                           RN => n6567, Q => registers_6_29_port);
   registers_reg_6_28_inst : HS65_LH_DFPRQX9 port map( D => n1622, CP => clk, 
                           RN => n6567, Q => registers_6_28_port);
   registers_reg_6_27_inst : HS65_LH_DFPRQX9 port map( D => n1621, CP => clk, 
                           RN => n6568, Q => registers_6_27_port);
   registers_reg_6_26_inst : HS65_LH_DFPRQX9 port map( D => n1620, CP => clk, 
                           RN => n6568, Q => registers_6_26_port);
   registers_reg_6_25_inst : HS65_LH_DFPRQX9 port map( D => n1619, CP => clk, 
                           RN => n6568, Q => registers_6_25_port);
   registers_reg_6_24_inst : HS65_LH_DFPRQX9 port map( D => n1618, CP => clk, 
                           RN => n6566, Q => registers_6_24_port);
   registers_reg_6_23_inst : HS65_LH_DFPRQX9 port map( D => n1617, CP => clk, 
                           RN => n6566, Q => registers_6_23_port);
   registers_reg_6_22_inst : HS65_LH_DFPRQX9 port map( D => n1616, CP => clk, 
                           RN => n6566, Q => registers_6_22_port);
   registers_reg_6_21_inst : HS65_LH_DFPRQX9 port map( D => n1615, CP => clk, 
                           RN => n6566, Q => registers_6_21_port);
   registers_reg_6_20_inst : HS65_LH_DFPRQX9 port map( D => n1614, CP => clk, 
                           RN => n6566, Q => registers_6_20_port);
   registers_reg_6_19_inst : HS65_LH_DFPRQX9 port map( D => n1613, CP => clk, 
                           RN => n6598, Q => registers_6_19_port);
   registers_reg_6_18_inst : HS65_LH_DFPRQX9 port map( D => n1612, CP => clk, 
                           RN => n6597, Q => registers_6_18_port);
   registers_reg_6_17_inst : HS65_LH_DFPRQX9 port map( D => n1611, CP => clk, 
                           RN => n6597, Q => registers_6_17_port);
   registers_reg_6_16_inst : HS65_LH_DFPRQX9 port map( D => n1610, CP => clk, 
                           RN => n6597, Q => registers_6_16_port);
   registers_reg_6_15_inst : HS65_LH_DFPRQX9 port map( D => n1609, CP => clk, 
                           RN => n6596, Q => registers_6_15_port);
   registers_reg_6_14_inst : HS65_LH_DFPRQX9 port map( D => n1608, CP => clk, 
                           RN => n6596, Q => registers_6_14_port);
   registers_reg_6_13_inst : HS65_LH_DFPRQX9 port map( D => n1607, CP => clk, 
                           RN => n6596, Q => registers_6_13_port);
   registers_reg_6_12_inst : HS65_LH_DFPRQX9 port map( D => n1606, CP => clk, 
                           RN => n6596, Q => registers_6_12_port);
   registers_reg_6_11_inst : HS65_LH_DFPRQX9 port map( D => n1605, CP => clk, 
                           RN => n6596, Q => registers_6_11_port);
   registers_reg_6_10_inst : HS65_LH_DFPRQX9 port map( D => n1604, CP => clk, 
                           RN => n6596, Q => registers_6_10_port);
   registers_reg_6_9_inst : HS65_LH_DFPRQX9 port map( D => n1603, CP => clk, RN
                           => n6596, Q => registers_6_9_port);
   registers_reg_6_8_inst : HS65_LH_DFPRQX9 port map( D => n1602, CP => clk, RN
                           => n6596, Q => registers_6_8_port);
   registers_reg_6_7_inst : HS65_LH_DFPRQX9 port map( D => n1601, CP => clk, RN
                           => n6595, Q => registers_6_7_port);
   registers_reg_6_6_inst : HS65_LH_DFPRQX9 port map( D => n1600, CP => clk, RN
                           => n6595, Q => registers_6_6_port);
   registers_reg_6_5_inst : HS65_LH_DFPRQX9 port map( D => n1599, CP => clk, RN
                           => n6595, Q => registers_6_5_port);
   registers_reg_6_4_inst : HS65_LH_DFPRQX9 port map( D => n1598, CP => clk, RN
                           => n6595, Q => registers_6_4_port);
   registers_reg_6_3_inst : HS65_LH_DFPRQX9 port map( D => n1597, CP => clk, RN
                           => n6595, Q => registers_6_3_port);
   registers_reg_6_2_inst : HS65_LH_DFPRQX9 port map( D => n1596, CP => clk, RN
                           => n6595, Q => registers_6_2_port);
   registers_reg_6_1_inst : HS65_LH_DFPRQX9 port map( D => n1595, CP => clk, RN
                           => n6595, Q => registers_6_1_port);
   registers_reg_6_0_inst : HS65_LH_DFPRQX9 port map( D => n1594, CP => clk, RN
                           => n6595, Q => registers_6_0_port);
   registers_reg_5_31_inst : HS65_LH_DFPRQX9 port map( D => n1593, CP => clk, 
                           RN => n6537, Q => registers_5_31_port);
   registers_reg_5_30_inst : HS65_LH_DFPRQX9 port map( D => n1592, CP => clk, 
                           RN => n6537, Q => registers_5_30_port);
   registers_reg_5_29_inst : HS65_LH_DFPRQX9 port map( D => n1591, CP => clk, 
                           RN => n6537, Q => registers_5_29_port);
   registers_reg_5_28_inst : HS65_LH_DFPRQX9 port map( D => n1590, CP => clk, 
                           RN => n6544, Q => registers_5_28_port);
   registers_reg_5_27_inst : HS65_LH_DFPRQX9 port map( D => n1589, CP => clk, 
                           RN => n6544, Q => registers_5_27_port);
   registers_reg_5_26_inst : HS65_LH_DFPRQX9 port map( D => n1588, CP => clk, 
                           RN => n6544, Q => registers_5_26_port);
   registers_reg_5_25_inst : HS65_LH_DFPRQX9 port map( D => n1587, CP => clk, 
                           RN => n6544, Q => registers_5_25_port);
   registers_reg_5_24_inst : HS65_LH_DFPRQX9 port map( D => n1586, CP => clk, 
                           RN => n6538, Q => registers_5_24_port);
   registers_reg_5_23_inst : HS65_LH_DFPRQX9 port map( D => n1585, CP => clk, 
                           RN => n6538, Q => registers_5_23_port);
   registers_reg_5_22_inst : HS65_LH_DFPRQX9 port map( D => n1584, CP => clk, 
                           RN => n6538, Q => registers_5_22_port);
   registers_reg_5_21_inst : HS65_LH_DFPRQX9 port map( D => n1583, CP => clk, 
                           RN => n6538, Q => registers_5_21_port);
   registers_reg_5_20_inst : HS65_LH_DFPRQX9 port map( D => n1582, CP => clk, 
                           RN => n6598, Q => registers_5_20_port);
   registers_reg_5_19_inst : HS65_LH_DFPRQX9 port map( D => n1581, CP => clk, 
                           RN => n6598, Q => registers_5_19_port);
   registers_reg_5_18_inst : HS65_LH_DFPRQX9 port map( D => n1580, CP => clk, 
                           RN => n6597, Q => registers_5_18_port);
   registers_reg_5_17_inst : HS65_LH_DFPRQX9 port map( D => n1579, CP => clk, 
                           RN => n6597, Q => registers_5_17_port);
   registers_reg_5_16_inst : HS65_LH_DFPRQX9 port map( D => n1578, CP => clk, 
                           RN => n6543, Q => registers_5_16_port);
   registers_reg_5_15_inst : HS65_LH_DFPRQX9 port map( D => n1577, CP => clk, 
                           RN => n6543, Q => registers_5_15_port);
   registers_reg_5_14_inst : HS65_LH_DFPRQX9 port map( D => n1576, CP => clk, 
                           RN => n6543, Q => registers_5_14_port);
   registers_reg_5_13_inst : HS65_LH_DFPRQX9 port map( D => n1575, CP => clk, 
                           RN => n6543, Q => registers_5_13_port);
   registers_reg_5_12_inst : HS65_LH_DFPRQX9 port map( D => n1574, CP => clk, 
                           RN => n6537, Q => registers_5_12_port);
   registers_reg_5_11_inst : HS65_LH_DFPRQX9 port map( D => n1573, CP => clk, 
                           RN => n6537, Q => registers_5_11_port);
   registers_reg_5_10_inst : HS65_LH_DFPRQX9 port map( D => n1572, CP => clk, 
                           RN => n6537, Q => registers_5_10_port);
   registers_reg_5_9_inst : HS65_LH_DFPRQX9 port map( D => n1571, CP => clk, RN
                           => n6537, Q => registers_5_9_port);
   registers_reg_5_8_inst : HS65_LH_DFPRQX9 port map( D => n1570, CP => clk, RN
                           => n6537, Q => registers_5_8_port);
   registers_reg_5_7_inst : HS65_LH_DFPRQX9 port map( D => n1569, CP => clk, RN
                           => n6537, Q => registers_5_7_port);
   registers_reg_5_6_inst : HS65_LH_DFPRQX9 port map( D => n1568, CP => clk, RN
                           => n6537, Q => registers_5_6_port);
   registers_reg_5_5_inst : HS65_LH_DFPRQX9 port map( D => n1567, CP => clk, RN
                           => n6537, Q => registers_5_5_port);
   registers_reg_5_4_inst : HS65_LH_DFPRQX9 port map( D => n1566, CP => clk, RN
                           => n6543, Q => registers_5_4_port);
   registers_reg_5_3_inst : HS65_LH_DFPRQX9 port map( D => n1565, CP => clk, RN
                           => n6543, Q => registers_5_3_port);
   registers_reg_5_2_inst : HS65_LH_DFPRQX9 port map( D => n1564, CP => clk, RN
                           => n6543, Q => registers_5_2_port);
   registers_reg_5_1_inst : HS65_LH_DFPRQX9 port map( D => n1563, CP => clk, RN
                           => n6543, Q => registers_5_1_port);
   registers_reg_5_0_inst : HS65_LH_DFPRQX9 port map( D => n1562, CP => clk, RN
                           => n6543, Q => registers_5_0_port);
   registers_reg_4_31_inst : HS65_LH_DFPRQX9 port map( D => n1561, CP => clk, 
                           RN => n6547, Q => registers_4_31_port);
   registers_reg_4_30_inst : HS65_LH_DFPRQX9 port map( D => n1560, CP => clk, 
                           RN => n6547, Q => registers_4_30_port);
   registers_reg_4_29_inst : HS65_LH_DFPRQX9 port map( D => n1559, CP => clk, 
                           RN => n6547, Q => registers_4_29_port);
   registers_reg_4_28_inst : HS65_LH_DFPRQX9 port map( D => n1558, CP => clk, 
                           RN => n6598, Q => registers_4_28_port);
   registers_reg_4_27_inst : HS65_LH_DFPRQX9 port map( D => n1557, CP => clk, 
                           RN => n6547, Q => registers_4_27_port);
   registers_reg_4_26_inst : HS65_LH_DFPRQX9 port map( D => n1556, CP => clk, 
                           RN => n6543, Q => registers_4_26_port);
   registers_reg_4_25_inst : HS65_LH_DFPRQX9 port map( D => n1555, CP => clk, 
                           RN => n6543, Q => registers_4_25_port);
   registers_reg_4_24_inst : HS65_LH_DFPRQX9 port map( D => n1554, CP => clk, 
                           RN => n6548, Q => registers_4_24_port);
   registers_reg_4_23_inst : HS65_LH_DFPRQX9 port map( D => n1553, CP => clk, 
                           RN => n6548, Q => registers_4_23_port);
   registers_reg_4_22_inst : HS65_LH_DFPRQX9 port map( D => n1552, CP => clk, 
                           RN => n6548, Q => registers_4_22_port);
   registers_reg_4_21_inst : HS65_LH_DFPRQX9 port map( D => n1551, CP => clk, 
                           RN => n6548, Q => registers_4_21_port);
   registers_reg_4_20_inst : HS65_LH_DFPRQX9 port map( D => n1550, CP => clk, 
                           RN => n6547, Q => registers_4_20_port);
   registers_reg_4_19_inst : HS65_LH_DFPRQX9 port map( D => n1549, CP => clk, 
                           RN => n6547, Q => registers_4_19_port);
   registers_reg_4_18_inst : HS65_LH_DFPRQX9 port map( D => n1548, CP => clk, 
                           RN => n6547, Q => registers_4_18_port);
   registers_reg_4_17_inst : HS65_LH_DFPRQX9 port map( D => n1547, CP => clk, 
                           RN => n6547, Q => registers_4_17_port);
   registers_reg_4_16_inst : HS65_LH_DFPRQX9 port map( D => n1546, CP => clk, 
                           RN => n6547, Q => registers_4_16_port);
   registers_reg_4_15_inst : HS65_LH_DFPRQX9 port map( D => n1545, CP => clk, 
                           RN => n6547, Q => registers_4_15_port);
   registers_reg_4_14_inst : HS65_LH_DFPRQX9 port map( D => n1544, CP => clk, 
                           RN => n6547, Q => registers_4_14_port);
   registers_reg_4_13_inst : HS65_LH_DFPRQX9 port map( D => n1543, CP => clk, 
                           RN => n6547, Q => registers_4_13_port);
   registers_reg_4_12_inst : HS65_LH_DFPRQX9 port map( D => n1542, CP => clk, 
                           RN => n6566, Q => registers_4_12_port);
   registers_reg_4_11_inst : HS65_LH_DFPRQX9 port map( D => n1541, CP => clk, 
                           RN => n6548, Q => registers_4_11_port);
   registers_reg_4_10_inst : HS65_LH_DFPRQX9 port map( D => n1540, CP => clk, 
                           RN => n6548, Q => registers_4_10_port);
   registers_reg_4_9_inst : HS65_LH_DFPRQX9 port map( D => n1539, CP => clk, RN
                           => n6548, Q => registers_4_9_port);
   registers_reg_4_8_inst : HS65_LH_DFPRQX9 port map( D => n1538, CP => clk, RN
                           => n6563, Q => registers_4_8_port);
   registers_reg_4_7_inst : HS65_LH_DFPRQX9 port map( D => n1537, CP => clk, RN
                           => n6563, Q => registers_4_7_port);
   registers_reg_4_6_inst : HS65_LH_DFPRQX9 port map( D => n1536, CP => clk, RN
                           => n6563, Q => registers_4_6_port);
   registers_reg_4_5_inst : HS65_LH_DFPRQX9 port map( D => n1535, CP => clk, RN
                           => n6563, Q => registers_4_5_port);
   registers_reg_4_4_inst : HS65_LH_DFPRQX9 port map( D => n1534, CP => clk, RN
                           => n6563, Q => registers_4_4_port);
   registers_reg_4_3_inst : HS65_LH_DFPRQX9 port map( D => n1533, CP => clk, RN
                           => n6563, Q => registers_4_3_port);
   registers_reg_4_2_inst : HS65_LH_DFPRQX9 port map( D => n1532, CP => clk, RN
                           => n6563, Q => registers_4_2_port);
   registers_reg_4_1_inst : HS65_LH_DFPRQX9 port map( D => n1531, CP => clk, RN
                           => n6563, Q => registers_4_1_port);
   registers_reg_4_0_inst : HS65_LH_DFPRQX9 port map( D => n1530, CP => clk, RN
                           => n6548, Q => registers_4_0_port);
   registers_reg_3_31_inst : HS65_LH_DFPRQX9 port map( D => n1529, CP => clk, 
                           RN => n6554, Q => registers_3_31_port);
   registers_reg_3_30_inst : HS65_LH_DFPRQX9 port map( D => n1528, CP => clk, 
                           RN => n6554, Q => registers_3_30_port);
   registers_reg_3_29_inst : HS65_LH_DFPRQX9 port map( D => n1527, CP => clk, 
                           RN => n6554, Q => registers_3_29_port);
   registers_reg_3_28_inst : HS65_LH_DFPRQX9 port map( D => n1526, CP => clk, 
                           RN => n6554, Q => registers_3_28_port);
   registers_reg_3_27_inst : HS65_LH_DFPRQX9 port map( D => n1525, CP => clk, 
                           RN => n6553, Q => registers_3_27_port);
   registers_reg_3_26_inst : HS65_LH_DFPRQX9 port map( D => n1524, CP => clk, 
                           RN => n6553, Q => registers_3_26_port);
   registers_reg_3_25_inst : HS65_LH_DFPRQX9 port map( D => n1523, CP => clk, 
                           RN => n6551, Q => registers_3_25_port);
   registers_reg_3_24_inst : HS65_LH_DFPRQX9 port map( D => n1522, CP => clk, 
                           RN => n6550, Q => registers_3_24_port);
   registers_reg_3_23_inst : HS65_LH_DFPRQX9 port map( D => n1521, CP => clk, 
                           RN => n6552, Q => registers_3_23_port);
   registers_reg_3_22_inst : HS65_LH_DFPRQX9 port map( D => n1520, CP => clk, 
                           RN => n6552, Q => registers_3_22_port);
   registers_reg_3_21_inst : HS65_LH_DFPRQX9 port map( D => n1519, CP => clk, 
                           RN => n6552, Q => registers_3_21_port);
   registers_reg_3_20_inst : HS65_LH_DFPRQX9 port map( D => n1518, CP => clk, 
                           RN => n6576, Q => registers_3_20_port);
   registers_reg_3_19_inst : HS65_LH_DFPRQX9 port map( D => n1517, CP => clk, 
                           RN => n6576, Q => registers_3_19_port);
   registers_reg_3_18_inst : HS65_LH_DFPRQX9 port map( D => n1516, CP => clk, 
                           RN => n6576, Q => registers_3_18_port);
   registers_reg_3_17_inst : HS65_LH_DFPRQX9 port map( D => n1515, CP => clk, 
                           RN => n6567, Q => registers_3_17_port);
   registers_reg_3_16_inst : HS65_LH_DFPRQX9 port map( D => n1514, CP => clk, 
                           RN => n6578, Q => registers_3_16_port);
   registers_reg_3_15_inst : HS65_LH_DFPRQX9 port map( D => n1513, CP => clk, 
                           RN => n6575, Q => registers_3_15_port);
   registers_reg_3_14_inst : HS65_LH_DFPRQX9 port map( D => n1512, CP => clk, 
                           RN => n6575, Q => registers_3_14_port);
   registers_reg_3_13_inst : HS65_LH_DFPRQX9 port map( D => n1511, CP => clk, 
                           RN => n6575, Q => registers_3_13_port);
   registers_reg_3_12_inst : HS65_LH_DFPRQX9 port map( D => n1510, CP => clk, 
                           RN => n6575, Q => registers_3_12_port);
   registers_reg_3_11_inst : HS65_LH_DFPRQX9 port map( D => n1509, CP => clk, 
                           RN => n6575, Q => registers_3_11_port);
   registers_reg_3_10_inst : HS65_LH_DFPRQX9 port map( D => n1508, CP => clk, 
                           RN => n6575, Q => registers_3_10_port);
   registers_reg_3_9_inst : HS65_LH_DFPRQX9 port map( D => n1507, CP => clk, RN
                           => n6575, Q => registers_3_9_port);
   registers_reg_3_8_inst : HS65_LH_DFPRQX9 port map( D => n1506, CP => clk, RN
                           => n6567, Q => registers_3_8_port);
   registers_reg_3_7_inst : HS65_LH_DFPRQX9 port map( D => n1505, CP => clk, RN
                           => n6565, Q => registers_3_7_port);
   registers_reg_3_6_inst : HS65_LH_DFPRQX9 port map( D => n1504, CP => clk, RN
                           => n6565, Q => registers_3_6_port);
   registers_reg_3_5_inst : HS65_LH_DFPRQX9 port map( D => n1503, CP => clk, RN
                           => n6565, Q => registers_3_5_port);
   registers_reg_3_4_inst : HS65_LH_DFPRQX9 port map( D => n1502, CP => clk, RN
                           => n6565, Q => registers_3_4_port);
   registers_reg_3_3_inst : HS65_LH_DFPRQX9 port map( D => n1501, CP => clk, RN
                           => n6565, Q => registers_3_3_port);
   registers_reg_3_2_inst : HS65_LH_DFPRQX9 port map( D => n1500, CP => clk, RN
                           => n6565, Q => registers_3_2_port);
   registers_reg_3_1_inst : HS65_LH_DFPRQX9 port map( D => n1499, CP => clk, RN
                           => n6565, Q => registers_3_1_port);
   registers_reg_3_0_inst : HS65_LH_DFPRQX9 port map( D => n1498, CP => clk, RN
                           => n6565, Q => registers_3_0_port);
   registers_reg_2_31_inst : HS65_LH_DFPRQX9 port map( D => n1497, CP => clk, 
                           RN => n6575, Q => registers_2_31_port);
   registers_reg_2_30_inst : HS65_LH_DFPRQX9 port map( D => n1496, CP => clk, 
                           RN => n6575, Q => registers_2_30_port);
   registers_reg_2_29_inst : HS65_LH_DFPRQX9 port map( D => n1495, CP => clk, 
                           RN => n6575, Q => registers_2_29_port);
   registers_reg_2_28_inst : HS65_LH_DFPRQX9 port map( D => n1494, CP => clk, 
                           RN => n6580, Q => registers_2_28_port);
   registers_reg_2_27_inst : HS65_LH_DFPRQX9 port map( D => n1493, CP => clk, 
                           RN => n6580, Q => registers_2_27_port);
   registers_reg_2_26_inst : HS65_LH_DFPRQX9 port map( D => n1492, CP => clk, 
                           RN => n6580, Q => registers_2_26_port);
   registers_reg_2_25_inst : HS65_LH_DFPRQX9 port map( D => n1491, CP => clk, 
                           RN => n6580, Q => registers_2_25_port);
   registers_reg_2_24_inst : HS65_LH_DFPRQX9 port map( D => n1490, CP => clk, 
                           RN => n6568, Q => registers_2_24_port);
   registers_reg_2_23_inst : HS65_LH_DFPRQX9 port map( D => n1489, CP => clk, 
                           RN => n6566, Q => registers_2_23_port);
   registers_reg_2_22_inst : HS65_LH_DFPRQX9 port map( D => n1488, CP => clk, 
                           RN => n6566, Q => registers_2_22_port);
   registers_reg_2_21_inst : HS65_LH_DFPRQX9 port map( D => n1487, CP => clk, 
                           RN => n6566, Q => registers_2_21_port);
   registers_reg_2_20_inst : HS65_LH_DFPRQX9 port map( D => n1486, CP => clk, 
                           RN => n6566, Q => registers_2_20_port);
   registers_reg_2_19_inst : HS65_LH_DFPRQX9 port map( D => n1485, CP => clk, 
                           RN => n6566, Q => registers_2_19_port);
   registers_reg_2_18_inst : HS65_LH_DFPRQX9 port map( D => n1484, CP => clk, 
                           RN => n6566, Q => registers_2_18_port);
   registers_reg_2_17_inst : HS65_LH_DFPRQX9 port map( D => n1483, CP => clk, 
                           RN => n6579, Q => registers_2_17_port);
   registers_reg_2_16_inst : HS65_LH_DFPRQX9 port map( D => n1482, CP => clk, 
                           RN => n6579, Q => registers_2_16_port);
   registers_reg_2_15_inst : HS65_LH_DFPRQX9 port map( D => n1481, CP => clk, 
                           RN => n6578, Q => registers_2_15_port);
   registers_reg_2_14_inst : HS65_LH_DFPRQX9 port map( D => n1480, CP => clk, 
                           RN => n6575, Q => registers_2_14_port);
   registers_reg_2_13_inst : HS65_LH_DFPRQX9 port map( D => n1479, CP => clk, 
                           RN => n6579, Q => registers_2_13_port);
   registers_reg_2_12_inst : HS65_LH_DFPRQX9 port map( D => n1478, CP => clk, 
                           RN => n6579, Q => registers_2_12_port);
   registers_reg_2_11_inst : HS65_LH_DFPRQX9 port map( D => n1477, CP => clk, 
                           RN => n6579, Q => registers_2_11_port);
   registers_reg_2_10_inst : HS65_LH_DFPRQX9 port map( D => n1476, CP => clk, 
                           RN => n6579, Q => registers_2_10_port);
   registers_reg_2_9_inst : HS65_LH_DFPRQX9 port map( D => n1475, CP => clk, RN
                           => n6579, Q => registers_2_9_port);
   registers_reg_2_8_inst : HS65_LH_DFPRQX9 port map( D => n1474, CP => clk, RN
                           => n6579, Q => registers_2_8_port);
   registers_reg_2_7_inst : HS65_LH_DFPRQX9 port map( D => n1473, CP => clk, RN
                           => n6579, Q => registers_2_7_port);
   registers_reg_2_6_inst : HS65_LH_DFPRQX9 port map( D => n1472, CP => clk, RN
                           => n6579, Q => registers_2_6_port);
   registers_reg_2_5_inst : HS65_LH_DFPRQX9 port map( D => n1471, CP => clk, RN
                           => n6567, Q => registers_2_5_port);
   registers_reg_2_4_inst : HS65_LH_DFPRQX9 port map( D => n1470, CP => clk, RN
                           => n6567, Q => registers_2_4_port);
   registers_reg_2_3_inst : HS65_LH_DFPRQX9 port map( D => n1469, CP => clk, RN
                           => n6567, Q => registers_2_3_port);
   registers_reg_2_2_inst : HS65_LH_DFPRQX9 port map( D => n1468, CP => clk, RN
                           => n6567, Q => registers_2_2_port);
   registers_reg_2_1_inst : HS65_LH_DFPRQX9 port map( D => n1467, CP => clk, RN
                           => n6567, Q => registers_2_1_port);
   registers_reg_2_0_inst : HS65_LH_DFPRQX9 port map( D => n1466, CP => clk, RN
                           => n6567, Q => registers_2_0_port);
   registers_reg_1_31_inst : HS65_LH_DFPRQX9 port map( D => n1465, CP => clk, 
                           RN => n6582, Q => registers_1_31_port);
   registers_reg_1_30_inst : HS65_LH_DFPRQX9 port map( D => n1464, CP => clk, 
                           RN => n6582, Q => registers_1_30_port);
   registers_reg_1_29_inst : HS65_LH_DFPRQX9 port map( D => n1463, CP => clk, 
                           RN => n6582, Q => registers_1_29_port);
   registers_reg_1_28_inst : HS65_LH_DFPRQX9 port map( D => n1462, CP => clk, 
                           RN => n6582, Q => registers_1_28_port);
   registers_reg_1_27_inst : HS65_LH_DFPRQX9 port map( D => n1461, CP => clk, 
                           RN => n6575, Q => registers_1_27_port);
   registers_reg_1_26_inst : HS65_LH_DFPRQX9 port map( D => n1460, CP => clk, 
                           RN => n6576, Q => registers_1_26_port);
   registers_reg_1_25_inst : HS65_LH_DFPRQX9 port map( D => n1459, CP => clk, 
                           RN => n6581, Q => registers_1_25_port);
   registers_reg_1_24_inst : HS65_LH_DFPRQX9 port map( D => n1458, CP => clk, 
                           RN => n6581, Q => registers_1_24_port);
   registers_reg_1_23_inst : HS65_LH_DFPRQX9 port map( D => n1457, CP => clk, 
                           RN => n6581, Q => registers_1_23_port);
   registers_reg_1_22_inst : HS65_LH_DFPRQX9 port map( D => n1456, CP => clk, 
                           RN => n6581, Q => registers_1_22_port);
   registers_reg_1_21_inst : HS65_LH_DFPRQX9 port map( D => n1455, CP => clk, 
                           RN => n6581, Q => registers_1_21_port);
   registers_reg_1_20_inst : HS65_LH_DFPRQX9 port map( D => n1454, CP => clk, 
                           RN => n6581, Q => registers_1_20_port);
   registers_reg_1_19_inst : HS65_LH_DFPRQX9 port map( D => n1453, CP => clk, 
                           RN => n6581, Q => registers_1_19_port);
   registers_reg_1_18_inst : HS65_LH_DFPRQX9 port map( D => n1452, CP => clk, 
                           RN => n6581, Q => registers_1_18_port);
   registers_reg_1_17_inst : HS65_LH_DFPRQX9 port map( D => n1451, CP => clk, 
                           RN => n6581, Q => registers_1_17_port);
   registers_reg_1_16_inst : HS65_LH_DFPRQX9 port map( D => n1450, CP => clk, 
                           RN => n6581, Q => registers_1_16_port);
   registers_reg_1_15_inst : HS65_LH_DFPRQX9 port map( D => n1449, CP => clk, 
                           RN => n6581, Q => registers_1_15_port);
   registers_reg_1_14_inst : HS65_LH_DFPRQX9 port map( D => n1448, CP => clk, 
                           RN => n6581, Q => registers_1_14_port);
   registers_reg_1_13_inst : HS65_LH_DFPRQX9 port map( D => n1447, CP => clk, 
                           RN => n6564, Q => registers_1_13_port);
   registers_reg_1_12_inst : HS65_LH_DFPRQX9 port map( D => n1446, CP => clk, 
                           RN => n6564, Q => registers_1_12_port);
   registers_reg_1_11_inst : HS65_LH_DFPRQX9 port map( D => n1445, CP => clk, 
                           RN => n6564, Q => registers_1_11_port);
   registers_reg_1_10_inst : HS65_LH_DFPRQX9 port map( D => n1444, CP => clk, 
                           RN => n6564, Q => registers_1_10_port);
   registers_reg_1_9_inst : HS65_LH_DFPRQX9 port map( D => n1443, CP => clk, RN
                           => n6560, Q => registers_1_9_port);
   registers_reg_1_8_inst : HS65_LH_DFPRQX9 port map( D => n1442, CP => clk, RN
                           => n6560, Q => registers_1_8_port);
   registers_reg_1_7_inst : HS65_LH_DFPRQX9 port map( D => n1441, CP => clk, RN
                           => n6560, Q => registers_1_7_port);
   registers_reg_1_6_inst : HS65_LH_DFPRQX9 port map( D => n1440, CP => clk, RN
                           => n6560, Q => registers_1_6_port);
   registers_reg_1_5_inst : HS65_LH_DFPRQX9 port map( D => n1439, CP => clk, RN
                           => n6560, Q => registers_1_5_port);
   registers_reg_1_4_inst : HS65_LH_DFPRQX9 port map( D => n1438, CP => clk, RN
                           => n6560, Q => registers_1_4_port);
   registers_reg_1_3_inst : HS65_LH_DFPRQX9 port map( D => n1437, CP => clk, RN
                           => n6560, Q => registers_1_3_port);
   registers_reg_1_2_inst : HS65_LH_DFPRQX9 port map( D => n1436, CP => clk, RN
                           => n6560, Q => registers_1_2_port);
   registers_reg_1_1_inst : HS65_LH_DFPRQX9 port map( D => n1435, CP => clk, RN
                           => n6558, Q => registers_1_1_port);
   registers_reg_1_0_inst : HS65_LH_DFPRQX9 port map( D => n1434, CP => clk, RN
                           => n6543, Q => registers_1_0_port);
   registers_reg_27_31_inst : HS65_LH_DFPRQNX9 port map( D => n2297, CP => clk,
                           RN => n6616, QN => n65);
   registers_reg_27_30_inst : HS65_LH_DFPRQNX9 port map( D => n2296, CP => clk,
                           RN => n6616, QN => n66);
   registers_reg_27_29_inst : HS65_LH_DFPRQNX9 port map( D => n2295, CP => clk,
                           RN => n6616, QN => n67);
   registers_reg_27_28_inst : HS65_LH_DFPRQNX9 port map( D => n2294, CP => clk,
                           RN => n6616, QN => n68);
   registers_reg_27_27_inst : HS65_LH_DFPRQNX9 port map( D => n2293, CP => clk,
                           RN => n6616, QN => n69);
   registers_reg_27_26_inst : HS65_LH_DFPRQNX9 port map( D => n2292, CP => clk,
                           RN => n6616, QN => n70);
   registers_reg_27_25_inst : HS65_LH_DFPRQNX9 port map( D => n2291, CP => clk,
                           RN => n6616, QN => n71);
   registers_reg_27_24_inst : HS65_LH_DFPRQNX9 port map( D => n2290, CP => clk,
                           RN => n6616, QN => n72);
   registers_reg_27_23_inst : HS65_LH_DFPRQNX9 port map( D => n2289, CP => clk,
                           RN => n6615, QN => n73);
   registers_reg_27_22_inst : HS65_LH_DFPRQNX9 port map( D => n2288, CP => clk,
                           RN => n6615, QN => n74);
   registers_reg_27_21_inst : HS65_LH_DFPRQNX9 port map( D => n2287, CP => clk,
                           RN => n6615, QN => n75);
   registers_reg_27_20_inst : HS65_LH_DFPRQNX9 port map( D => n2286, CP => clk,
                           RN => n6615, QN => n76);
   registers_reg_27_19_inst : HS65_LH_DFPRQNX9 port map( D => n2285, CP => clk,
                           RN => n6615, QN => n77);
   registers_reg_27_18_inst : HS65_LH_DFPRQNX9 port map( D => n2284, CP => clk,
                           RN => n6615, QN => n78);
   registers_reg_27_17_inst : HS65_LH_DFPRQNX9 port map( D => n2283, CP => clk,
                           RN => n6615, QN => n79);
   registers_reg_27_16_inst : HS65_LH_DFPRQNX9 port map( D => n2282, CP => clk,
                           RN => n6615, QN => n80);
   registers_reg_27_15_inst : HS65_LH_DFPRQNX9 port map( D => n2281, CP => clk,
                           RN => n6615, QN => n81);
   registers_reg_27_14_inst : HS65_LH_DFPRQNX9 port map( D => n2280, CP => clk,
                           RN => n6615, QN => n82);
   registers_reg_27_13_inst : HS65_LH_DFPRQNX9 port map( D => n2279, CP => clk,
                           RN => n6615, QN => n83);
   registers_reg_27_12_inst : HS65_LH_DFPRQNX9 port map( D => n2278, CP => clk,
                           RN => n6615, QN => n84);
   registers_reg_27_11_inst : HS65_LH_DFPRQNX9 port map( D => n2277, CP => clk,
                           RN => n6615, QN => n85);
   registers_reg_27_10_inst : HS65_LH_DFPRQNX9 port map( D => n2276, CP => clk,
                           RN => n6615, QN => n86);
   registers_reg_27_9_inst : HS65_LH_DFPRQNX9 port map( D => n2275, CP => clk, 
                           RN => n6614, QN => n87);
   registers_reg_27_8_inst : HS65_LH_DFPRQNX9 port map( D => n2274, CP => clk, 
                           RN => n6614, QN => n88);
   registers_reg_27_7_inst : HS65_LH_DFPRQNX9 port map( D => n2273, CP => clk, 
                           RN => n6614, QN => n89);
   registers_reg_27_6_inst : HS65_LH_DFPRQNX9 port map( D => n2272, CP => clk, 
                           RN => n6614, QN => n90);
   registers_reg_27_5_inst : HS65_LH_DFPRQNX9 port map( D => n2271, CP => clk, 
                           RN => n6614, QN => n91);
   registers_reg_27_4_inst : HS65_LH_DFPRQNX9 port map( D => n2270, CP => clk, 
                           RN => n6614, QN => n92);
   registers_reg_27_3_inst : HS65_LH_DFPRQNX9 port map( D => n2269, CP => clk, 
                           RN => n6614, QN => n93);
   registers_reg_27_2_inst : HS65_LH_DFPRQNX9 port map( D => n2268, CP => clk, 
                           RN => n6614, QN => n94);
   registers_reg_27_1_inst : HS65_LH_DFPRQNX9 port map( D => n2267, CP => clk, 
                           RN => n6614, QN => n95);
   registers_reg_27_0_inst : HS65_LH_DFPRQNX9 port map( D => n2266, CP => clk, 
                           RN => n6614, QN => n96);
   registers_reg_28_31_inst : HS65_LH_DFPRQNX9 port map( D => n2329, CP => clk,
                           RN => n6611, QN => n33);
   registers_reg_28_30_inst : HS65_LH_DFPRQNX9 port map( D => n2328, CP => clk,
                           RN => n6611, QN => n34);
   registers_reg_28_29_inst : HS65_LH_DFPRQNX9 port map( D => n2327, CP => clk,
                           RN => n6611, QN => n35);
   registers_reg_28_28_inst : HS65_LH_DFPRQNX9 port map( D => n2326, CP => clk,
                           RN => n6611, QN => n36);
   registers_reg_28_27_inst : HS65_LH_DFPRQNX9 port map( D => n2325, CP => clk,
                           RN => n6611, QN => n37);
   registers_reg_28_26_inst : HS65_LH_DFPRQNX9 port map( D => n2324, CP => clk,
                           RN => n6611, QN => n38);
   registers_reg_28_25_inst : HS65_LH_DFPRQNX9 port map( D => n2323, CP => clk,
                           RN => n6611, QN => n39);
   registers_reg_28_24_inst : HS65_LH_DFPRQNX9 port map( D => n2322, CP => clk,
                           RN => n6611, QN => n40);
   registers_reg_28_23_inst : HS65_LH_DFPRQNX9 port map( D => n2321, CP => clk,
                           RN => n6611, QN => n41);
   registers_reg_28_22_inst : HS65_LH_DFPRQNX9 port map( D => n2320, CP => clk,
                           RN => n6611, QN => n42);
   registers_reg_28_21_inst : HS65_LH_DFPRQNX9 port map( D => n2319, CP => clk,
                           RN => n6611, QN => n43);
   registers_reg_28_20_inst : HS65_LH_DFPRQNX9 port map( D => n2318, CP => clk,
                           RN => n6611, QN => n44);
   registers_reg_28_19_inst : HS65_LH_DFPRQNX9 port map( D => n2317, CP => clk,
                           RN => n6611, QN => n45);
   registers_reg_28_18_inst : HS65_LH_DFPRQNX9 port map( D => n2316, CP => clk,
                           RN => n6611, QN => n46);
   registers_reg_28_17_inst : HS65_LH_DFPRQNX9 port map( D => n2315, CP => clk,
                           RN => n6610, QN => n47);
   registers_reg_28_16_inst : HS65_LH_DFPRQNX9 port map( D => n2314, CP => clk,
                           RN => n6610, QN => n48);
   registers_reg_28_15_inst : HS65_LH_DFPRQNX9 port map( D => n2313, CP => clk,
                           RN => n6610, QN => n49);
   registers_reg_28_14_inst : HS65_LH_DFPRQNX9 port map( D => n2312, CP => clk,
                           RN => n6610, QN => n50);
   registers_reg_28_13_inst : HS65_LH_DFPRQNX9 port map( D => n2311, CP => clk,
                           RN => n6610, QN => n51);
   registers_reg_28_12_inst : HS65_LH_DFPRQNX9 port map( D => n2310, CP => clk,
                           RN => n6610, QN => n52);
   registers_reg_28_11_inst : HS65_LH_DFPRQNX9 port map( D => n2309, CP => clk,
                           RN => n6610, QN => n53);
   registers_reg_28_10_inst : HS65_LH_DFPRQNX9 port map( D => n2308, CP => clk,
                           RN => n6610, QN => n54);
   registers_reg_28_9_inst : HS65_LH_DFPRQNX9 port map( D => n2307, CP => clk, 
                           RN => n6610, QN => n55);
   registers_reg_28_8_inst : HS65_LH_DFPRQNX9 port map( D => n2306, CP => clk, 
                           RN => n6610, QN => n56);
   registers_reg_28_7_inst : HS65_LH_DFPRQNX9 port map( D => n2305, CP => clk, 
                           RN => n6610, QN => n57);
   registers_reg_28_6_inst : HS65_LH_DFPRQNX9 port map( D => n2304, CP => clk, 
                           RN => n6610, QN => n58);
   registers_reg_28_5_inst : HS65_LH_DFPRQNX9 port map( D => n2303, CP => clk, 
                           RN => n6610, QN => n59);
   registers_reg_28_4_inst : HS65_LH_DFPRQNX9 port map( D => n2302, CP => clk, 
                           RN => n6610, QN => n60);
   registers_reg_28_3_inst : HS65_LH_DFPRQNX9 port map( D => n2301, CP => clk, 
                           RN => n6609, QN => n61);
   registers_reg_28_2_inst : HS65_LH_DFPRQNX9 port map( D => n2300, CP => clk, 
                           RN => n6609, QN => n62);
   registers_reg_28_1_inst : HS65_LH_DFPRQNX9 port map( D => n2299, CP => clk, 
                           RN => n6609, QN => n63);
   registers_reg_28_0_inst : HS65_LH_DFPRQNX9 port map( D => n2298, CP => clk, 
                           RN => n6609, QN => n64);
   registers_reg_14_31_inst : HS65_LH_DFPRQNX9 port map( D => n1881, CP => clk,
                           RN => n6609, QN => n161);
   registers_reg_14_30_inst : HS65_LH_DFPRQNX9 port map( D => n1880, CP => clk,
                           RN => n6609, QN => n162);
   registers_reg_14_29_inst : HS65_LH_DFPRQNX9 port map( D => n1879, CP => clk,
                           RN => n6609, QN => n163);
   registers_reg_14_28_inst : HS65_LH_DFPRQNX9 port map( D => n1878, CP => clk,
                           RN => n6609, QN => n164);
   registers_reg_14_27_inst : HS65_LH_DFPRQNX9 port map( D => n1877, CP => clk,
                           RN => n6609, QN => n165);
   registers_reg_14_26_inst : HS65_LH_DFPRQNX9 port map( D => n1876, CP => clk,
                           RN => n6609, QN => n166);
   registers_reg_14_25_inst : HS65_LH_DFPRQNX9 port map( D => n1875, CP => clk,
                           RN => n6609, QN => n167);
   registers_reg_14_24_inst : HS65_LH_DFPRQNX9 port map( D => n1874, CP => clk,
                           RN => n6609, QN => n168);
   registers_reg_14_23_inst : HS65_LH_DFPRQNX9 port map( D => n1873, CP => clk,
                           RN => n6609, QN => n169);
   registers_reg_14_22_inst : HS65_LH_DFPRQNX9 port map( D => n1872, CP => clk,
                           RN => n6609, QN => n170);
   registers_reg_14_21_inst : HS65_LH_DFPRQNX9 port map( D => n1871, CP => clk,
                           RN => n6608, QN => n171);
   registers_reg_14_20_inst : HS65_LH_DFPRQNX9 port map( D => n1870, CP => clk,
                           RN => n6608, QN => n172);
   registers_reg_14_19_inst : HS65_LH_DFPRQNX9 port map( D => n1869, CP => clk,
                           RN => n6608, QN => n173);
   registers_reg_14_18_inst : HS65_LH_DFPRQNX9 port map( D => n1868, CP => clk,
                           RN => n6608, QN => n174);
   registers_reg_14_17_inst : HS65_LH_DFPRQNX9 port map( D => n1867, CP => clk,
                           RN => n6608, QN => n175);
   registers_reg_14_16_inst : HS65_LH_DFPRQNX9 port map( D => n1866, CP => clk,
                           RN => n6608, QN => n176);
   registers_reg_14_15_inst : HS65_LH_DFPRQNX9 port map( D => n1865, CP => clk,
                           RN => n6608, QN => n177);
   registers_reg_14_14_inst : HS65_LH_DFPRQNX9 port map( D => n1864, CP => clk,
                           RN => n6608, QN => n178);
   registers_reg_14_13_inst : HS65_LH_DFPRQNX9 port map( D => n1863, CP => clk,
                           RN => n6608, QN => n179);
   registers_reg_14_12_inst : HS65_LH_DFPRQNX9 port map( D => n1862, CP => clk,
                           RN => n6608, QN => n180);
   registers_reg_14_11_inst : HS65_LH_DFPRQNX9 port map( D => n1861, CP => clk,
                           RN => n6608, QN => n181);
   registers_reg_14_10_inst : HS65_LH_DFPRQNX9 port map( D => n1860, CP => clk,
                           RN => n6608, QN => n182);
   registers_reg_14_9_inst : HS65_LH_DFPRQNX9 port map( D => n1859, CP => clk, 
                           RN => n6608, QN => n183);
   registers_reg_14_8_inst : HS65_LH_DFPRQNX9 port map( D => n1858, CP => clk, 
                           RN => n6608, QN => n184);
   registers_reg_14_7_inst : HS65_LH_DFPRQNX9 port map( D => n1857, CP => clk, 
                           RN => n6607, QN => n185);
   registers_reg_14_6_inst : HS65_LH_DFPRQNX9 port map( D => n1856, CP => clk, 
                           RN => n6607, QN => n186);
   registers_reg_14_5_inst : HS65_LH_DFPRQNX9 port map( D => n1855, CP => clk, 
                           RN => n6607, QN => n187);
   registers_reg_14_4_inst : HS65_LH_DFPRQNX9 port map( D => n1854, CP => clk, 
                           RN => n6607, QN => n188);
   registers_reg_14_3_inst : HS65_LH_DFPRQNX9 port map( D => n1853, CP => clk, 
                           RN => n6607, QN => n189);
   registers_reg_14_2_inst : HS65_LH_DFPRQNX9 port map( D => n1852, CP => clk, 
                           RN => n6607, QN => n190);
   registers_reg_14_1_inst : HS65_LH_DFPRQNX9 port map( D => n1851, CP => clk, 
                           RN => n6607, QN => n191);
   registers_reg_14_0_inst : HS65_LH_DFPRQNX9 port map( D => n1850, CP => clk, 
                           RN => n6607, QN => n192);
   registers_reg_26_31_inst : HS65_LH_DFPRQNX9 port map( D => n2265, CP => clk,
                           RN => n6607, QN => n97);
   registers_reg_26_30_inst : HS65_LH_DFPRQNX9 port map( D => n2264, CP => clk,
                           RN => n6607, QN => n98);
   registers_reg_26_29_inst : HS65_LH_DFPRQNX9 port map( D => n2263, CP => clk,
                           RN => n6607, QN => n99);
   registers_reg_26_28_inst : HS65_LH_DFPRQNX9 port map( D => n2262, CP => clk,
                           RN => n6607, QN => n100);
   registers_reg_26_27_inst : HS65_LH_DFPRQNX9 port map( D => n2261, CP => clk,
                           RN => n6607, QN => n101);
   registers_reg_26_26_inst : HS65_LH_DFPRQNX9 port map( D => n2260, CP => clk,
                           RN => n6607, QN => n102);
   registers_reg_26_25_inst : HS65_LH_DFPRQNX9 port map( D => n2259, CP => clk,
                           RN => n6606, QN => n103);
   registers_reg_26_24_inst : HS65_LH_DFPRQNX9 port map( D => n2258, CP => clk,
                           RN => n6606, QN => n104);
   registers_reg_26_23_inst : HS65_LH_DFPRQNX9 port map( D => n2257, CP => clk,
                           RN => n6606, QN => n105);
   registers_reg_26_22_inst : HS65_LH_DFPRQNX9 port map( D => n2256, CP => clk,
                           RN => n6606, QN => n106);
   registers_reg_26_21_inst : HS65_LH_DFPRQNX9 port map( D => n2255, CP => clk,
                           RN => n6606, QN => n107);
   registers_reg_26_20_inst : HS65_LH_DFPRQNX9 port map( D => n2254, CP => clk,
                           RN => n6606, QN => n108);
   registers_reg_26_19_inst : HS65_LH_DFPRQNX9 port map( D => n2253, CP => clk,
                           RN => n6606, QN => n109);
   registers_reg_26_18_inst : HS65_LH_DFPRQNX9 port map( D => n2252, CP => clk,
                           RN => n6606, QN => n110);
   registers_reg_26_17_inst : HS65_LH_DFPRQNX9 port map( D => n2251, CP => clk,
                           RN => n6606, QN => n111);
   registers_reg_26_16_inst : HS65_LH_DFPRQNX9 port map( D => n2250, CP => clk,
                           RN => n6606, QN => n112);
   registers_reg_26_15_inst : HS65_LH_DFPRQNX9 port map( D => n2249, CP => clk,
                           RN => n6606, QN => n113);
   registers_reg_26_14_inst : HS65_LH_DFPRQNX9 port map( D => n2248, CP => clk,
                           RN => n6606, QN => n114);
   registers_reg_26_13_inst : HS65_LH_DFPRQNX9 port map( D => n2247, CP => clk,
                           RN => n6606, QN => n115);
   registers_reg_26_12_inst : HS65_LH_DFPRQNX9 port map( D => n2246, CP => clk,
                           RN => n6606, QN => n116);
   registers_reg_26_11_inst : HS65_LH_DFPRQNX9 port map( D => n2245, CP => clk,
                           RN => n6605, QN => n117);
   registers_reg_26_10_inst : HS65_LH_DFPRQNX9 port map( D => n2244, CP => clk,
                           RN => n6605, QN => n118);
   registers_reg_26_9_inst : HS65_LH_DFPRQNX9 port map( D => n2243, CP => clk, 
                           RN => n6605, QN => n119);
   registers_reg_26_8_inst : HS65_LH_DFPRQNX9 port map( D => n2242, CP => clk, 
                           RN => n6605, QN => n120);
   registers_reg_26_7_inst : HS65_LH_DFPRQNX9 port map( D => n2241, CP => clk, 
                           RN => n6605, QN => n121);
   registers_reg_26_6_inst : HS65_LH_DFPRQNX9 port map( D => n2240, CP => clk, 
                           RN => n6605, QN => n122);
   registers_reg_26_5_inst : HS65_LH_DFPRQNX9 port map( D => n2239, CP => clk, 
                           RN => n6605, QN => n123);
   registers_reg_26_4_inst : HS65_LH_DFPRQNX9 port map( D => n2238, CP => clk, 
                           RN => n6605, QN => n124);
   registers_reg_26_3_inst : HS65_LH_DFPRQNX9 port map( D => n2237, CP => clk, 
                           RN => n6605, QN => n125);
   registers_reg_26_2_inst : HS65_LH_DFPRQNX9 port map( D => n2236, CP => clk, 
                           RN => n6605, QN => n126);
   registers_reg_26_1_inst : HS65_LH_DFPRQNX9 port map( D => n2235, CP => clk, 
                           RN => n6605, QN => n127);
   registers_reg_26_0_inst : HS65_LH_DFPRQNX9 port map( D => n2234, CP => clk, 
                           RN => n6605, QN => n128);
   registers_reg_29_31_inst : HS65_LH_DFPRQNX9 port map( D => n2361, CP => clk,
                           RN => n6605, QN => n1);
   registers_reg_29_30_inst : HS65_LH_DFPRQNX9 port map( D => n2360, CP => clk,
                           RN => n6605, QN => n2);
   registers_reg_29_29_inst : HS65_LH_DFPRQNX9 port map( D => n2359, CP => clk,
                           RN => n6604, QN => n3);
   registers_reg_29_28_inst : HS65_LH_DFPRQNX9 port map( D => n2358, CP => clk,
                           RN => n6604, QN => n4);
   registers_reg_29_27_inst : HS65_LH_DFPRQNX9 port map( D => n2357, CP => clk,
                           RN => n6604, QN => n5);
   registers_reg_29_26_inst : HS65_LH_DFPRQNX9 port map( D => n2356, CP => clk,
                           RN => n6604, QN => n6);
   registers_reg_29_25_inst : HS65_LH_DFPRQNX9 port map( D => n2355, CP => clk,
                           RN => n6604, QN => n7);
   registers_reg_29_24_inst : HS65_LH_DFPRQNX9 port map( D => n2354, CP => clk,
                           RN => n6604, QN => n8);
   registers_reg_29_23_inst : HS65_LH_DFPRQNX9 port map( D => n2353, CP => clk,
                           RN => n6604, QN => n9);
   registers_reg_29_22_inst : HS65_LH_DFPRQNX9 port map( D => n2352, CP => clk,
                           RN => n6604, QN => n10);
   registers_reg_29_21_inst : HS65_LH_DFPRQNX9 port map( D => n2351, CP => clk,
                           RN => n6604, QN => n11);
   registers_reg_29_20_inst : HS65_LH_DFPRQNX9 port map( D => n2350, CP => clk,
                           RN => n6604, QN => n12);
   registers_reg_29_19_inst : HS65_LH_DFPRQNX9 port map( D => n2349, CP => clk,
                           RN => n6604, QN => n13);
   registers_reg_29_18_inst : HS65_LH_DFPRQNX9 port map( D => n2348, CP => clk,
                           RN => n6604, QN => n14);
   registers_reg_29_17_inst : HS65_LH_DFPRQNX9 port map( D => n2347, CP => clk,
                           RN => n6604, QN => n15);
   registers_reg_29_16_inst : HS65_LH_DFPRQNX9 port map( D => n2346, CP => clk,
                           RN => n6604, QN => n16);
   registers_reg_29_15_inst : HS65_LH_DFPRQNX9 port map( D => n2345, CP => clk,
                           RN => n6603, QN => n17);
   registers_reg_29_14_inst : HS65_LH_DFPRQNX9 port map( D => n2344, CP => clk,
                           RN => n6603, QN => n18);
   registers_reg_29_13_inst : HS65_LH_DFPRQNX9 port map( D => n2343, CP => clk,
                           RN => n6603, QN => n19);
   registers_reg_29_12_inst : HS65_LH_DFPRQNX9 port map( D => n2342, CP => clk,
                           RN => n6603, QN => n20);
   registers_reg_29_11_inst : HS65_LH_DFPRQNX9 port map( D => n2341, CP => clk,
                           RN => n6603, QN => n21);
   registers_reg_29_10_inst : HS65_LH_DFPRQNX9 port map( D => n2340, CP => clk,
                           RN => n6603, QN => n22);
   registers_reg_29_9_inst : HS65_LH_DFPRQNX9 port map( D => n2339, CP => clk, 
                           RN => n6603, QN => n23);
   registers_reg_29_8_inst : HS65_LH_DFPRQNX9 port map( D => n2338, CP => clk, 
                           RN => n6603, QN => n24);
   registers_reg_29_7_inst : HS65_LH_DFPRQNX9 port map( D => n2337, CP => clk, 
                           RN => n6603, QN => n25);
   registers_reg_29_6_inst : HS65_LH_DFPRQNX9 port map( D => n2336, CP => clk, 
                           RN => n6603, QN => n26);
   registers_reg_29_5_inst : HS65_LH_DFPRQNX9 port map( D => n2335, CP => clk, 
                           RN => n6603, QN => n27);
   registers_reg_29_4_inst : HS65_LH_DFPRQNX9 port map( D => n2334, CP => clk, 
                           RN => n6603, QN => n28);
   registers_reg_29_3_inst : HS65_LH_DFPRQNX9 port map( D => n2333, CP => clk, 
                           RN => n6603, QN => n29);
   registers_reg_29_2_inst : HS65_LH_DFPRQNX9 port map( D => n2332, CP => clk, 
                           RN => n6603, QN => n30);
   registers_reg_29_1_inst : HS65_LH_DFPRQNX9 port map( D => n2331, CP => clk, 
                           RN => n6602, QN => n31);
   registers_reg_29_0_inst : HS65_LH_DFPRQNX9 port map( D => n2330, CP => clk, 
                           RN => n6602, QN => n32);
   registers_reg_8_31_inst : HS65_LH_DFPRQNX9 port map( D => n1689, CP => clk, 
                           RN => n6600, QN => n225);
   registers_reg_8_30_inst : HS65_LH_DFPRQNX9 port map( D => n1688, CP => clk, 
                           RN => n6600, QN => n226);
   registers_reg_8_29_inst : HS65_LH_DFPRQNX9 port map( D => n1687, CP => clk, 
                           RN => n6600, QN => n227);
   registers_reg_8_28_inst : HS65_LH_DFPRQNX9 port map( D => n1686, CP => clk, 
                           RN => n6600, QN => n228);
   registers_reg_8_27_inst : HS65_LH_DFPRQNX9 port map( D => n1685, CP => clk, 
                           RN => n6600, QN => n229);
   registers_reg_8_26_inst : HS65_LH_DFPRQNX9 port map( D => n1684, CP => clk, 
                           RN => n6600, QN => n230);
   registers_reg_8_25_inst : HS65_LH_DFPRQNX9 port map( D => n1683, CP => clk, 
                           RN => n6600, QN => n231);
   registers_reg_8_24_inst : HS65_LH_DFPRQNX9 port map( D => n1682, CP => clk, 
                           RN => n6600, QN => n232);
   registers_reg_8_23_inst : HS65_LH_DFPRQNX9 port map( D => n1681, CP => clk, 
                           RN => n6599, QN => n233);
   registers_reg_8_22_inst : HS65_LH_DFPRQNX9 port map( D => n1680, CP => clk, 
                           RN => n6599, QN => n234);
   registers_reg_8_21_inst : HS65_LH_DFPRQNX9 port map( D => n1679, CP => clk, 
                           RN => n6599, QN => n235);
   registers_reg_8_20_inst : HS65_LH_DFPRQNX9 port map( D => n1678, CP => clk, 
                           RN => n6599, QN => n236);
   registers_reg_8_19_inst : HS65_LH_DFPRQNX9 port map( D => n1677, CP => clk, 
                           RN => n6599, QN => n237);
   registers_reg_8_18_inst : HS65_LH_DFPRQNX9 port map( D => n1676, CP => clk, 
                           RN => n6599, QN => n238);
   registers_reg_8_17_inst : HS65_LH_DFPRQNX9 port map( D => n1675, CP => clk, 
                           RN => n6599, QN => n239);
   registers_reg_8_16_inst : HS65_LH_DFPRQNX9 port map( D => n1674, CP => clk, 
                           RN => n6599, QN => n240);
   registers_reg_8_15_inst : HS65_LH_DFPRQNX9 port map( D => n1673, CP => clk, 
                           RN => n6599, QN => n241);
   registers_reg_8_14_inst : HS65_LH_DFPRQNX9 port map( D => n1672, CP => clk, 
                           RN => n6599, QN => n242);
   registers_reg_8_13_inst : HS65_LH_DFPRQNX9 port map( D => n1671, CP => clk, 
                           RN => n6599, QN => n243);
   registers_reg_8_12_inst : HS65_LH_DFPRQNX9 port map( D => n1670, CP => clk, 
                           RN => n6599, QN => n244);
   registers_reg_8_11_inst : HS65_LH_DFPRQNX9 port map( D => n1669, CP => clk, 
                           RN => n6599, QN => n245);
   registers_reg_8_10_inst : HS65_LH_DFPRQNX9 port map( D => n1668, CP => clk, 
                           RN => n6599, QN => n246);
   registers_reg_8_9_inst : HS65_LH_DFPRQNX9 port map( D => n1667, CP => clk, 
                           RN => n6598, QN => n247);
   registers_reg_8_8_inst : HS65_LH_DFPRQNX9 port map( D => n1666, CP => clk, 
                           RN => n6598, QN => n248);
   registers_reg_8_7_inst : HS65_LH_DFPRQNX9 port map( D => n1665, CP => clk, 
                           RN => n6598, QN => n249);
   registers_reg_8_6_inst : HS65_LH_DFPRQNX9 port map( D => n1664, CP => clk, 
                           RN => n6598, QN => n250);
   registers_reg_8_5_inst : HS65_LH_DFPRQNX9 port map( D => n1663, CP => clk, 
                           RN => n6598, QN => n251);
   registers_reg_8_4_inst : HS65_LH_DFPRQNX9 port map( D => n1662, CP => clk, 
                           RN => n6598, QN => n252);
   registers_reg_8_3_inst : HS65_LH_DFPRQNX9 port map( D => n1661, CP => clk, 
                           RN => n6598, QN => n253);
   registers_reg_8_2_inst : HS65_LH_DFPRQNX9 port map( D => n1660, CP => clk, 
                           RN => n6598, QN => n254);
   registers_reg_8_1_inst : HS65_LH_DFPRQNX9 port map( D => n1659, CP => clk, 
                           RN => n6598, QN => n255);
   registers_reg_8_0_inst : HS65_LH_DFPRQNX9 port map( D => n1658, CP => clk, 
                           RN => n6598, QN => n256);
   registers_reg_15_31_inst : HS65_LH_DFPRQNX9 port map( D => n1913, CP => clk,
                           RN => n6614, QN => n129);
   registers_reg_15_30_inst : HS65_LH_DFPRQNX9 port map( D => n1912, CP => clk,
                           RN => n6614, QN => n130);
   registers_reg_15_29_inst : HS65_LH_DFPRQNX9 port map( D => n1911, CP => clk,
                           RN => n6614, QN => n131);
   registers_reg_15_28_inst : HS65_LH_DFPRQNX9 port map( D => n1910, CP => clk,
                           RN => n6614, QN => n132);
   registers_reg_15_27_inst : HS65_LH_DFPRQNX9 port map( D => n1909, CP => clk,
                           RN => n6613, QN => n133);
   registers_reg_15_26_inst : HS65_LH_DFPRQNX9 port map( D => n1908, CP => clk,
                           RN => n6613, QN => n134);
   registers_reg_15_25_inst : HS65_LH_DFPRQNX9 port map( D => n1907, CP => clk,
                           RN => n6613, QN => n135);
   registers_reg_15_24_inst : HS65_LH_DFPRQNX9 port map( D => n1906, CP => clk,
                           RN => n6613, QN => n136);
   registers_reg_15_23_inst : HS65_LH_DFPRQNX9 port map( D => n1905, CP => clk,
                           RN => n6613, QN => n137);
   registers_reg_15_22_inst : HS65_LH_DFPRQNX9 port map( D => n1904, CP => clk,
                           RN => n6613, QN => n138);
   registers_reg_15_21_inst : HS65_LH_DFPRQNX9 port map( D => n1903, CP => clk,
                           RN => n6613, QN => n139);
   registers_reg_15_20_inst : HS65_LH_DFPRQNX9 port map( D => n1902, CP => clk,
                           RN => n6613, QN => n140);
   registers_reg_15_19_inst : HS65_LH_DFPRQNX9 port map( D => n1901, CP => clk,
                           RN => n6613, QN => n141);
   registers_reg_15_18_inst : HS65_LH_DFPRQNX9 port map( D => n1900, CP => clk,
                           RN => n6613, QN => n142);
   registers_reg_15_17_inst : HS65_LH_DFPRQNX9 port map( D => n1899, CP => clk,
                           RN => n6613, QN => n143);
   registers_reg_15_16_inst : HS65_LH_DFPRQNX9 port map( D => n1898, CP => clk,
                           RN => n6613, QN => n144);
   registers_reg_15_15_inst : HS65_LH_DFPRQNX9 port map( D => n1897, CP => clk,
                           RN => n6613, QN => n145);
   registers_reg_15_14_inst : HS65_LH_DFPRQNX9 port map( D => n1896, CP => clk,
                           RN => n6613, QN => n146);
   registers_reg_15_13_inst : HS65_LH_DFPRQNX9 port map( D => n1895, CP => clk,
                           RN => n6612, QN => n147);
   registers_reg_15_12_inst : HS65_LH_DFPRQNX9 port map( D => n1894, CP => clk,
                           RN => n6612, QN => n148);
   registers_reg_15_11_inst : HS65_LH_DFPRQNX9 port map( D => n1893, CP => clk,
                           RN => n6612, QN => n149);
   registers_reg_15_10_inst : HS65_LH_DFPRQNX9 port map( D => n1892, CP => clk,
                           RN => n6612, QN => n150);
   registers_reg_15_9_inst : HS65_LH_DFPRQNX9 port map( D => n1891, CP => clk, 
                           RN => n6612, QN => n151);
   registers_reg_15_8_inst : HS65_LH_DFPRQNX9 port map( D => n1890, CP => clk, 
                           RN => n6612, QN => n152);
   registers_reg_15_7_inst : HS65_LH_DFPRQNX9 port map( D => n1889, CP => clk, 
                           RN => n6612, QN => n153);
   registers_reg_15_6_inst : HS65_LH_DFPRQNX9 port map( D => n1888, CP => clk, 
                           RN => n6612, QN => n154);
   registers_reg_15_5_inst : HS65_LH_DFPRQNX9 port map( D => n1887, CP => clk, 
                           RN => n6612, QN => n155);
   registers_reg_15_4_inst : HS65_LH_DFPRQNX9 port map( D => n1886, CP => clk, 
                           RN => n6612, QN => n156);
   registers_reg_15_3_inst : HS65_LH_DFPRQNX9 port map( D => n1885, CP => clk, 
                           RN => n6612, QN => n157);
   registers_reg_15_2_inst : HS65_LH_DFPRQNX9 port map( D => n1884, CP => clk, 
                           RN => n6612, QN => n158);
   registers_reg_15_1_inst : HS65_LH_DFPRQNX9 port map( D => n1883, CP => clk, 
                           RN => n6612, QN => n159);
   registers_reg_15_0_inst : HS65_LH_DFPRQNX9 port map( D => n1882, CP => clk, 
                           RN => n6612, QN => n160);
   registers_reg_9_31_inst : HS65_LH_DFPRQNX9 port map( D => n1721, CP => clk, 
                           RN => n6602, QN => n193);
   registers_reg_9_30_inst : HS65_LH_DFPRQNX9 port map( D => n1720, CP => clk, 
                           RN => n6602, QN => n194);
   registers_reg_9_29_inst : HS65_LH_DFPRQNX9 port map( D => n1719, CP => clk, 
                           RN => n6602, QN => n195);
   registers_reg_9_28_inst : HS65_LH_DFPRQNX9 port map( D => n1718, CP => clk, 
                           RN => n6602, QN => n196);
   registers_reg_9_27_inst : HS65_LH_DFPRQNX9 port map( D => n1717, CP => clk, 
                           RN => n6602, QN => n197);
   registers_reg_9_26_inst : HS65_LH_DFPRQNX9 port map( D => n1716, CP => clk, 
                           RN => n6602, QN => n198);
   registers_reg_9_25_inst : HS65_LH_DFPRQNX9 port map( D => n1715, CP => clk, 
                           RN => n6602, QN => n199);
   registers_reg_9_24_inst : HS65_LH_DFPRQNX9 port map( D => n1714, CP => clk, 
                           RN => n6602, QN => n200);
   registers_reg_9_23_inst : HS65_LH_DFPRQNX9 port map( D => n1713, CP => clk, 
                           RN => n6602, QN => n201);
   registers_reg_9_22_inst : HS65_LH_DFPRQNX9 port map( D => n1712, CP => clk, 
                           RN => n6602, QN => n202);
   registers_reg_9_21_inst : HS65_LH_DFPRQNX9 port map( D => n1711, CP => clk, 
                           RN => n6602, QN => n203);
   registers_reg_9_20_inst : HS65_LH_DFPRQNX9 port map( D => n1710, CP => clk, 
                           RN => n6602, QN => n204);
   registers_reg_9_19_inst : HS65_LH_DFPRQNX9 port map( D => n1709, CP => clk, 
                           RN => n6601, QN => n205);
   registers_reg_9_18_inst : HS65_LH_DFPRQNX9 port map( D => n1708, CP => clk, 
                           RN => n6601, QN => n206);
   registers_reg_9_17_inst : HS65_LH_DFPRQNX9 port map( D => n1707, CP => clk, 
                           RN => n6601, QN => n207);
   registers_reg_9_16_inst : HS65_LH_DFPRQNX9 port map( D => n1706, CP => clk, 
                           RN => n6601, QN => n208);
   registers_reg_9_15_inst : HS65_LH_DFPRQNX9 port map( D => n1705, CP => clk, 
                           RN => n6601, QN => n209);
   registers_reg_9_14_inst : HS65_LH_DFPRQNX9 port map( D => n1704, CP => clk, 
                           RN => n6601, QN => n210);
   registers_reg_9_13_inst : HS65_LH_DFPRQNX9 port map( D => n1703, CP => clk, 
                           RN => n6601, QN => n211);
   registers_reg_9_12_inst : HS65_LH_DFPRQNX9 port map( D => n1702, CP => clk, 
                           RN => n6601, QN => n212);
   registers_reg_9_11_inst : HS65_LH_DFPRQNX9 port map( D => n1701, CP => clk, 
                           RN => n6601, QN => n213);
   registers_reg_9_10_inst : HS65_LH_DFPRQNX9 port map( D => n1700, CP => clk, 
                           RN => n6601, QN => n214);
   registers_reg_9_9_inst : HS65_LH_DFPRQNX9 port map( D => n1699, CP => clk, 
                           RN => n6601, QN => n215);
   registers_reg_9_8_inst : HS65_LH_DFPRQNX9 port map( D => n1698, CP => clk, 
                           RN => n6601, QN => n216);
   registers_reg_9_7_inst : HS65_LH_DFPRQNX9 port map( D => n1697, CP => clk, 
                           RN => n6601, QN => n217);
   registers_reg_9_6_inst : HS65_LH_DFPRQNX9 port map( D => n1696, CP => clk, 
                           RN => n6601, QN => n218);
   registers_reg_9_5_inst : HS65_LH_DFPRQNX9 port map( D => n1695, CP => clk, 
                           RN => n6600, QN => n219);
   registers_reg_9_4_inst : HS65_LH_DFPRQNX9 port map( D => n1694, CP => clk, 
                           RN => n6600, QN => n220);
   registers_reg_9_3_inst : HS65_LH_DFPRQNX9 port map( D => n1693, CP => clk, 
                           RN => n6600, QN => n221);
   registers_reg_9_2_inst : HS65_LH_DFPRQNX9 port map( D => n1692, CP => clk, 
                           RN => n6600, QN => n222);
   registers_reg_9_1_inst : HS65_LH_DFPRQNX9 port map( D => n1691, CP => clk, 
                           RN => n6600, QN => n223);
   registers_reg_9_0_inst : HS65_LH_DFPRQNX9 port map( D => n1690, CP => clk, 
                           RN => n6600, QN => n224);
   U3 : HS65_LH_AND2X4 port map( A => n2824, B => n2825, Z => n6167);
   U4 : HS65_LH_AND2X4 port map( A => n2827, B => n2825, Z => n6168);
   U5 : HS65_LH_AND2X4 port map( A => n2850, B => n2829, Z => n6169);
   U6 : HS65_LH_AND2X4 port map( A => n2850, B => n2833, Z => n6170);
   U7 : HS65_LH_AND2X4 port map( A => n2841, B => n2833, Z => n6171);
   U8 : HS65_LH_AND2X4 port map( A => n2841, B => n2831, Z => n6172);
   U9 : HS65_LH_AND2X4 port map( A => n2841, B => n2829, Z => n6173);
   U10 : HS65_LH_AND2X4 port map( A => n2841, B => n2824, Z => n6174);
   U11 : HS65_LH_AND2X4 port map( A => n2841, B => n2827, Z => n6175);
   U12 : HS65_LH_AND2X4 port map( A => n2859, B => n2831, Z => n6176);
   U13 : HS65_LH_AND2X4 port map( A => n2859, B => n2833, Z => n6177);
   U14 : HS65_LH_AND2X4 port map( A => n2859, B => n2835, Z => n6178);
   U15 : HS65_LH_AND2X4 port map( A => n2859, B => n2829, Z => n6179);
   U16 : HS65_LH_AND2X4 port map( A => n2859, B => n2837, Z => n6180);
   U17 : HS65_LH_AND2X4 port map( A => n2859, B => n2824, Z => n6181);
   U18 : HS65_LH_AND2X4 port map( A => n1323, B => n1330, Z => n882);
   U19 : HS65_LH_AND2X4 port map( A => n2806, B => n2819, Z => n1373);
   U20 : HS65_LH_AND2X4 port map( A => n1322, B => n1327, Z => n862);
   U21 : HS65_LH_AND2X4 port map( A => n1326, B => n1327, Z => n857);
   U22 : HS65_LH_AND2X4 port map( A => n1329, B => n1327, Z => n868);
   U23 : HS65_LH_AND2X4 port map( A => n1329, B => n1323, Z => n870);
   U24 : HS65_LH_AND2X4 port map( A => n1326, B => n1323, Z => n866);
   U25 : HS65_LH_AND2X4 port map( A => n1324, B => n1323, Z => n865);
   U26 : HS65_LH_AND2X4 port map( A => n2822, B => n2806, Z => n1381);
   U27 : HS65_LH_AND2X4 port map( A => n2810, B => n2806, Z => n1354);
   U28 : HS65_LH_AND2X4 port map( A => n2813, B => n2806, Z => n1359);
   U29 : HS65_LH_AND2X4 port map( A => n2811, B => n2806, Z => n1355);
   U30 : HS65_LH_AND2X4 port map( A => n2811, B => n2808, Z => n1353);
   U31 : HS65_LH_AND2X4 port map( A => n2805, B => n2808, Z => n1348);
   U32 : HS65_LH_AND2X4 port map( A => n2813, B => n2808, Z => n1357);
   U33 : HS65_LH_AND2X4 port map( A => n2810, B => n2808, Z => n1356);
   U34 : HS65_LH_AND2X4 port map( A => n1330, B => n1325, Z => n881);
   U35 : HS65_LH_AND2X4 port map( A => n1338, B => n1325, Z => n888);
   U36 : HS65_LH_AND2X4 port map( A => n1331, B => n1325, Z => n892);
   U37 : HS65_LH_AND2X4 port map( A => n1329, B => n1325, Z => n871);
   U38 : HS65_LH_AND2X4 port map( A => n1326, B => n1325, Z => n869);
   U39 : HS65_LH_AND2X4 port map( A => n1322, B => n1325, Z => n864);
   U40 : HS65_LH_AND2X4 port map( A => n2805, B => n2812, Z => n1352);
   U41 : HS65_LH_AND2X4 port map( A => n2813, B => n2812, Z => n1361);
   U42 : HS65_LH_AND2X4 port map( A => n2810, B => n2812, Z => n1360);
   U43 : HS65_LH_AND2X4 port map( A => n2812, B => n2822, Z => n1380);
   U44 : HS65_LH_AND2X4 port map( A => n2820, B => n2807, Z => n1367);
   U45 : HS65_LH_AND2X4 port map( A => n2813, B => n2807, Z => n1362);
   U46 : HS65_LH_AND2X4 port map( A => n2811, B => n2807, Z => n1358);
   U47 : HS65_LH_AND2X4 port map( A => n1324, B => n1328, Z => n886);
   U48 : HS65_LH_AND2X4 port map( A => n1329, B => n1328, Z => n863);
   U49 : HS65_LH_AND2X4 port map( A => n1326, B => n1328, Z => n856);
   U50 : HS65_LH_AND2X4 port map( A => n1327, B => n1331, Z => n891);
   U51 : HS65_LH_AND2X4 port map( A => n1327, B => n1330, Z => n861);
   U52 : HS65_LH_AND2X4 port map( A => n1323, B => n1331, Z => n867);
   U53 : HS65_LH_AND2X4 port map( A => n2808, B => n2819, Z => n1372);
   U54 : HS65_LH_AND2X4 port map( A => n2812, B => n2809, Z => n1379);
   U55 : HS65_LH_AND2X4 port map( A => n2812, B => n2819, Z => n1377);
   U56 : HS65_LH_AND2X4 port map( A => n2806, B => n2809, Z => n1378);
   U57 : HS65_LH_AND2X4 port map( A => n2808, B => n2809, Z => n1347);
   U58 : HS65_LH_AND2X4 port map( A => n1325, B => n1337, Z => n876);
   U59 : HS65_LH_AND2X4 port map( A => n1327, B => n1337, Z => n889);
   U60 : HS65_LH_AND2X4 port map( A => n1323, B => n1337, Z => n890);
   U61 : HS65_LH_AND2X4 port map( A => n2812, B => n2811, Z => n1384);
   U62 : HS65_LH_AND2X4 port map( A => n1328, B => n1338, Z => n877);
   U63 : HS65_LH_AND2X4 port map( A => n1323, B => n1338, Z => n887);
   U64 : HS65_LH_AND2X4 port map( A => n1327, B => n1338, Z => n893);
   U65 : HS65_LH_AND2X4 port map( A => n2808, B => n2820, Z => n1368);
   U66 : HS65_LH_AND2X4 port map( A => n2806, B => n2820, Z => n1383);
   U67 : HS65_LH_AND2X4 port map( A => n2812, B => n2820, Z => n1382);
   U68 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => n795, C => 
                           regfile_i(38), Z => n2841);
   U69 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => n811, C => 
                           regfile_i(39), Z => n2850);
   U70 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => n795, C => n811, Z 
                           => n2825);
   U71 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => regfile_i(38), C => 
                           regfile_i(39), Z => n2859);
   U72 : HS65_LH_IVX9 port map( A => regfile_i(1), Z => n848);
   U73 : HS65_LH_IVX9 port map( A => regfile_i(2), Z => n847);
   U74 : HS65_LH_BFX9 port map( A => n6626, Z => n6598);
   U75 : HS65_LH_BFX9 port map( A => n6625, Z => n6599);
   U76 : HS65_LH_BFX9 port map( A => n6625, Z => n6600);
   U77 : HS65_LH_BFX9 port map( A => n6624, Z => n6601);
   U78 : HS65_LH_BFX9 port map( A => n6624, Z => n6602);
   U79 : HS65_LH_BFX9 port map( A => n6623, Z => n6603);
   U80 : HS65_LH_BFX9 port map( A => n6623, Z => n6604);
   U81 : HS65_LH_BFX9 port map( A => n6622, Z => n6605);
   U82 : HS65_LH_BFX9 port map( A => n6622, Z => n6606);
   U83 : HS65_LH_BFX9 port map( A => n6621, Z => n6607);
   U84 : HS65_LH_BFX9 port map( A => n6621, Z => n6608);
   U85 : HS65_LH_BFX9 port map( A => n6620, Z => n6609);
   U86 : HS65_LH_BFX9 port map( A => n6620, Z => n6610);
   U87 : HS65_LH_BFX9 port map( A => n6619, Z => n6611);
   U88 : HS65_LH_BFX9 port map( A => n6619, Z => n6612);
   U89 : HS65_LH_BFX9 port map( A => n6618, Z => n6613);
   U90 : HS65_LH_BFX9 port map( A => n6618, Z => n6614);
   U91 : HS65_LH_BFX9 port map( A => n6617, Z => n6615);
   U92 : HS65_LH_BFX9 port map( A => n6634, Z => n6581);
   U93 : HS65_LH_BFX9 port map( A => n6637, Z => n6575);
   U94 : HS65_LH_BFX9 port map( A => n6651, Z => n6547);
   U95 : HS65_LH_BFX9 port map( A => n6653, Z => n6543);
   U96 : HS65_LH_BFX9 port map( A => n6642, Z => n6566);
   U97 : HS65_LH_BFX9 port map( A => n6641, Z => n6567);
   U98 : HS65_LH_BFX9 port map( A => n6642, Z => n6565);
   U99 : HS65_LH_BFX9 port map( A => n6656, Z => n6537);
   U100 : HS65_LH_BFX9 port map( A => n6643, Z => n6564);
   U101 : HS65_LH_BFX9 port map( A => n6643, Z => n6563);
   U102 : HS65_LH_BFX9 port map( A => n6649, Z => n6551);
   U103 : HS65_LH_BFX9 port map( A => n6650, Z => n6549);
   U104 : HS65_LH_BFX9 port map( A => n6652, Z => n6546);
   U105 : HS65_LH_BFX9 port map( A => n6652, Z => n6545);
   U106 : HS65_LH_BFX9 port map( A => n6653, Z => n6544);
   U107 : HS65_LH_BFX9 port map( A => n6644, Z => n6562);
   U108 : HS65_LH_BFX9 port map( A => n6645, Z => n6560);
   U109 : HS65_LH_BFX9 port map( A => n6644, Z => n6561);
   U110 : HS65_LH_BFX9 port map( A => n6645, Z => n6559);
   U111 : HS65_LH_BFX9 port map( A => n6648, Z => n6554);
   U112 : HS65_LH_BFX9 port map( A => n6648, Z => n6553);
   U113 : HS65_LH_BFX9 port map( A => n6646, Z => n6558);
   U114 : HS65_LH_BFX9 port map( A => n6647, Z => n6556);
   U115 : HS65_LH_BFX9 port map( A => n6646, Z => n6557);
   U116 : HS65_LH_BFX9 port map( A => n6647, Z => n6555);
   U117 : HS65_LH_BFX9 port map( A => n6649, Z => n6552);
   U118 : HS65_LH_BFX9 port map( A => n6650, Z => n6550);
   U119 : HS65_LH_BFX9 port map( A => n6651, Z => n6548);
   U120 : HS65_LH_BFX9 port map( A => n6631, Z => n6587);
   U121 : HS65_LH_BFX9 port map( A => n6636, Z => n6577);
   U122 : HS65_LH_BFX9 port map( A => n6637, Z => n6576);
   U123 : HS65_LH_BFX9 port map( A => n6638, Z => n6574);
   U124 : HS65_LH_BFX9 port map( A => n6638, Z => n6573);
   U125 : HS65_LH_BFX9 port map( A => n6655, Z => n6540);
   U126 : HS65_LH_BFX9 port map( A => n6654, Z => n6542);
   U127 : HS65_LH_BFX9 port map( A => n6654, Z => n6541);
   U128 : HS65_LH_BFX9 port map( A => n6656, Z => n6538);
   U129 : HS65_LH_BFX9 port map( A => n6626, Z => n6597);
   U130 : HS65_LH_BFX9 port map( A => n6627, Z => n6596);
   U131 : HS65_LH_BFX9 port map( A => n6627, Z => n6595);
   U132 : HS65_LH_BFX9 port map( A => n6628, Z => n6594);
   U133 : HS65_LH_BFX9 port map( A => n6628, Z => n6593);
   U134 : HS65_LH_BFX9 port map( A => n6629, Z => n6592);
   U135 : HS65_LH_BFX9 port map( A => n6630, Z => n6590);
   U136 : HS65_LH_BFX9 port map( A => n6629, Z => n6591);
   U137 : HS65_LH_BFX9 port map( A => n6631, Z => n6588);
   U138 : HS65_LH_BFX9 port map( A => n6630, Z => n6589);
   U139 : HS65_LH_BFX9 port map( A => n6632, Z => n6586);
   U140 : HS65_LH_BFX9 port map( A => n6634, Z => n6582);
   U141 : HS65_LH_BFX9 port map( A => n6632, Z => n6585);
   U142 : HS65_LH_BFX9 port map( A => n6635, Z => n6579);
   U143 : HS65_LH_BFX9 port map( A => n6633, Z => n6584);
   U144 : HS65_LH_BFX9 port map( A => n6633, Z => n6583);
   U145 : HS65_LH_BFX9 port map( A => n6635, Z => n6580);
   U146 : HS65_LH_BFX9 port map( A => n6636, Z => n6578);
   U147 : HS65_LH_BFX9 port map( A => n6641, Z => n6568);
   U148 : HS65_LH_BFX9 port map( A => n6639, Z => n6572);
   U149 : HS65_LH_BFX9 port map( A => n6640, Z => n6570);
   U150 : HS65_LH_BFX9 port map( A => n6639, Z => n6571);
   U151 : HS65_LH_BFX9 port map( A => n6640, Z => n6569);
   U152 : HS65_LH_BFX9 port map( A => n6655, Z => n6539);
   U153 : HS65_LH_BFX9 port map( A => n6617, Z => n6616);
   U154 : HS65_LH_IVX9 port map( A => n6239, Z => n6238);
   U155 : HS65_LH_IVX9 port map( A => n6239, Z => n6237);
   U156 : HS65_LH_IVX9 port map( A => n6259, Z => n6258);
   U157 : HS65_LH_IVX9 port map( A => n6259, Z => n6257);
   U158 : HS65_LH_IVX9 port map( A => n6264, Z => n6263);
   U159 : HS65_LH_IVX9 port map( A => n6264, Z => n6262);
   U160 : HS65_LH_IVX9 port map( A => n6209, Z => n6208);
   U161 : HS65_LH_IVX9 port map( A => n6209, Z => n6207);
   U162 : HS65_LH_IVX9 port map( A => n6299, Z => n6298);
   U163 : HS65_LH_IVX9 port map( A => n6299, Z => n6297);
   U164 : HS65_LH_IVX9 port map( A => n6304, Z => n6303);
   U165 : HS65_LH_IVX9 port map( A => n6304, Z => n6302);
   U166 : HS65_LH_IVX9 port map( A => n6229, Z => n6228);
   U167 : HS65_LH_IVX9 port map( A => n6229, Z => n6227);
   U168 : HS65_LH_IVX9 port map( A => n6269, Z => n6268);
   U169 : HS65_LH_IVX9 port map( A => n6269, Z => n6267);
   U170 : HS65_LH_BFX9 port map( A => n1373, Z => n6367);
   U171 : HS65_LH_BFX9 port map( A => n1373, Z => n6368);
   U172 : HS65_LH_BFX9 port map( A => n882, Z => n6460);
   U173 : HS65_LH_BFX9 port map( A => n882, Z => n6461);
   U174 : HS65_LH_IVX9 port map( A => n6324, Z => n6323);
   U175 : HS65_LH_IVX9 port map( A => n6324, Z => n6322);
   U176 : HS65_LH_IVX9 port map( A => n6309, Z => n6308);
   U177 : HS65_LH_IVX9 port map( A => n6309, Z => n6307);
   U178 : HS65_LH_IVX9 port map( A => n6319, Z => n6318);
   U179 : HS65_LH_IVX9 port map( A => n6319, Z => n6317);
   U180 : HS65_LH_IVX9 port map( A => n6314, Z => n6313);
   U181 : HS65_LH_IVX9 port map( A => n6314, Z => n6312);
   U182 : HS65_LH_IVX9 port map( A => n6219, Z => n6218);
   U183 : HS65_LH_IVX9 port map( A => n6219, Z => n6217);
   U184 : HS65_LH_IVX9 port map( A => n6224, Z => n6223);
   U185 : HS65_LH_IVX9 port map( A => n6224, Z => n6222);
   U186 : HS65_LH_IVX9 port map( A => n6249, Z => n6248);
   U187 : HS65_LH_IVX9 port map( A => n6249, Z => n6247);
   U188 : HS65_LH_IVX9 port map( A => n6254, Z => n6253);
   U189 : HS65_LH_IVX9 port map( A => n6254, Z => n6252);
   U190 : HS65_LH_BFX9 port map( A => n6168, Z => n6330);
   U191 : HS65_LH_BFX9 port map( A => n6167, Z => n6335);
   U192 : HS65_LH_BFX9 port map( A => n6171, Z => n6275);
   U193 : HS65_LH_BFX9 port map( A => n6172, Z => n6280);
   U194 : HS65_LH_BFX9 port map( A => n6173, Z => n6285);
   U195 : HS65_LH_BFX9 port map( A => n6175, Z => n6290);
   U196 : HS65_LH_BFX9 port map( A => n6174, Z => n6295);
   U197 : HS65_LH_BFX9 port map( A => n6180, Z => n6185);
   U198 : HS65_LH_BFX9 port map( A => n6181, Z => n6215);
   U199 : HS65_LH_BFX9 port map( A => n6170, Z => n6235);
   U200 : HS65_LH_BFX9 port map( A => n6169, Z => n6245);
   U201 : HS65_LH_BFX9 port map( A => n6178, Z => n6190);
   U202 : HS65_LH_BFX9 port map( A => n6177, Z => n6195);
   U203 : HS65_LH_BFX9 port map( A => n6176, Z => n6200);
   U204 : HS65_LH_BFX9 port map( A => n6179, Z => n6205);
   U205 : HS65_LH_BFX9 port map( A => n1373, Z => n6369);
   U206 : HS65_LH_BFX9 port map( A => n882, Z => n6462);
   U207 : HS65_LH_IVX9 port map( A => n6234, Z => n6232);
   U208 : HS65_LH_IVX9 port map( A => n6234, Z => n6233);
   U209 : HS65_LH_IVX9 port map( A => n6244, Z => n6242);
   U210 : HS65_LH_IVX9 port map( A => n6244, Z => n6243);
   U211 : HS65_LH_IVX9 port map( A => n6189, Z => n6187);
   U212 : HS65_LH_IVX9 port map( A => n6189, Z => n6188);
   U213 : HS65_LH_IVX9 port map( A => n6194, Z => n6192);
   U214 : HS65_LH_IVX9 port map( A => n6194, Z => n6193);
   U215 : HS65_LH_IVX9 port map( A => n6199, Z => n6197);
   U216 : HS65_LH_IVX9 port map( A => n6199, Z => n6198);
   U217 : HS65_LH_IVX9 port map( A => n6204, Z => n6202);
   U218 : HS65_LH_IVX9 port map( A => n6204, Z => n6203);
   U219 : HS65_LH_IVX9 port map( A => n6274, Z => n6272);
   U220 : HS65_LH_IVX9 port map( A => n6274, Z => n6273);
   U221 : HS65_LH_IVX9 port map( A => n6279, Z => n6277);
   U222 : HS65_LH_IVX9 port map( A => n6279, Z => n6278);
   U223 : HS65_LH_IVX9 port map( A => n6284, Z => n6282);
   U224 : HS65_LH_IVX9 port map( A => n6284, Z => n6283);
   U225 : HS65_LH_IVX9 port map( A => n6289, Z => n6287);
   U226 : HS65_LH_IVX9 port map( A => n6289, Z => n6288);
   U227 : HS65_LH_IVX9 port map( A => n6294, Z => n6292);
   U228 : HS65_LH_IVX9 port map( A => n6294, Z => n6293);
   U229 : HS65_LH_IVX9 port map( A => n6184, Z => n6182);
   U230 : HS65_LH_IVX9 port map( A => n6184, Z => n6183);
   U231 : HS65_LH_IVX9 port map( A => n6214, Z => n6212);
   U232 : HS65_LH_IVX9 port map( A => n6214, Z => n6213);
   U233 : HS65_LH_IVX9 port map( A => n6329, Z => n6327);
   U234 : HS65_LH_IVX9 port map( A => n6329, Z => n6328);
   U235 : HS65_LH_IVX9 port map( A => n6334, Z => n6332);
   U236 : HS65_LH_IVX9 port map( A => n6334, Z => n6333);
   U237 : HS65_LH_BFX9 port map( A => n6168, Z => n6331);
   U238 : HS65_LH_BFX9 port map( A => n6167, Z => n6336);
   U239 : HS65_LH_BFX9 port map( A => n6171, Z => n6276);
   U240 : HS65_LH_BFX9 port map( A => n6172, Z => n6281);
   U241 : HS65_LH_BFX9 port map( A => n6173, Z => n6286);
   U242 : HS65_LH_BFX9 port map( A => n6175, Z => n6291);
   U243 : HS65_LH_BFX9 port map( A => n6174, Z => n6296);
   U244 : HS65_LH_BFX9 port map( A => n6180, Z => n6186);
   U245 : HS65_LH_BFX9 port map( A => n6181, Z => n6216);
   U246 : HS65_LH_BFX9 port map( A => n6170, Z => n6236);
   U247 : HS65_LH_BFX9 port map( A => n6169, Z => n6246);
   U248 : HS65_LH_BFX9 port map( A => n6178, Z => n6191);
   U249 : HS65_LH_BFX9 port map( A => n6177, Z => n6196);
   U250 : HS65_LH_BFX9 port map( A => n6176, Z => n6201);
   U251 : HS65_LH_BFX9 port map( A => n6179, Z => n6206);
   U252 : HS65_LH_BFX9 port map( A => n6659, Z => n6642);
   U253 : HS65_LH_BFX9 port map( A => n6659, Z => n6643);
   U254 : HS65_LH_BFX9 port map( A => n6657, Z => n6652);
   U255 : HS65_LH_BFX9 port map( A => n6657, Z => n6653);
   U256 : HS65_LH_BFX9 port map( A => n6659, Z => n6644);
   U257 : HS65_LH_BFX9 port map( A => n6659, Z => n6645);
   U258 : HS65_LH_BFX9 port map( A => n6658, Z => n6648);
   U259 : HS65_LH_BFX9 port map( A => n6659, Z => n6646);
   U260 : HS65_LH_BFX9 port map( A => n6658, Z => n6647);
   U261 : HS65_LH_BFX9 port map( A => n6658, Z => n6649);
   U262 : HS65_LH_BFX9 port map( A => n6658, Z => n6650);
   U263 : HS65_LH_BFX9 port map( A => n6658, Z => n6651);
   U264 : HS65_LH_BFX9 port map( A => n6660, Z => n6637);
   U265 : HS65_LH_BFX9 port map( A => n6660, Z => n6638);
   U266 : HS65_LH_BFX9 port map( A => n6657, Z => n6654);
   U267 : HS65_LH_BFX9 port map( A => n6657, Z => n6656);
   U268 : HS65_LH_BFX9 port map( A => n6662, Z => n6627);
   U269 : HS65_LH_BFX9 port map( A => n6662, Z => n6628);
   U270 : HS65_LH_BFX9 port map( A => n6662, Z => n6629);
   U271 : HS65_LH_BFX9 port map( A => n6662, Z => n6631);
   U272 : HS65_LH_BFX9 port map( A => n6662, Z => n6630);
   U273 : HS65_LH_BFX9 port map( A => n6661, Z => n6634);
   U274 : HS65_LH_BFX9 port map( A => n6661, Z => n6632);
   U275 : HS65_LH_BFX9 port map( A => n6661, Z => n6633);
   U276 : HS65_LH_BFX9 port map( A => n6661, Z => n6635);
   U277 : HS65_LH_BFX9 port map( A => n6661, Z => n6636);
   U278 : HS65_LH_BFX9 port map( A => n6660, Z => n6641);
   U279 : HS65_LH_BFX9 port map( A => n6660, Z => n6639);
   U280 : HS65_LH_BFX9 port map( A => n6660, Z => n6640);
   U281 : HS65_LH_BFX9 port map( A => n6657, Z => n6655);
   U282 : HS65_LH_BFX9 port map( A => n6663, Z => n6625);
   U283 : HS65_LH_BFX9 port map( A => n6663, Z => n6624);
   U284 : HS65_LH_BFX9 port map( A => n6663, Z => n6623);
   U285 : HS65_LH_BFX9 port map( A => n6663, Z => n6622);
   U286 : HS65_LH_BFX9 port map( A => n6664, Z => n6621);
   U287 : HS65_LH_BFX9 port map( A => n6664, Z => n6620);
   U288 : HS65_LH_BFX9 port map( A => n6664, Z => n6619);
   U289 : HS65_LH_BFX9 port map( A => n6664, Z => n6618);
   U290 : HS65_LH_BFX9 port map( A => n6664, Z => n6617);
   U291 : HS65_LH_BFX9 port map( A => n6663, Z => n6626);
   U292 : HS65_LH_BFX9 port map( A => n2853, Z => n6239);
   U293 : HS65_LH_BFX9 port map( A => n2848, Z => n6259);
   U294 : HS65_LH_BFX9 port map( A => n2847, Z => n6264);
   U295 : HS65_LH_BFX9 port map( A => n2860, Z => n6209);
   U296 : HS65_LH_BFX9 port map( A => n2857, Z => n6219);
   U297 : HS65_LH_BFX9 port map( A => n2856, Z => n6224);
   U298 : HS65_LH_BFX9 port map( A => n2851, Z => n6249);
   U299 : HS65_LH_BFX9 port map( A => n2849, Z => n6254);
   U300 : HS65_LH_BFX9 port map( A => n2855, Z => n6229);
   U301 : HS65_LH_BFX9 port map( A => n2846, Z => n6269);
   U302 : HS65_LH_BFX9 port map( A => n2828, Z => n6324);
   U303 : HS65_LH_BFX9 port map( A => n2834, Z => n6309);
   U304 : HS65_LH_BFX9 port map( A => n2830, Z => n6319);
   U305 : HS65_LH_BFX9 port map( A => n2832, Z => n6314);
   U306 : HS65_LH_BFX9 port map( A => n2838, Z => n6299);
   U307 : HS65_LH_BFX9 port map( A => n2836, Z => n6304);
   U308 : HS65_LH_BFX9 port map( A => n2857, Z => n6220);
   U309 : HS65_LH_BFX9 port map( A => n2856, Z => n6225);
   U310 : HS65_LH_BFX9 port map( A => n2851, Z => n6250);
   U311 : HS65_LH_BFX9 port map( A => n2849, Z => n6255);
   U312 : HS65_LH_BFX9 port map( A => n2855, Z => n6230);
   U313 : HS65_LH_BFX9 port map( A => n2846, Z => n6270);
   U314 : HS65_LH_BFX9 port map( A => n2828, Z => n6325);
   U315 : HS65_LH_BFX9 port map( A => n2834, Z => n6310);
   U316 : HS65_LH_BFX9 port map( A => n2830, Z => n6320);
   U317 : HS65_LH_BFX9 port map( A => n2832, Z => n6315);
   U318 : HS65_LH_BFX9 port map( A => n2838, Z => n6300);
   U319 : HS65_LH_BFX9 port map( A => n2836, Z => n6305);
   U320 : HS65_LH_BFX9 port map( A => n2853, Z => n6240);
   U321 : HS65_LH_BFX9 port map( A => n2848, Z => n6260);
   U322 : HS65_LH_BFX9 port map( A => n2847, Z => n6265);
   U323 : HS65_LH_BFX9 port map( A => n2860, Z => n6210);
   U324 : HS65_LH_BFX9 port map( A => n1352, Z => n6415);
   U325 : HS65_LH_BFX9 port map( A => n1352, Z => n6416);
   U326 : HS65_LH_BFX9 port map( A => n861, Z => n6508);
   U327 : HS65_LH_BFX9 port map( A => n861, Z => n6509);
   U328 : HS65_LH_BFX9 port map( A => n6168, Z => n6329);
   U329 : HS65_LH_BFX9 port map( A => n6167, Z => n6334);
   U330 : HS65_LH_BFX9 port map( A => n6171, Z => n6274);
   U331 : HS65_LH_BFX9 port map( A => n6172, Z => n6279);
   U332 : HS65_LH_BFX9 port map( A => n6173, Z => n6284);
   U333 : HS65_LH_BFX9 port map( A => n6175, Z => n6289);
   U334 : HS65_LH_BFX9 port map( A => n6174, Z => n6294);
   U335 : HS65_LH_BFX9 port map( A => n6180, Z => n6184);
   U336 : HS65_LH_BFX9 port map( A => n6181, Z => n6214);
   U337 : HS65_LH_BFX9 port map( A => n6170, Z => n6234);
   U338 : HS65_LH_BFX9 port map( A => n6169, Z => n6244);
   U339 : HS65_LH_BFX9 port map( A => n6178, Z => n6189);
   U340 : HS65_LH_BFX9 port map( A => n6177, Z => n6194);
   U341 : HS65_LH_BFX9 port map( A => n6176, Z => n6199);
   U342 : HS65_LH_BFX9 port map( A => n6179, Z => n6204);
   U343 : HS65_LH_BFX9 port map( A => n1353, Z => n6412);
   U344 : HS65_LH_BFX9 port map( A => n1353, Z => n6413);
   U345 : HS65_LH_BFX9 port map( A => n1354, Z => n6409);
   U346 : HS65_LH_BFX9 port map( A => n1354, Z => n6410);
   U347 : HS65_LH_BFX9 port map( A => n862, Z => n6505);
   U348 : HS65_LH_BFX9 port map( A => n862, Z => n6506);
   U349 : HS65_LH_BFX9 port map( A => n863, Z => n6502);
   U350 : HS65_LH_BFX9 port map( A => n863, Z => n6503);
   U351 : HS65_LH_BFX9 port map( A => n881, Z => n6463);
   U352 : HS65_LH_BFX9 port map( A => n856, Z => n6520);
   U353 : HS65_LH_BFX9 port map( A => n881, Z => n6464);
   U354 : HS65_LH_BFX9 port map( A => n856, Z => n6521);
   U355 : HS65_LH_BFX9 port map( A => n1372, Z => n6370);
   U356 : HS65_LH_BFX9 port map( A => n1367, Z => n6382);
   U357 : HS65_LH_BFX9 port map( A => n1347, Z => n6427);
   U358 : HS65_LH_BFX9 port map( A => n1372, Z => n6371);
   U359 : HS65_LH_BFX9 port map( A => n1367, Z => n6383);
   U360 : HS65_LH_BFX9 port map( A => n1347, Z => n6428);
   U361 : HS65_LH_BFX9 port map( A => n885, Z => n6454);
   U362 : HS65_LH_BFX9 port map( A => n885, Z => n6455);
   U363 : HS65_LH_BFX9 port map( A => n860, Z => n6511);
   U364 : HS65_LH_BFX9 port map( A => n860, Z => n6512);
   U365 : HS65_LH_BFX9 port map( A => n880, Z => n6466);
   U366 : HS65_LH_BFX9 port map( A => n880, Z => n6467);
   U367 : HS65_LH_BFX9 port map( A => n1348, Z => n6424);
   U368 : HS65_LH_BFX9 port map( A => n1348, Z => n6425);
   U369 : HS65_LH_BFX9 port map( A => n1368, Z => n6379);
   U370 : HS65_LH_BFX9 port map( A => n1368, Z => n6380);
   U371 : HS65_LH_BFX9 port map( A => n876, Z => n6475);
   U372 : HS65_LH_BFX9 port map( A => n876, Z => n6476);
   U373 : HS65_LH_BFX9 port map( A => n879, Z => n6469);
   U374 : HS65_LH_BFX9 port map( A => n879, Z => n6470);
   U375 : HS65_LH_BFX9 port map( A => n1371, Z => n6373);
   U376 : HS65_LH_BFX9 port map( A => n1371, Z => n6374);
   U377 : HS65_LH_BFX9 port map( A => n877, Z => n6472);
   U378 : HS65_LH_BFX9 port map( A => n857, Z => n6517);
   U379 : HS65_LH_BFX9 port map( A => n877, Z => n6473);
   U380 : HS65_LH_BFX9 port map( A => n857, Z => n6518);
   U381 : HS65_LH_BFX9 port map( A => n1376, Z => n6361);
   U382 : HS65_LH_BFX9 port map( A => n1351, Z => n6418);
   U383 : HS65_LH_BFX9 port map( A => n1376, Z => n6362);
   U384 : HS65_LH_BFX9 port map( A => n1351, Z => n6419);
   U385 : HS65_LH_BFX9 port map( A => n859, Z => n6514);
   U386 : HS65_LH_BFX9 port map( A => n859, Z => n6515);
   U387 : HS65_LH_BFX9 port map( A => n884, Z => n6457);
   U388 : HS65_LH_BFX9 port map( A => n884, Z => n6458);
   U389 : HS65_LH_BFX9 port map( A => n2853, Z => n6241);
   U390 : HS65_LH_BFX9 port map( A => n2848, Z => n6261);
   U391 : HS65_LH_BFX9 port map( A => n2847, Z => n6266);
   U392 : HS65_LH_BFX9 port map( A => n1352, Z => n6417);
   U393 : HS65_LH_BFX9 port map( A => n861, Z => n6510);
   U394 : HS65_LH_BFX9 port map( A => n2860, Z => n6211);
   U395 : HS65_LH_BFX9 port map( A => n1375, Z => n6364);
   U396 : HS65_LH_BFX9 port map( A => n1370, Z => n6376);
   U397 : HS65_LH_BFX9 port map( A => n1350, Z => n6421);
   U398 : HS65_LH_BFX9 port map( A => n1375, Z => n6365);
   U399 : HS65_LH_BFX9 port map( A => n1370, Z => n6377);
   U400 : HS65_LH_BFX9 port map( A => n1350, Z => n6422);
   U401 : HS65_LH_BFX9 port map( A => n1353, Z => n6414);
   U402 : HS65_LH_BFX9 port map( A => n862, Z => n6507);
   U403 : HS65_LH_BFX9 port map( A => n2857, Z => n6221);
   U404 : HS65_LH_BFX9 port map( A => n2856, Z => n6226);
   U405 : HS65_LH_BFX9 port map( A => n2851, Z => n6251);
   U406 : HS65_LH_BFX9 port map( A => n2849, Z => n6256);
   U407 : HS65_LH_BFX9 port map( A => n2855, Z => n6231);
   U408 : HS65_LH_BFX9 port map( A => n2846, Z => n6271);
   U409 : HS65_LH_BFX9 port map( A => n2828, Z => n6326);
   U410 : HS65_LH_BFX9 port map( A => n2834, Z => n6311);
   U411 : HS65_LH_BFX9 port map( A => n2830, Z => n6321);
   U412 : HS65_LH_BFX9 port map( A => n2832, Z => n6316);
   U413 : HS65_LH_BFX9 port map( A => n2838, Z => n6301);
   U414 : HS65_LH_BFX9 port map( A => n2836, Z => n6306);
   U415 : HS65_LH_BFX9 port map( A => n863, Z => n6504);
   U416 : HS65_LH_BFX9 port map( A => n888, Z => n6445);
   U417 : HS65_LH_BFX9 port map( A => n866, Z => n6493);
   U418 : HS65_LH_BFX9 port map( A => n888, Z => n6446);
   U419 : HS65_LH_BFX9 port map( A => n866, Z => n6494);
   U420 : HS65_LH_BFX9 port map( A => n1379, Z => n6352);
   U421 : HS65_LH_BFX9 port map( A => n1383, Z => n6340);
   U422 : HS65_LH_BFX9 port map( A => n1361, Z => n6388);
   U423 : HS65_LH_BFX9 port map( A => n1357, Z => n6400);
   U424 : HS65_LH_BFX9 port map( A => n1379, Z => n6353);
   U425 : HS65_LH_BFX9 port map( A => n1383, Z => n6341);
   U426 : HS65_LH_BFX9 port map( A => n1361, Z => n6389);
   U427 : HS65_LH_BFX9 port map( A => n1357, Z => n6401);
   U428 : HS65_LH_BFX9 port map( A => n886, Z => n6451);
   U429 : HS65_LH_BFX9 port map( A => n886, Z => n6452);
   U430 : HS65_LH_BFX9 port map( A => n1381, Z => n6346);
   U431 : HS65_LH_BFX9 port map( A => n1381, Z => n6347);
   U432 : HS65_LH_BFX9 port map( A => n1377, Z => n6358);
   U433 : HS65_LH_BFX9 port map( A => n1359, Z => n6394);
   U434 : HS65_LH_BFX9 port map( A => n1355, Z => n6406);
   U435 : HS65_LH_BFX9 port map( A => n1377, Z => n6359);
   U436 : HS65_LH_BFX9 port map( A => n1359, Z => n6395);
   U437 : HS65_LH_BFX9 port map( A => n1355, Z => n6407);
   U438 : HS65_LH_BFX9 port map( A => n865, Z => n6496);
   U439 : HS65_LH_BFX9 port map( A => n865, Z => n6497);
   U440 : HS65_LH_BFX9 port map( A => n1378, Z => n6355);
   U441 : HS65_LH_BFX9 port map( A => n1382, Z => n6343);
   U442 : HS65_LH_BFX9 port map( A => n1360, Z => n6391);
   U443 : HS65_LH_BFX9 port map( A => n1356, Z => n6403);
   U444 : HS65_LH_BFX9 port map( A => n1378, Z => n6356);
   U445 : HS65_LH_BFX9 port map( A => n1382, Z => n6344);
   U446 : HS65_LH_BFX9 port map( A => n1360, Z => n6392);
   U447 : HS65_LH_BFX9 port map( A => n1356, Z => n6404);
   U448 : HS65_LH_BFX9 port map( A => n893, Z => n6430);
   U449 : HS65_LH_BFX9 port map( A => n893, Z => n6431);
   U450 : HS65_LH_BFX9 port map( A => n1380, Z => n6349);
   U451 : HS65_LH_BFX9 port map( A => n1384, Z => n6337);
   U452 : HS65_LH_BFX9 port map( A => n1362, Z => n6385);
   U453 : HS65_LH_BFX9 port map( A => n1358, Z => n6397);
   U454 : HS65_LH_BFX9 port map( A => n1380, Z => n6350);
   U455 : HS65_LH_BFX9 port map( A => n1384, Z => n6338);
   U456 : HS65_LH_BFX9 port map( A => n1362, Z => n6386);
   U457 : HS65_LH_BFX9 port map( A => n1358, Z => n6398);
   U458 : HS65_LH_BFX9 port map( A => n876, Z => n6477);
   U459 : HS65_LH_BFX9 port map( A => n889, Z => n6442);
   U460 : HS65_LH_BFX9 port map( A => n871, Z => n6478);
   U461 : HS65_LH_BFX9 port map( A => n867, Z => n6490);
   U462 : HS65_LH_BFX9 port map( A => n889, Z => n6443);
   U463 : HS65_LH_BFX9 port map( A => n871, Z => n6479);
   U464 : HS65_LH_BFX9 port map( A => n867, Z => n6491);
   U465 : HS65_LH_BFX9 port map( A => n887, Z => n6448);
   U466 : HS65_LH_BFX9 port map( A => n891, Z => n6436);
   U467 : HS65_LH_BFX9 port map( A => n869, Z => n6484);
   U468 : HS65_LH_BFX9 port map( A => n887, Z => n6449);
   U469 : HS65_LH_BFX9 port map( A => n891, Z => n6437);
   U470 : HS65_LH_BFX9 port map( A => n869, Z => n6485);
   U471 : HS65_LH_BFX9 port map( A => n879, Z => n6471);
   U472 : HS65_LH_BFX9 port map( A => n884, Z => n6459);
   U473 : HS65_LH_BFX9 port map( A => n859, Z => n6516);
   U474 : HS65_LH_BFX9 port map( A => n890, Z => n6439);
   U475 : HS65_LH_BFX9 port map( A => n868, Z => n6487);
   U476 : HS65_LH_BFX9 port map( A => n864, Z => n6499);
   U477 : HS65_LH_BFX9 port map( A => n890, Z => n6440);
   U478 : HS65_LH_BFX9 port map( A => n868, Z => n6488);
   U479 : HS65_LH_BFX9 port map( A => n864, Z => n6500);
   U480 : HS65_LH_BFX9 port map( A => n1354, Z => n6411);
   U481 : HS65_LH_BFX9 port map( A => n892, Z => n6433);
   U482 : HS65_LH_BFX9 port map( A => n870, Z => n6481);
   U483 : HS65_LH_BFX9 port map( A => n892, Z => n6434);
   U484 : HS65_LH_BFX9 port map( A => n870, Z => n6482);
   U485 : HS65_LH_BFX9 port map( A => n1375, Z => n6366);
   U486 : HS65_LH_BFX9 port map( A => n1370, Z => n6378);
   U487 : HS65_LH_BFX9 port map( A => n1350, Z => n6423);
   U488 : HS65_LH_BFX9 port map( A => n881, Z => n6465);
   U489 : HS65_LH_BFX9 port map( A => n856, Z => n6522);
   U490 : HS65_LH_BFX9 port map( A => n1372, Z => n6372);
   U491 : HS65_LH_BFX9 port map( A => n1367, Z => n6384);
   U492 : HS65_LH_BFX9 port map( A => n1347, Z => n6429);
   U493 : HS65_LH_BFX9 port map( A => n885, Z => n6456);
   U494 : HS65_LH_BFX9 port map( A => n860, Z => n6513);
   U495 : HS65_LH_BFX9 port map( A => n880, Z => n6468);
   U496 : HS65_LH_BFX9 port map( A => n1371, Z => n6375);
   U497 : HS65_LH_BFX9 port map( A => n1351, Z => n6420);
   U498 : HS65_LH_BFX9 port map( A => n1376, Z => n6363);
   U499 : HS65_LH_BFX9 port map( A => n1348, Z => n6426);
   U500 : HS65_LH_BFX9 port map( A => n1368, Z => n6381);
   U501 : HS65_LH_BFX9 port map( A => n877, Z => n6474);
   U502 : HS65_LH_BFX9 port map( A => n857, Z => n6519);
   U503 : HS65_LH_BFX9 port map( A => n865, Z => n6498);
   U504 : HS65_LH_BFX9 port map( A => n1378, Z => n6357);
   U505 : HS65_LH_BFX9 port map( A => n1382, Z => n6345);
   U506 : HS65_LH_BFX9 port map( A => n1360, Z => n6393);
   U507 : HS65_LH_BFX9 port map( A => n1356, Z => n6405);
   U508 : HS65_LH_BFX9 port map( A => n893, Z => n6432);
   U509 : HS65_LH_BFX9 port map( A => n1380, Z => n6351);
   U510 : HS65_LH_BFX9 port map( A => n1384, Z => n6339);
   U511 : HS65_LH_BFX9 port map( A => n1362, Z => n6387);
   U512 : HS65_LH_BFX9 port map( A => n1358, Z => n6399);
   U513 : HS65_LH_BFX9 port map( A => n889, Z => n6444);
   U514 : HS65_LH_BFX9 port map( A => n871, Z => n6480);
   U515 : HS65_LH_BFX9 port map( A => n867, Z => n6492);
   U516 : HS65_LH_BFX9 port map( A => n887, Z => n6450);
   U517 : HS65_LH_BFX9 port map( A => n891, Z => n6438);
   U518 : HS65_LH_BFX9 port map( A => n869, Z => n6486);
   U519 : HS65_LH_BFX9 port map( A => n890, Z => n6441);
   U520 : HS65_LH_BFX9 port map( A => n868, Z => n6489);
   U521 : HS65_LH_BFX9 port map( A => n864, Z => n6501);
   U522 : HS65_LH_BFX9 port map( A => n892, Z => n6435);
   U523 : HS65_LH_BFX9 port map( A => n870, Z => n6483);
   U524 : HS65_LH_BFX9 port map( A => n888, Z => n6447);
   U525 : HS65_LH_BFX9 port map( A => n866, Z => n6495);
   U526 : HS65_LH_BFX9 port map( A => n1379, Z => n6354);
   U527 : HS65_LH_BFX9 port map( A => n1383, Z => n6342);
   U528 : HS65_LH_BFX9 port map( A => n1361, Z => n6390);
   U529 : HS65_LH_BFX9 port map( A => n1357, Z => n6402);
   U530 : HS65_LH_BFX9 port map( A => n886, Z => n6453);
   U531 : HS65_LH_BFX9 port map( A => n1381, Z => n6348);
   U532 : HS65_LH_BFX9 port map( A => n1377, Z => n6360);
   U533 : HS65_LH_BFX9 port map( A => n1359, Z => n6396);
   U534 : HS65_LH_BFX9 port map( A => n1355, Z => n6408);
   U535 : HS65_LH_BFX9 port map( A => n6533, Z => n6659);
   U536 : HS65_LH_BFX9 port map( A => n6533, Z => n6658);
   U537 : HS65_LH_BFX9 port map( A => n6534, Z => n6662);
   U538 : HS65_LH_BFX9 port map( A => n6534, Z => n6661);
   U539 : HS65_LH_BFX9 port map( A => n6534, Z => n6660);
   U540 : HS65_LH_BFX9 port map( A => n6533, Z => n6657);
   U541 : HS65_LH_BFX9 port map( A => n6535, Z => n6664);
   U542 : HS65_LH_BFX9 port map( A => n6535, Z => n6663);
   U543 : HS65_LH_OAI22X6 port map( A => n6303, B => n288, C => n846, D => 
                           n6304, Z => n2202);
   U544 : HS65_LH_OAI22X6 port map( A => n6302, B => n287, C => n845, D => 
                           n6305, Z => n2203);
   U545 : HS65_LH_OAI22X6 port map( A => n6303, B => n286, C => n844, D => 
                           n6305, Z => n2204);
   U546 : HS65_LH_OAI22X6 port map( A => n6302, B => n285, C => n843, D => 
                           n6305, Z => n2205);
   U547 : HS65_LH_OAI22X6 port map( A => n6303, B => n284, C => n842, D => 
                           n6305, Z => n2206);
   U548 : HS65_LH_OAI22X6 port map( A => n6302, B => n283, C => n841, D => 
                           n6305, Z => n2207);
   U549 : HS65_LH_OAI22X6 port map( A => n6303, B => n282, C => n840, D => 
                           n6305, Z => n2208);
   U550 : HS65_LH_OAI22X6 port map( A => n6302, B => n281, C => n839, D => 
                           n6305, Z => n2209);
   U551 : HS65_LH_OAI22X6 port map( A => n6303, B => n280, C => n838, D => 
                           n6305, Z => n2210);
   U552 : HS65_LH_OAI22X6 port map( A => n6303, B => n279, C => n837, D => 
                           n6305, Z => n2211);
   U553 : HS65_LH_OAI22X6 port map( A => n6303, B => n278, C => n836, D => 
                           n6305, Z => n2212);
   U554 : HS65_LH_OAI22X6 port map( A => n6303, B => n277, C => n835, D => 
                           n6305, Z => n2213);
   U555 : HS65_LH_OAI22X6 port map( A => n6303, B => n276, C => n834, D => 
                           n6305, Z => n2214);
   U556 : HS65_LH_OAI22X6 port map( A => n6303, B => n275, C => n833, D => 
                           n6305, Z => n2215);
   U557 : HS65_LH_OAI22X6 port map( A => n6303, B => n274, C => n832, D => 
                           n6305, Z => n2216);
   U558 : HS65_LH_OAI22X6 port map( A => n6303, B => n273, C => n831, D => 
                           n6305, Z => n2217);
   U559 : HS65_LH_OAI22X6 port map( A => n6303, B => n272, C => n830, D => 
                           n6305, Z => n2218);
   U560 : HS65_LH_OAI22X6 port map( A => n6303, B => n271, C => n829, D => 
                           n6305, Z => n2219);
   U561 : HS65_LH_OAI22X6 port map( A => n6303, B => n270, C => n828, D => 
                           n6305, Z => n2220);
   U562 : HS65_LH_OAI22X6 port map( A => n6303, B => n269, C => n827, D => 
                           n6305, Z => n2221);
   U563 : HS65_LH_OAI22X6 port map( A => n6302, B => n268, C => n826, D => 
                           n6306, Z => n2222);
   U564 : HS65_LH_OAI22X6 port map( A => n6302, B => n267, C => n825, D => 
                           n6306, Z => n2223);
   U565 : HS65_LH_OAI22X6 port map( A => n6302, B => n266, C => n824, D => 
                           n6306, Z => n2224);
   U566 : HS65_LH_OAI22X6 port map( A => n6302, B => n265, C => n823, D => 
                           n6306, Z => n2225);
   U567 : HS65_LH_OAI22X6 port map( A => n6302, B => n264, C => n822, D => 
                           n6306, Z => n2226);
   U568 : HS65_LH_OAI22X6 port map( A => n6302, B => n263, C => n821, D => 
                           n6306, Z => n2227);
   U569 : HS65_LH_OAI22X6 port map( A => n6302, B => n262, C => n820, D => 
                           n6306, Z => n2228);
   U570 : HS65_LH_OAI22X6 port map( A => n6302, B => n261, C => n819, D => 
                           n6306, Z => n2229);
   U571 : HS65_LH_OAI22X6 port map( A => n6302, B => n260, C => n818, D => 
                           n6306, Z => n2230);
   U572 : HS65_LH_OAI22X6 port map( A => n6302, B => n259, C => n817, D => 
                           n6306, Z => n2231);
   U573 : HS65_LH_OAI22X6 port map( A => n6302, B => n258, C => n816, D => 
                           n6306, Z => n2232);
   U574 : HS65_LH_OAI22X6 port map( A => n6302, B => n257, C => n815, D => 
                           n6306, Z => n2233);
   U575 : HS65_LH_OAI22X6 port map( A => n6228, B => n480, C => n846, D => 
                           n6229, Z => n1722);
   U576 : HS65_LH_OAI22X6 port map( A => n6227, B => n479, C => n845, D => 
                           n6230, Z => n1723);
   U577 : HS65_LH_OAI22X6 port map( A => n6228, B => n478, C => n844, D => 
                           n6230, Z => n1724);
   U578 : HS65_LH_OAI22X6 port map( A => n6227, B => n477, C => n843, D => 
                           n6230, Z => n1725);
   U579 : HS65_LH_OAI22X6 port map( A => n6228, B => n476, C => n842, D => 
                           n6230, Z => n1726);
   U580 : HS65_LH_OAI22X6 port map( A => n6227, B => n475, C => n841, D => 
                           n6230, Z => n1727);
   U581 : HS65_LH_OAI22X6 port map( A => n6228, B => n474, C => n840, D => 
                           n6230, Z => n1728);
   U582 : HS65_LH_OAI22X6 port map( A => n6227, B => n473, C => n839, D => 
                           n6230, Z => n1729);
   U583 : HS65_LH_OAI22X6 port map( A => n6228, B => n472, C => n838, D => 
                           n6230, Z => n1730);
   U584 : HS65_LH_OAI22X6 port map( A => n6228, B => n471, C => n837, D => 
                           n6230, Z => n1731);
   U585 : HS65_LH_OAI22X6 port map( A => n6228, B => n470, C => n836, D => 
                           n6230, Z => n1732);
   U586 : HS65_LH_OAI22X6 port map( A => n6228, B => n469, C => n835, D => 
                           n6230, Z => n1733);
   U587 : HS65_LH_OAI22X6 port map( A => n6228, B => n468, C => n834, D => 
                           n6230, Z => n1734);
   U588 : HS65_LH_OAI22X6 port map( A => n6228, B => n467, C => n833, D => 
                           n6230, Z => n1735);
   U589 : HS65_LH_OAI22X6 port map( A => n6228, B => n466, C => n832, D => 
                           n6230, Z => n1736);
   U590 : HS65_LH_OAI22X6 port map( A => n6228, B => n465, C => n831, D => 
                           n6230, Z => n1737);
   U591 : HS65_LH_OAI22X6 port map( A => n6228, B => n464, C => n830, D => 
                           n6230, Z => n1738);
   U592 : HS65_LH_OAI22X6 port map( A => n6228, B => n463, C => n829, D => 
                           n6230, Z => n1739);
   U593 : HS65_LH_OAI22X6 port map( A => n6228, B => n462, C => n828, D => 
                           n6230, Z => n1740);
   U594 : HS65_LH_OAI22X6 port map( A => n6228, B => n461, C => n827, D => 
                           n6230, Z => n1741);
   U595 : HS65_LH_OAI22X6 port map( A => n6227, B => n460, C => n826, D => 
                           n6231, Z => n1742);
   U596 : HS65_LH_OAI22X6 port map( A => n6227, B => n459, C => n825, D => 
                           n6231, Z => n1743);
   U597 : HS65_LH_OAI22X6 port map( A => n6227, B => n458, C => n824, D => 
                           n6231, Z => n1744);
   U598 : HS65_LH_OAI22X6 port map( A => n6227, B => n457, C => n823, D => 
                           n6231, Z => n1745);
   U599 : HS65_LH_OAI22X6 port map( A => n6227, B => n456, C => n822, D => 
                           n6231, Z => n1746);
   U600 : HS65_LH_OAI22X6 port map( A => n6227, B => n455, C => n821, D => 
                           n6231, Z => n1747);
   U601 : HS65_LH_OAI22X6 port map( A => n6227, B => n454, C => n820, D => 
                           n6231, Z => n1748);
   U602 : HS65_LH_OAI22X6 port map( A => n6227, B => n453, C => n819, D => 
                           n6231, Z => n1749);
   U603 : HS65_LH_OAI22X6 port map( A => n6227, B => n452, C => n818, D => 
                           n6231, Z => n1750);
   U604 : HS65_LH_OAI22X6 port map( A => n6227, B => n451, C => n817, D => 
                           n6231, Z => n1751);
   U605 : HS65_LH_OAI22X6 port map( A => n6227, B => n450, C => n816, D => 
                           n6231, Z => n1752);
   U606 : HS65_LH_OAI22X6 port map( A => n6227, B => n449, C => n815, D => 
                           n6231, Z => n1753);
   U607 : HS65_LH_OAI22X6 port map( A => n6268, B => n352, C => n846, D => 
                           n6269, Z => n1978);
   U608 : HS65_LH_OAI22X6 port map( A => n6267, B => n351, C => n845, D => 
                           n6270, Z => n1979);
   U609 : HS65_LH_OAI22X6 port map( A => n6268, B => n350, C => n844, D => 
                           n6270, Z => n1980);
   U610 : HS65_LH_OAI22X6 port map( A => n6267, B => n349, C => n843, D => 
                           n6270, Z => n1981);
   U611 : HS65_LH_OAI22X6 port map( A => n6268, B => n348, C => n842, D => 
                           n6270, Z => n1982);
   U612 : HS65_LH_OAI22X6 port map( A => n6267, B => n347, C => n841, D => 
                           n6270, Z => n1983);
   U613 : HS65_LH_OAI22X6 port map( A => n6268, B => n346, C => n840, D => 
                           n6270, Z => n1984);
   U614 : HS65_LH_OAI22X6 port map( A => n6267, B => n345, C => n839, D => 
                           n6270, Z => n1985);
   U615 : HS65_LH_OAI22X6 port map( A => n6268, B => n344, C => n838, D => 
                           n6270, Z => n1986);
   U616 : HS65_LH_OAI22X6 port map( A => n6268, B => n343, C => n837, D => 
                           n6270, Z => n1987);
   U617 : HS65_LH_OAI22X6 port map( A => n6268, B => n342, C => n836, D => 
                           n6270, Z => n1988);
   U618 : HS65_LH_OAI22X6 port map( A => n6268, B => n341, C => n835, D => 
                           n6270, Z => n1989);
   U619 : HS65_LH_OAI22X6 port map( A => n6268, B => n340, C => n834, D => 
                           n6270, Z => n1990);
   U620 : HS65_LH_OAI22X6 port map( A => n6268, B => n339, C => n833, D => 
                           n6270, Z => n1991);
   U621 : HS65_LH_OAI22X6 port map( A => n6268, B => n338, C => n832, D => 
                           n6270, Z => n1992);
   U622 : HS65_LH_OAI22X6 port map( A => n6268, B => n337, C => n831, D => 
                           n6270, Z => n1993);
   U623 : HS65_LH_OAI22X6 port map( A => n6268, B => n336, C => n830, D => 
                           n6270, Z => n1994);
   U624 : HS65_LH_OAI22X6 port map( A => n6268, B => n335, C => n829, D => 
                           n6270, Z => n1995);
   U625 : HS65_LH_OAI22X6 port map( A => n6268, B => n334, C => n828, D => 
                           n6270, Z => n1996);
   U626 : HS65_LH_OAI22X6 port map( A => n6268, B => n333, C => n827, D => 
                           n6270, Z => n1997);
   U627 : HS65_LH_OAI22X6 port map( A => n6267, B => n332, C => n826, D => 
                           n6271, Z => n1998);
   U628 : HS65_LH_OAI22X6 port map( A => n6267, B => n331, C => n825, D => 
                           n6271, Z => n1999);
   U629 : HS65_LH_OAI22X6 port map( A => n6267, B => n330, C => n824, D => 
                           n6271, Z => n2000);
   U630 : HS65_LH_OAI22X6 port map( A => n6267, B => n329, C => n823, D => 
                           n6271, Z => n2001);
   U631 : HS65_LH_OAI22X6 port map( A => n6267, B => n328, C => n822, D => 
                           n6271, Z => n2002);
   U632 : HS65_LH_OAI22X6 port map( A => n6267, B => n327, C => n821, D => 
                           n6271, Z => n2003);
   U633 : HS65_LH_OAI22X6 port map( A => n6267, B => n326, C => n820, D => 
                           n6271, Z => n2004);
   U634 : HS65_LH_OAI22X6 port map( A => n6267, B => n325, C => n819, D => 
                           n6271, Z => n2005);
   U635 : HS65_LH_OAI22X6 port map( A => n6267, B => n324, C => n818, D => 
                           n6271, Z => n2006);
   U636 : HS65_LH_OAI22X6 port map( A => n6267, B => n323, C => n817, D => 
                           n6271, Z => n2007);
   U637 : HS65_LH_OAI22X6 port map( A => n6267, B => n322, C => n816, D => 
                           n6271, Z => n2008);
   U638 : HS65_LH_OAI22X6 port map( A => n6267, B => n321, C => n815, D => 
                           n6271, Z => n2009);
   U639 : HS65_LH_OAI22X6 port map( A => n6298, B => n320, C => n846, D => 
                           n6299, Z => n2170);
   U640 : HS65_LH_OAI22X6 port map( A => n6297, B => n319, C => n845, D => 
                           n6300, Z => n2171);
   U641 : HS65_LH_OAI22X6 port map( A => n6298, B => n318, C => n844, D => 
                           n6300, Z => n2172);
   U642 : HS65_LH_OAI22X6 port map( A => n6297, B => n317, C => n843, D => 
                           n6300, Z => n2173);
   U643 : HS65_LH_OAI22X6 port map( A => n6298, B => n316, C => n842, D => 
                           n6300, Z => n2174);
   U644 : HS65_LH_OAI22X6 port map( A => n6297, B => n315, C => n841, D => 
                           n6300, Z => n2175);
   U645 : HS65_LH_OAI22X6 port map( A => n6298, B => n314, C => n840, D => 
                           n6300, Z => n2176);
   U646 : HS65_LH_OAI22X6 port map( A => n6297, B => n313, C => n839, D => 
                           n6300, Z => n2177);
   U647 : HS65_LH_OAI22X6 port map( A => n6298, B => n312, C => n838, D => 
                           n6300, Z => n2178);
   U648 : HS65_LH_OAI22X6 port map( A => n6298, B => n311, C => n837, D => 
                           n6300, Z => n2179);
   U649 : HS65_LH_OAI22X6 port map( A => n6298, B => n310, C => n836, D => 
                           n6300, Z => n2180);
   U650 : HS65_LH_OAI22X6 port map( A => n6298, B => n309, C => n835, D => 
                           n6300, Z => n2181);
   U651 : HS65_LH_OAI22X6 port map( A => n6298, B => n308, C => n834, D => 
                           n6300, Z => n2182);
   U652 : HS65_LH_OAI22X6 port map( A => n6298, B => n307, C => n833, D => 
                           n6300, Z => n2183);
   U653 : HS65_LH_OAI22X6 port map( A => n6298, B => n306, C => n832, D => 
                           n6300, Z => n2184);
   U654 : HS65_LH_OAI22X6 port map( A => n6298, B => n305, C => n831, D => 
                           n6300, Z => n2185);
   U655 : HS65_LH_OAI22X6 port map( A => n6298, B => n304, C => n830, D => 
                           n6300, Z => n2186);
   U656 : HS65_LH_OAI22X6 port map( A => n6298, B => n303, C => n829, D => 
                           n6300, Z => n2187);
   U657 : HS65_LH_OAI22X6 port map( A => n6298, B => n302, C => n828, D => 
                           n6300, Z => n2188);
   U658 : HS65_LH_OAI22X6 port map( A => n6298, B => n301, C => n827, D => 
                           n6300, Z => n2189);
   U659 : HS65_LH_OAI22X6 port map( A => n6297, B => n300, C => n826, D => 
                           n6301, Z => n2190);
   U660 : HS65_LH_OAI22X6 port map( A => n6297, B => n299, C => n825, D => 
                           n6301, Z => n2191);
   U661 : HS65_LH_OAI22X6 port map( A => n6297, B => n298, C => n824, D => 
                           n6301, Z => n2192);
   U662 : HS65_LH_OAI22X6 port map( A => n6297, B => n297, C => n823, D => 
                           n6301, Z => n2193);
   U663 : HS65_LH_OAI22X6 port map( A => n6297, B => n296, C => n822, D => 
                           n6301, Z => n2194);
   U664 : HS65_LH_OAI22X6 port map( A => n6297, B => n295, C => n821, D => 
                           n6301, Z => n2195);
   U665 : HS65_LH_OAI22X6 port map( A => n6297, B => n294, C => n820, D => 
                           n6301, Z => n2196);
   U666 : HS65_LH_OAI22X6 port map( A => n6297, B => n293, C => n819, D => 
                           n6301, Z => n2197);
   U667 : HS65_LH_OAI22X6 port map( A => n6297, B => n292, C => n818, D => 
                           n6301, Z => n2198);
   U668 : HS65_LH_OAI22X6 port map( A => n6297, B => n291, C => n817, D => 
                           n6301, Z => n2199);
   U669 : HS65_LH_OAI22X6 port map( A => n6297, B => n290, C => n816, D => 
                           n6301, Z => n2200);
   U670 : HS65_LH_OAI22X6 port map( A => n6297, B => n289, C => n815, D => 
                           n6301, Z => n2201);
   U671 : HS65_LH_OAI22X6 port map( A => n846, B => n6239, C => n6238, D => 
                           n448, Z => n1786);
   U672 : HS65_LH_OAI22X6 port map( A => n846, B => n6259, C => n6258, D => 
                           n416, Z => n1914);
   U673 : HS65_LH_OAI22X6 port map( A => n846, B => n6264, C => n6263, D => 
                           n384, Z => n1946);
   U674 : HS65_LH_OAI22X6 port map( A => n846, B => n6209, C => n6208, D => 
                           n512, Z => n1594);
   U675 : HS65_LH_OAI22X6 port map( A => n845, B => n6240, C => n6237, D => 
                           n447, Z => n1787);
   U676 : HS65_LH_OAI22X6 port map( A => n844, B => n6240, C => n6238, D => 
                           n446, Z => n1788);
   U677 : HS65_LH_OAI22X6 port map( A => n843, B => n6240, C => n6237, D => 
                           n445, Z => n1789);
   U678 : HS65_LH_OAI22X6 port map( A => n842, B => n6240, C => n6238, D => 
                           n444, Z => n1790);
   U679 : HS65_LH_OAI22X6 port map( A => n841, B => n6240, C => n6237, D => 
                           n443, Z => n1791);
   U680 : HS65_LH_OAI22X6 port map( A => n840, B => n6240, C => n6238, D => 
                           n442, Z => n1792);
   U681 : HS65_LH_OAI22X6 port map( A => n839, B => n6240, C => n6238, D => 
                           n441, Z => n1793);
   U682 : HS65_LH_OAI22X6 port map( A => n838, B => n6240, C => n6238, D => 
                           n440, Z => n1794);
   U683 : HS65_LH_OAI22X6 port map( A => n837, B => n6240, C => n6238, D => 
                           n439, Z => n1795);
   U684 : HS65_LH_OAI22X6 port map( A => n836, B => n6240, C => n6238, D => 
                           n438, Z => n1796);
   U685 : HS65_LH_OAI22X6 port map( A => n835, B => n6240, C => n6238, D => 
                           n437, Z => n1797);
   U686 : HS65_LH_OAI22X6 port map( A => n834, B => n6240, C => n6238, D => 
                           n436, Z => n1798);
   U687 : HS65_LH_OAI22X6 port map( A => n833, B => n6240, C => n6238, D => 
                           n435, Z => n1799);
   U688 : HS65_LH_OAI22X6 port map( A => n832, B => n6240, C => n6238, D => 
                           n434, Z => n1800);
   U689 : HS65_LH_OAI22X6 port map( A => n831, B => n6240, C => n6238, D => 
                           n433, Z => n1801);
   U690 : HS65_LH_OAI22X6 port map( A => n830, B => n6240, C => n6238, D => 
                           n432, Z => n1802);
   U691 : HS65_LH_OAI22X6 port map( A => n829, B => n6240, C => n6238, D => 
                           n431, Z => n1803);
   U692 : HS65_LH_OAI22X6 port map( A => n828, B => n6240, C => n6238, D => 
                           n430, Z => n1804);
   U693 : HS65_LH_OAI22X6 port map( A => n845, B => n6260, C => n6257, D => 
                           n415, Z => n1915);
   U694 : HS65_LH_OAI22X6 port map( A => n844, B => n6260, C => n6258, D => 
                           n414, Z => n1916);
   U695 : HS65_LH_OAI22X6 port map( A => n843, B => n6260, C => n6257, D => 
                           n413, Z => n1917);
   U696 : HS65_LH_OAI22X6 port map( A => n842, B => n6260, C => n6258, D => 
                           n412, Z => n1918);
   U697 : HS65_LH_OAI22X6 port map( A => n841, B => n6260, C => n6257, D => 
                           n411, Z => n1919);
   U698 : HS65_LH_OAI22X6 port map( A => n840, B => n6260, C => n6258, D => 
                           n410, Z => n1920);
   U699 : HS65_LH_OAI22X6 port map( A => n839, B => n6260, C => n6258, D => 
                           n409, Z => n1921);
   U700 : HS65_LH_OAI22X6 port map( A => n838, B => n6260, C => n6258, D => 
                           n408, Z => n1922);
   U701 : HS65_LH_OAI22X6 port map( A => n837, B => n6260, C => n6258, D => 
                           n407, Z => n1923);
   U702 : HS65_LH_OAI22X6 port map( A => n836, B => n6260, C => n6258, D => 
                           n406, Z => n1924);
   U703 : HS65_LH_OAI22X6 port map( A => n835, B => n6260, C => n6258, D => 
                           n405, Z => n1925);
   U704 : HS65_LH_OAI22X6 port map( A => n834, B => n6260, C => n6258, D => 
                           n404, Z => n1926);
   U705 : HS65_LH_OAI22X6 port map( A => n833, B => n6260, C => n6258, D => 
                           n403, Z => n1927);
   U706 : HS65_LH_OAI22X6 port map( A => n832, B => n6260, C => n6258, D => 
                           n402, Z => n1928);
   U707 : HS65_LH_OAI22X6 port map( A => n831, B => n6260, C => n6258, D => 
                           n401, Z => n1929);
   U708 : HS65_LH_OAI22X6 port map( A => n830, B => n6260, C => n6258, D => 
                           n400, Z => n1930);
   U709 : HS65_LH_OAI22X6 port map( A => n829, B => n6260, C => n6258, D => 
                           n399, Z => n1931);
   U710 : HS65_LH_OAI22X6 port map( A => n828, B => n6260, C => n6258, D => 
                           n398, Z => n1932);
   U711 : HS65_LH_OAI22X6 port map( A => n845, B => n6265, C => n6262, D => 
                           n383, Z => n1947);
   U712 : HS65_LH_OAI22X6 port map( A => n844, B => n6265, C => n6263, D => 
                           n382, Z => n1948);
   U713 : HS65_LH_OAI22X6 port map( A => n843, B => n6265, C => n6262, D => 
                           n381, Z => n1949);
   U714 : HS65_LH_OAI22X6 port map( A => n842, B => n6265, C => n6263, D => 
                           n380, Z => n1950);
   U715 : HS65_LH_OAI22X6 port map( A => n841, B => n6265, C => n6262, D => 
                           n379, Z => n1951);
   U716 : HS65_LH_OAI22X6 port map( A => n840, B => n6265, C => n6263, D => 
                           n378, Z => n1952);
   U717 : HS65_LH_OAI22X6 port map( A => n839, B => n6265, C => n6263, D => 
                           n377, Z => n1953);
   U718 : HS65_LH_OAI22X6 port map( A => n838, B => n6265, C => n6263, D => 
                           n376, Z => n1954);
   U719 : HS65_LH_OAI22X6 port map( A => n837, B => n6265, C => n6263, D => 
                           n375, Z => n1955);
   U720 : HS65_LH_OAI22X6 port map( A => n836, B => n6265, C => n6263, D => 
                           n374, Z => n1956);
   U721 : HS65_LH_OAI22X6 port map( A => n835, B => n6265, C => n6263, D => 
                           n373, Z => n1957);
   U722 : HS65_LH_OAI22X6 port map( A => n834, B => n6265, C => n6263, D => 
                           n372, Z => n1958);
   U723 : HS65_LH_OAI22X6 port map( A => n833, B => n6265, C => n6263, D => 
                           n371, Z => n1959);
   U724 : HS65_LH_OAI22X6 port map( A => n832, B => n6265, C => n6263, D => 
                           n370, Z => n1960);
   U725 : HS65_LH_OAI22X6 port map( A => n831, B => n6265, C => n6263, D => 
                           n369, Z => n1961);
   U726 : HS65_LH_OAI22X6 port map( A => n830, B => n6265, C => n6263, D => 
                           n368, Z => n1962);
   U727 : HS65_LH_OAI22X6 port map( A => n829, B => n6265, C => n6263, D => 
                           n367, Z => n1963);
   U728 : HS65_LH_OAI22X6 port map( A => n828, B => n6265, C => n6263, D => 
                           n366, Z => n1964);
   U729 : HS65_LH_OAI22X6 port map( A => n845, B => n6210, C => n6207, D => 
                           n511, Z => n1595);
   U730 : HS65_LH_OAI22X6 port map( A => n844, B => n6210, C => n6208, D => 
                           n510, Z => n1596);
   U731 : HS65_LH_OAI22X6 port map( A => n843, B => n6210, C => n6207, D => 
                           n509, Z => n1597);
   U732 : HS65_LH_OAI22X6 port map( A => n842, B => n6210, C => n6208, D => 
                           n508, Z => n1598);
   U733 : HS65_LH_OAI22X6 port map( A => n841, B => n6210, C => n6207, D => 
                           n507, Z => n1599);
   U734 : HS65_LH_OAI22X6 port map( A => n840, B => n6210, C => n6208, D => 
                           n506, Z => n1600);
   U735 : HS65_LH_OAI22X6 port map( A => n839, B => n6210, C => n6208, D => 
                           n505, Z => n1601);
   U736 : HS65_LH_OAI22X6 port map( A => n838, B => n6210, C => n6208, D => 
                           n504, Z => n1602);
   U737 : HS65_LH_OAI22X6 port map( A => n837, B => n6210, C => n6208, D => 
                           n503, Z => n1603);
   U738 : HS65_LH_OAI22X6 port map( A => n836, B => n6210, C => n6208, D => 
                           n502, Z => n1604);
   U739 : HS65_LH_OAI22X6 port map( A => n835, B => n6210, C => n6208, D => 
                           n501, Z => n1605);
   U740 : HS65_LH_OAI22X6 port map( A => n834, B => n6210, C => n6208, D => 
                           n500, Z => n1606);
   U741 : HS65_LH_OAI22X6 port map( A => n833, B => n6210, C => n6208, D => 
                           n499, Z => n1607);
   U742 : HS65_LH_OAI22X6 port map( A => n832, B => n6210, C => n6208, D => 
                           n498, Z => n1608);
   U743 : HS65_LH_OAI22X6 port map( A => n831, B => n6210, C => n6208, D => 
                           n497, Z => n1609);
   U744 : HS65_LH_OAI22X6 port map( A => n830, B => n6210, C => n6208, D => 
                           n496, Z => n1610);
   U745 : HS65_LH_OAI22X6 port map( A => n829, B => n6210, C => n6208, D => 
                           n495, Z => n1611);
   U746 : HS65_LH_OAI22X6 port map( A => n828, B => n6210, C => n6208, D => 
                           n494, Z => n1612);
   U747 : HS65_LH_OAI22X6 port map( A => n827, B => n6241, C => n6237, D => 
                           n429, Z => n1805);
   U748 : HS65_LH_OAI22X6 port map( A => n826, B => n6241, C => n6237, D => 
                           n428, Z => n1806);
   U749 : HS65_LH_OAI22X6 port map( A => n825, B => n6241, C => n6237, D => 
                           n427, Z => n1807);
   U750 : HS65_LH_OAI22X6 port map( A => n824, B => n6241, C => n6237, D => 
                           n426, Z => n1808);
   U751 : HS65_LH_OAI22X6 port map( A => n823, B => n6241, C => n6237, D => 
                           n425, Z => n1809);
   U752 : HS65_LH_OAI22X6 port map( A => n822, B => n6241, C => n6237, D => 
                           n424, Z => n1810);
   U753 : HS65_LH_OAI22X6 port map( A => n821, B => n6241, C => n6237, D => 
                           n423, Z => n1811);
   U754 : HS65_LH_OAI22X6 port map( A => n820, B => n6241, C => n6237, D => 
                           n422, Z => n1812);
   U755 : HS65_LH_OAI22X6 port map( A => n819, B => n6241, C => n6237, D => 
                           n421, Z => n1813);
   U756 : HS65_LH_OAI22X6 port map( A => n818, B => n6241, C => n6237, D => 
                           n420, Z => n1814);
   U757 : HS65_LH_OAI22X6 port map( A => n817, B => n6241, C => n6237, D => 
                           n419, Z => n1815);
   U758 : HS65_LH_OAI22X6 port map( A => n816, B => n6241, C => n6237, D => 
                           n418, Z => n1816);
   U759 : HS65_LH_OAI22X6 port map( A => n815, B => n6241, C => n6237, D => 
                           n417, Z => n1817);
   U760 : HS65_LH_OAI22X6 port map( A => n827, B => n6261, C => n6257, D => 
                           n397, Z => n1933);
   U761 : HS65_LH_OAI22X6 port map( A => n826, B => n6261, C => n6257, D => 
                           n396, Z => n1934);
   U762 : HS65_LH_OAI22X6 port map( A => n825, B => n6261, C => n6257, D => 
                           n395, Z => n1935);
   U763 : HS65_LH_OAI22X6 port map( A => n824, B => n6261, C => n6257, D => 
                           n394, Z => n1936);
   U764 : HS65_LH_OAI22X6 port map( A => n823, B => n6261, C => n6257, D => 
                           n393, Z => n1937);
   U765 : HS65_LH_OAI22X6 port map( A => n822, B => n6261, C => n6257, D => 
                           n392, Z => n1938);
   U766 : HS65_LH_OAI22X6 port map( A => n821, B => n6261, C => n6257, D => 
                           n391, Z => n1939);
   U767 : HS65_LH_OAI22X6 port map( A => n820, B => n6261, C => n6257, D => 
                           n390, Z => n1940);
   U768 : HS65_LH_OAI22X6 port map( A => n819, B => n6261, C => n6257, D => 
                           n389, Z => n1941);
   U769 : HS65_LH_OAI22X6 port map( A => n818, B => n6261, C => n6257, D => 
                           n388, Z => n1942);
   U770 : HS65_LH_OAI22X6 port map( A => n817, B => n6261, C => n6257, D => 
                           n387, Z => n1943);
   U771 : HS65_LH_OAI22X6 port map( A => n816, B => n6261, C => n6257, D => 
                           n386, Z => n1944);
   U772 : HS65_LH_OAI22X6 port map( A => n815, B => n6261, C => n6257, D => 
                           n385, Z => n1945);
   U773 : HS65_LH_OAI22X6 port map( A => n827, B => n6266, C => n6262, D => 
                           n365, Z => n1965);
   U774 : HS65_LH_OAI22X6 port map( A => n826, B => n6266, C => n6262, D => 
                           n364, Z => n1966);
   U775 : HS65_LH_OAI22X6 port map( A => n825, B => n6266, C => n6262, D => 
                           n363, Z => n1967);
   U776 : HS65_LH_OAI22X6 port map( A => n824, B => n6266, C => n6262, D => 
                           n362, Z => n1968);
   U777 : HS65_LH_OAI22X6 port map( A => n823, B => n6266, C => n6262, D => 
                           n361, Z => n1969);
   U778 : HS65_LH_OAI22X6 port map( A => n822, B => n6266, C => n6262, D => 
                           n360, Z => n1970);
   U779 : HS65_LH_OAI22X6 port map( A => n821, B => n6266, C => n6262, D => 
                           n359, Z => n1971);
   U780 : HS65_LH_OAI22X6 port map( A => n820, B => n6266, C => n6262, D => 
                           n358, Z => n1972);
   U781 : HS65_LH_OAI22X6 port map( A => n819, B => n6266, C => n6262, D => 
                           n357, Z => n1973);
   U782 : HS65_LH_OAI22X6 port map( A => n818, B => n6266, C => n6262, D => 
                           n356, Z => n1974);
   U783 : HS65_LH_OAI22X6 port map( A => n817, B => n6266, C => n6262, D => 
                           n355, Z => n1975);
   U784 : HS65_LH_OAI22X6 port map( A => n816, B => n6266, C => n6262, D => 
                           n354, Z => n1976);
   U785 : HS65_LH_OAI22X6 port map( A => n815, B => n6266, C => n6262, D => 
                           n353, Z => n1977);
   U786 : HS65_LH_OAI22X6 port map( A => n827, B => n6211, C => n6207, D => 
                           n493, Z => n1613);
   U787 : HS65_LH_OAI22X6 port map( A => n826, B => n6211, C => n6207, D => 
                           n492, Z => n1614);
   U788 : HS65_LH_OAI22X6 port map( A => n825, B => n6211, C => n6207, D => 
                           n491, Z => n1615);
   U789 : HS65_LH_OAI22X6 port map( A => n824, B => n6211, C => n6207, D => 
                           n490, Z => n1616);
   U790 : HS65_LH_OAI22X6 port map( A => n823, B => n6211, C => n6207, D => 
                           n489, Z => n1617);
   U791 : HS65_LH_OAI22X6 port map( A => n822, B => n6211, C => n6207, D => 
                           n488, Z => n1618);
   U792 : HS65_LH_OAI22X6 port map( A => n821, B => n6211, C => n6207, D => 
                           n487, Z => n1619);
   U793 : HS65_LH_OAI22X6 port map( A => n820, B => n6211, C => n6207, D => 
                           n486, Z => n1620);
   U794 : HS65_LH_OAI22X6 port map( A => n819, B => n6211, C => n6207, D => 
                           n485, Z => n1621);
   U795 : HS65_LH_OAI22X6 port map( A => n818, B => n6211, C => n6207, D => 
                           n484, Z => n1622);
   U796 : HS65_LH_OAI22X6 port map( A => n817, B => n6211, C => n6207, D => 
                           n483, Z => n1623);
   U797 : HS65_LH_OAI22X6 port map( A => n816, B => n6211, C => n6207, D => 
                           n482, Z => n1624);
   U798 : HS65_LH_OAI22X6 port map( A => n815, B => n6211, C => n6207, D => 
                           n481, Z => n1625);
   U799 : HS65_LH_NAND2X7 port map( A => n1327, B => n1324, Z => n885);
   U800 : HS65_LH_NAND2X7 port map( A => n1328, B => n1337, Z => n879);
   U801 : HS65_LH_NAND2X7 port map( A => n2822, B => n2807, Z => n1375);
   U802 : HS65_LH_NAND2X7 port map( A => n2809, B => n2807, Z => n1371);
   U803 : HS65_LH_NAND2X7 port map( A => n2819, B => n2807, Z => n1370);
   U804 : HS65_LH_NAND2X7 port map( A => n2805, B => n2807, Z => n1350);
   U805 : HS65_LH_NAND2X7 port map( A => n1322, B => n1323, Z => n860);
   U806 : HS65_LH_NAND2X7 port map( A => n2805, B => n2806, Z => n1351);
   U807 : HS65_LH_NAND2X7 port map( A => n2822, B => n2808, Z => n1376);
   U808 : HS65_LH_NAND2X7 port map( A => n1330, B => n1328, Z => n884);
   U809 : HS65_LH_NAND2X7 port map( A => n1331, B => n1328, Z => n880);
   U810 : HS65_LH_NAND2X7 port map( A => n1324, B => n1325, Z => n859);
   U811 : HS65_LH_NAND2X7 port map( A => n2829, B => n2825, Z => n2828);
   U812 : HS65_LH_NAND2X7 port map( A => n2835, B => n2825, Z => n2834);
   U813 : HS65_LH_NAND2X7 port map( A => n2831, B => n2825, Z => n2830);
   U814 : HS65_LH_NAND2X7 port map( A => n2833, B => n2825, Z => n2832);
   U815 : HS65_LH_NAND2X7 port map( A => n2839, B => n2825, Z => n2838);
   U816 : HS65_LH_NAND2X7 port map( A => n2837, B => n2825, Z => n2836);
   U817 : HS65_LH_NAND2X7 port map( A => n2841, B => n2839, Z => n2848);
   U818 : HS65_LH_NAND2X7 port map( A => n2841, B => n2837, Z => n2847);
   U819 : HS65_LH_NAND2X7 port map( A => n2841, B => n2835, Z => n2846);
   U820 : HS65_LH_NAND2X7 port map( A => n2850, B => n2839, Z => n2857);
   U821 : HS65_LH_NAND2X7 port map( A => n2850, B => n2837, Z => n2856);
   U822 : HS65_LH_NAND2X7 port map( A => n2850, B => n2827, Z => n2851);
   U823 : HS65_LH_NAND2X7 port map( A => n2850, B => n2824, Z => n2849);
   U824 : HS65_LH_NAND2X7 port map( A => n2850, B => n2835, Z => n2855);
   U825 : HS65_LH_NAND2X7 port map( A => n2850, B => n2831, Z => n2853);
   U826 : HS65_LH_NOR3X4 port map( A => n813, B => n814, C => n812, Z => n2824)
                           ;
   U827 : HS65_LH_NAND2X7 port map( A => n2859, B => n2827, Z => n2860);
   U828 : HS65_LH_NOR3X4 port map( A => n775, B => n774, C => n778, Z => n1330)
                           ;
   U829 : HS65_LH_NOR3X4 port map( A => n769, B => n770, C => n773, Z => n2819)
                           ;
   U830 : HS65_LH_NOR2X6 port map( A => n776, B => n777, Z => n1323);
   U831 : HS65_LH_NOR2X6 port map( A => n771, B => n772, Z => n2806);
   U832 : HS65_LH_OAI22X6 port map( A => n6469, B => n406, C => n6466, D => 
                           n374, Z => n1312);
   U833 : HS65_LH_BFX9 port map( A => n847, Z => n6531);
   U834 : HS65_LH_BFX9 port map( A => n847, Z => n6530);
   U835 : HS65_LH_BFX9 port map( A => n848, Z => n6525);
   U836 : HS65_LH_BFX9 port map( A => n848, Z => n6527);
   U837 : HS65_LH_BFX9 port map( A => n848, Z => n6526);
   U838 : HS65_LH_BFX9 port map( A => n847, Z => n6528);
   U839 : HS65_LH_BFX9 port map( A => n847, Z => n6529);
   U840 : HS65_LH_BFX9 port map( A => n847, Z => n6532);
   U841 : HS65_LH_BFX9 port map( A => n848, Z => n6523);
   U842 : HS65_LH_BFX9 port map( A => n848, Z => n6524);
   U843 : HS65_LH_OAI21X3 port map( A => n6525, B => n846, C => n1314, Z => 
                           regfile_o(0));
   U844 : HS65_LH_OAI21X3 port map( A => n1315, B => n1316, C => n6523, Z => 
                           n1314);
   U845 : HS65_LH_NAND4ABX3 port map( A => n1317, B => n1318, C => n1319, D => 
                           n1320, Z => n1316);
   U846 : HS65_LH_NAND4ABX3 port map( A => n1332, B => n1333, C => n1334, D => 
                           n1335, Z => n1315);
   U847 : HS65_LH_OAI21X3 port map( A => n6527, B => n845, C => n1160, Z => 
                           regfile_o(1));
   U848 : HS65_LH_OAI21X3 port map( A => n1161, B => n1162, C => n6524, Z => 
                           n1160);
   U849 : HS65_LH_NAND4ABX3 port map( A => n1163, B => n1164, C => n1165, D => 
                           n1166, Z => n1162);
   U850 : HS65_LH_NAND4ABX3 port map( A => n1168, B => n1169, C => n1170, D => 
                           n1171, Z => n1161);
   U851 : HS65_LH_OAI21X3 port map( A => n6526, B => n844, C => n1006, Z => 
                           regfile_o(2));
   U852 : HS65_LH_OAI21X3 port map( A => n1007, B => n1008, C => n6525, Z => 
                           n1006);
   U853 : HS65_LH_NAND4ABX3 port map( A => n1009, B => n1010, C => n1011, D => 
                           n1012, Z => n1008);
   U854 : HS65_LH_NAND4ABX3 port map( A => n1014, B => n1015, C => n1016, D => 
                           n1017, Z => n1007);
   U855 : HS65_LH_OAI21X3 port map( A => n6525, B => n843, C => n964, Z => 
                           regfile_o(3));
   U856 : HS65_LH_OAI21X3 port map( A => n965, B => n966, C => n6524, Z => n964
                           );
   U857 : HS65_LH_NAND4ABX3 port map( A => n967, B => n968, C => n969, D => 
                           n970, Z => n966);
   U858 : HS65_LH_NAND4ABX3 port map( A => n972, B => n973, C => n974, D => 
                           n975, Z => n965);
   U859 : HS65_LH_OAI21X3 port map( A => n6526, B => n842, C => n950, Z => 
                           regfile_o(4));
   U860 : HS65_LH_OAI21X3 port map( A => n951, B => n952, C => n6524, Z => n950
                           );
   U861 : HS65_LH_NAND4ABX3 port map( A => n953, B => n954, C => n955, D => 
                           n956, Z => n952);
   U862 : HS65_LH_NAND4ABX3 port map( A => n958, B => n959, C => n960, D => 
                           n961, Z => n951);
   U863 : HS65_LH_OAI21X3 port map( A => n6525, B => n841, C => n936, Z => 
                           regfile_o(5));
   U864 : HS65_LH_OAI21X3 port map( A => n937, B => n938, C => n6524, Z => n936
                           );
   U865 : HS65_LH_NAND4ABX3 port map( A => n939, B => n940, C => n941, D => 
                           n942, Z => n938);
   U866 : HS65_LH_NAND4ABX3 port map( A => n944, B => n945, C => n946, D => 
                           n947, Z => n937);
   U867 : HS65_LH_OAI21X3 port map( A => n6525, B => n840, C => n922, Z => 
                           regfile_o(6));
   U868 : HS65_LH_OAI21X3 port map( A => n923, B => n924, C => n6523, Z => n922
                           );
   U869 : HS65_LH_NAND4ABX3 port map( A => n925, B => n926, C => n927, D => 
                           n928, Z => n924);
   U870 : HS65_LH_NAND4ABX3 port map( A => n930, B => n931, C => n932, D => 
                           n933, Z => n923);
   U871 : HS65_LH_OAI21X3 port map( A => n6526, B => n839, C => n908, Z => 
                           regfile_o(7));
   U872 : HS65_LH_OAI21X3 port map( A => n909, B => n910, C => n6523, Z => n908
                           );
   U873 : HS65_LH_NAND4ABX3 port map( A => n911, B => n912, C => n913, D => 
                           n914, Z => n910);
   U874 : HS65_LH_NAND4ABX3 port map( A => n916, B => n917, C => n918, D => 
                           n919, Z => n909);
   U875 : HS65_LH_OAI21X3 port map( A => n6525, B => n838, C => n894, Z => 
                           regfile_o(8));
   U876 : HS65_LH_OAI21X3 port map( A => n895, B => n896, C => n6523, Z => n894
                           );
   U877 : HS65_LH_NAND4ABX3 port map( A => n897, B => n898, C => n899, D => 
                           n900, Z => n896);
   U878 : HS65_LH_NAND4ABX3 port map( A => n902, B => n903, C => n904, D => 
                           n905, Z => n895);
   U879 : HS65_LH_OAI21X3 port map( A => n6526, B => n837, C => n849, Z => 
                           regfile_o(9));
   U880 : HS65_LH_OAI21X3 port map( A => n850, B => n851, C => n6523, Z => n849
                           );
   U881 : HS65_LH_NAND4ABX3 port map( A => n852, B => n853, C => n854, D => 
                           n855, Z => n851);
   U882 : HS65_LH_NAND4ABX3 port map( A => n872, B => n873, C => n874, D => 
                           n875, Z => n850);
   U883 : HS65_LH_OAI21X3 port map( A => n848, B => n836, C => n1300, Z => 
                           regfile_o(10));
   U884 : HS65_LH_OAI21X3 port map( A => n1301, B => n1302, C => n6523, Z => 
                           n1300);
   U885 : HS65_LH_NAND4ABX3 port map( A => n1303, B => n1304, C => n1305, D => 
                           n1306, Z => n1302);
   U886 : HS65_LH_OAI21X3 port map( A => n6527, B => n835, C => n1286, Z => 
                           regfile_o(11));
   U887 : HS65_LH_OAI21X3 port map( A => n1287, B => n1288, C => n6523, Z => 
                           n1286);
   U888 : HS65_LH_NAND4ABX3 port map( A => n1289, B => n1290, C => n1291, D => 
                           n1292, Z => n1288);
   U889 : HS65_LH_NAND4ABX3 port map( A => n1294, B => n1295, C => n1296, D => 
                           n1297, Z => n1287);
   U890 : HS65_LH_OAI21X3 port map( A => n6527, B => n834, C => n1272, Z => 
                           regfile_o(12));
   U891 : HS65_LH_OAI21X3 port map( A => n1273, B => n1274, C => n6523, Z => 
                           n1272);
   U892 : HS65_LH_NAND4ABX3 port map( A => n1275, B => n1276, C => n1277, D => 
                           n1278, Z => n1274);
   U893 : HS65_LH_NAND4ABX3 port map( A => n1280, B => n1281, C => n1282, D => 
                           n1283, Z => n1273);
   U894 : HS65_LH_OAI21X3 port map( A => n6527, B => n833, C => n1258, Z => 
                           regfile_o(13));
   U895 : HS65_LH_OAI21X3 port map( A => n1259, B => n1260, C => n6523, Z => 
                           n1258);
   U896 : HS65_LH_NAND4ABX3 port map( A => n1261, B => n1262, C => n1263, D => 
                           n1264, Z => n1260);
   U897 : HS65_LH_NAND4ABX3 port map( A => n1266, B => n1267, C => n1268, D => 
                           n1269, Z => n1259);
   U898 : HS65_LH_OAI21X3 port map( A => n6527, B => n832, C => n1244, Z => 
                           regfile_o(14));
   U899 : HS65_LH_OAI21X3 port map( A => n1245, B => n1246, C => n6523, Z => 
                           n1244);
   U900 : HS65_LH_NAND4ABX3 port map( A => n1247, B => n1248, C => n1249, D => 
                           n1250, Z => n1246);
   U901 : HS65_LH_NAND4ABX3 port map( A => n1252, B => n1253, C => n1254, D => 
                           n1255, Z => n1245);
   U902 : HS65_LH_OAI21X3 port map( A => n6527, B => n831, C => n1230, Z => 
                           regfile_o(15));
   U903 : HS65_LH_OAI21X3 port map( A => n1231, B => n1232, C => n6523, Z => 
                           n1230);
   U904 : HS65_LH_NAND4ABX3 port map( A => n1233, B => n1234, C => n1235, D => 
                           n1236, Z => n1232);
   U905 : HS65_LH_NAND4ABX3 port map( A => n1238, B => n1239, C => n1240, D => 
                           n1241, Z => n1231);
   U906 : HS65_LH_OAI21X3 port map( A => n6527, B => n830, C => n1216, Z => 
                           regfile_o(16));
   U907 : HS65_LH_OAI21X3 port map( A => n1217, B => n1218, C => n6523, Z => 
                           n1216);
   U908 : HS65_LH_NAND4ABX3 port map( A => n1219, B => n1220, C => n1221, D => 
                           n1222, Z => n1218);
   U909 : HS65_LH_NAND4ABX3 port map( A => n1224, B => n1225, C => n1226, D => 
                           n1227, Z => n1217);
   U910 : HS65_LH_OAI21X3 port map( A => n6527, B => n829, C => n1202, Z => 
                           regfile_o(17));
   U911 : HS65_LH_OAI21X3 port map( A => n1203, B => n1204, C => n6524, Z => 
                           n1202);
   U912 : HS65_LH_NAND4ABX3 port map( A => n1205, B => n1206, C => n1207, D => 
                           n1208, Z => n1204);
   U913 : HS65_LH_NAND4ABX3 port map( A => n1210, B => n1211, C => n1212, D => 
                           n1213, Z => n1203);
   U914 : HS65_LH_OAI21X3 port map( A => n6527, B => n828, C => n1188, Z => 
                           regfile_o(18));
   U915 : HS65_LH_OAI21X3 port map( A => n1189, B => n1190, C => n6524, Z => 
                           n1188);
   U916 : HS65_LH_NAND4ABX3 port map( A => n1191, B => n1192, C => n1193, D => 
                           n1194, Z => n1190);
   U917 : HS65_LH_NAND4ABX3 port map( A => n1196, B => n1197, C => n1198, D => 
                           n1199, Z => n1189);
   U918 : HS65_LH_OAI21X3 port map( A => n6527, B => n827, C => n1174, Z => 
                           regfile_o(19));
   U919 : HS65_LH_OAI21X3 port map( A => n1175, B => n1176, C => n6524, Z => 
                           n1174);
   U920 : HS65_LH_NAND4ABX3 port map( A => n1177, B => n1178, C => n1179, D => 
                           n1180, Z => n1176);
   U921 : HS65_LH_NAND4ABX3 port map( A => n1182, B => n1183, C => n1184, D => 
                           n1185, Z => n1175);
   U922 : HS65_LH_OAI21X3 port map( A => n6527, B => n826, C => n1146, Z => 
                           regfile_o(20));
   U923 : HS65_LH_OAI21X3 port map( A => n1147, B => n1148, C => n6524, Z => 
                           n1146);
   U924 : HS65_LH_NAND4ABX3 port map( A => n1149, B => n1150, C => n1151, D => 
                           n1152, Z => n1148);
   U925 : HS65_LH_NAND4ABX3 port map( A => n1154, B => n1155, C => n1156, D => 
                           n1157, Z => n1147);
   U926 : HS65_LH_OAI21X3 port map( A => n6527, B => n825, C => n1132, Z => 
                           regfile_o(21));
   U927 : HS65_LH_OAI21X3 port map( A => n1133, B => n1134, C => n6524, Z => 
                           n1132);
   U928 : HS65_LH_NAND4ABX3 port map( A => n1135, B => n1136, C => n1137, D => 
                           n1138, Z => n1134);
   U929 : HS65_LH_NAND4ABX3 port map( A => n1140, B => n1141, C => n1142, D => 
                           n1143, Z => n1133);
   U930 : HS65_LH_OAI21X3 port map( A => n6527, B => n824, C => n1118, Z => 
                           regfile_o(22));
   U931 : HS65_LH_OAI21X3 port map( A => n1119, B => n1120, C => n6524, Z => 
                           n1118);
   U932 : HS65_LH_NAND4ABX3 port map( A => n1121, B => n1122, C => n1123, D => 
                           n1124, Z => n1120);
   U933 : HS65_LH_NAND4ABX3 port map( A => n1126, B => n1127, C => n1128, D => 
                           n1129, Z => n1119);
   U934 : HS65_LH_OAI21X3 port map( A => n6526, B => n823, C => n1104, Z => 
                           regfile_o(23));
   U935 : HS65_LH_OAI21X3 port map( A => n1105, B => n1106, C => n6524, Z => 
                           n1104);
   U936 : HS65_LH_NAND4ABX3 port map( A => n1107, B => n1108, C => n1109, D => 
                           n1110, Z => n1106);
   U937 : HS65_LH_NAND4ABX3 port map( A => n1112, B => n1113, C => n1114, D => 
                           n1115, Z => n1105);
   U938 : HS65_LH_OAI21X3 port map( A => n6526, B => n822, C => n1090, Z => 
                           regfile_o(24));
   U939 : HS65_LH_OAI21X3 port map( A => n1091, B => n1092, C => n6525, Z => 
                           n1090);
   U940 : HS65_LH_NAND4ABX3 port map( A => n1093, B => n1094, C => n1095, D => 
                           n1096, Z => n1092);
   U941 : HS65_LH_NAND4ABX3 port map( A => n1098, B => n1099, C => n1100, D => 
                           n1101, Z => n1091);
   U942 : HS65_LH_OAI21X3 port map( A => n6526, B => n821, C => n1076, Z => 
                           regfile_o(25));
   U943 : HS65_LH_OAI21X3 port map( A => n1077, B => n1078, C => n6525, Z => 
                           n1076);
   U944 : HS65_LH_NAND4ABX3 port map( A => n1079, B => n1080, C => n1081, D => 
                           n1082, Z => n1078);
   U945 : HS65_LH_NAND4ABX3 port map( A => n1084, B => n1085, C => n1086, D => 
                           n1087, Z => n1077);
   U946 : HS65_LH_OAI21X3 port map( A => n6526, B => n820, C => n1062, Z => 
                           regfile_o(26));
   U947 : HS65_LH_OAI21X3 port map( A => n1063, B => n1064, C => n6524, Z => 
                           n1062);
   U948 : HS65_LH_NAND4ABX3 port map( A => n1065, B => n1066, C => n1067, D => 
                           n1068, Z => n1064);
   U949 : HS65_LH_NAND4ABX3 port map( A => n1070, B => n1071, C => n1072, D => 
                           n1073, Z => n1063);
   U950 : HS65_LH_OAI21X3 port map( A => n6526, B => n819, C => n1048, Z => 
                           regfile_o(27));
   U951 : HS65_LH_OAI21X3 port map( A => n1049, B => n1050, C => n6525, Z => 
                           n1048);
   U952 : HS65_LH_NAND4ABX3 port map( A => n1051, B => n1052, C => n1053, D => 
                           n1054, Z => n1050);
   U953 : HS65_LH_NAND4ABX3 port map( A => n1056, B => n1057, C => n1058, D => 
                           n1059, Z => n1049);
   U954 : HS65_LH_OAI21X3 port map( A => n6526, B => n818, C => n1034, Z => 
                           regfile_o(28));
   U955 : HS65_LH_OAI21X3 port map( A => n1035, B => n1036, C => n6525, Z => 
                           n1034);
   U956 : HS65_LH_NAND4ABX3 port map( A => n1037, B => n1038, C => n1039, D => 
                           n1040, Z => n1036);
   U957 : HS65_LH_NAND4ABX3 port map( A => n1042, B => n1043, C => n1044, D => 
                           n1045, Z => n1035);
   U958 : HS65_LH_OAI21X3 port map( A => n6526, B => n817, C => n1020, Z => 
                           regfile_o(29));
   U959 : HS65_LH_OAI21X3 port map( A => n1021, B => n1022, C => n6525, Z => 
                           n1020);
   U960 : HS65_LH_NAND4ABX3 port map( A => n1023, B => n1024, C => n1025, D => 
                           n1026, Z => n1022);
   U961 : HS65_LH_NAND4ABX3 port map( A => n1028, B => n1029, C => n1030, D => 
                           n1031, Z => n1021);
   U962 : HS65_LH_OAI21X3 port map( A => n6526, B => n816, C => n992, Z => 
                           regfile_o(30));
   U963 : HS65_LH_OAI21X3 port map( A => n993, B => n994, C => n6525, Z => n992
                           );
   U964 : HS65_LH_NAND4ABX3 port map( A => n995, B => n996, C => n997, D => 
                           n998, Z => n994);
   U965 : HS65_LH_NAND4ABX3 port map( A => n1000, B => n1001, C => n1002, D => 
                           n1003, Z => n993);
   U966 : HS65_LH_OAI21X3 port map( A => n6526, B => n815, C => n978, Z => 
                           regfile_o(31));
   U967 : HS65_LH_OAI21X3 port map( A => n979, B => n980, C => n6525, Z => n978
                           );
   U968 : HS65_LH_NAND4ABX3 port map( A => n981, B => n982, C => n983, D => 
                           n984, Z => n980);
   U969 : HS65_LH_NAND4ABX3 port map( A => n986, B => n987, C => n988, D => 
                           n989, Z => n979);
   U970 : HS65_LH_OAI21X3 port map( A => n844, B => n6531, C => n2489, Z => 
                           regfile_o(34));
   U971 : HS65_LH_OAI21X3 port map( A => n2490, B => n2491, C => n6530, Z => 
                           n2489);
   U972 : HS65_LH_NAND4ABX3 port map( A => n2492, B => n2493, C => n2494, D => 
                           n2495, Z => n2491);
   U973 : HS65_LH_NAND4ABX3 port map( A => n2497, B => n2498, C => n2499, D => 
                           n2500, Z => n2490);
   U974 : HS65_LH_OAI21X3 port map( A => n842, B => n6531, C => n2433, Z => 
                           regfile_o(36));
   U975 : HS65_LH_OAI21X3 port map( A => n2434, B => n2435, C => n6529, Z => 
                           n2433);
   U976 : HS65_LH_NAND4ABX3 port map( A => n2436, B => n2437, C => n2438, D => 
                           n2439, Z => n2435);
   U977 : HS65_LH_NAND4ABX3 port map( A => n2441, B => n2442, C => n2443, D => 
                           n2444, Z => n2434);
   U978 : HS65_LH_OAI21X3 port map( A => n839, B => n6531, C => n1399, Z => 
                           regfile_o(39));
   U979 : HS65_LH_OAI21X3 port map( A => n1400, B => n1401, C => n6528, Z => 
                           n1399);
   U980 : HS65_LH_NAND4ABX3 port map( A => n1402, B => n1403, C => n1404, D => 
                           n1405, Z => n1401);
   U981 : HS65_LH_NAND4ABX3 port map( A => n1407, B => n1408, C => n1409, D => 
                           n1410, Z => n1400);
   U982 : HS65_LH_OAI21X3 port map( A => n837, B => n6531, C => n1340, Z => 
                           regfile_o(41));
   U983 : HS65_LH_OAI21X3 port map( A => n1341, B => n1342, C => n6528, Z => 
                           n1340);
   U984 : HS65_LH_NAND4ABX3 port map( A => n1343, B => n1344, C => n1345, D => 
                           n1346, Z => n1342);
   U985 : HS65_LH_NAND4ABX3 port map( A => n1363, B => n1364, C => n1365, D => 
                           n1366, Z => n1341);
   U986 : HS65_LH_OAI21X3 port map( A => n824, B => n6531, C => n2601, Z => 
                           regfile_o(54));
   U987 : HS65_LH_OAI21X3 port map( A => n2602, B => n2603, C => n6529, Z => 
                           n2601);
   U988 : HS65_LH_NAND4ABX3 port map( A => n2604, B => n2605, C => n2606, D => 
                           n2607, Z => n2603);
   U989 : HS65_LH_NAND4ABX3 port map( A => n2609, B => n2610, C => n2611, D => 
                           n2612, Z => n2602);
   U990 : HS65_LH_OAI21X3 port map( A => n823, B => n6531, C => n2587, Z => 
                           regfile_o(55));
   U991 : HS65_LH_OAI21X3 port map( A => n2588, B => n2589, C => n6529, Z => 
                           n2587);
   U992 : HS65_LH_NAND4ABX3 port map( A => n2590, B => n2591, C => n2592, D => 
                           n2593, Z => n2589);
   U993 : HS65_LH_NAND4ABX3 port map( A => n2595, B => n2596, C => n2597, D => 
                           n2598, Z => n2588);
   U994 : HS65_LH_OAI21X3 port map( A => n822, B => n6531, C => n2573, Z => 
                           regfile_o(56));
   U995 : HS65_LH_OAI21X3 port map( A => n2574, B => n2575, C => n6530, Z => 
                           n2573);
   U996 : HS65_LH_NAND4ABX3 port map( A => n2576, B => n2577, C => n2578, D => 
                           n2579, Z => n2575);
   U997 : HS65_LH_NAND4ABX3 port map( A => n2581, B => n2582, C => n2583, D => 
                           n2584, Z => n2574);
   U998 : HS65_LH_OAI21X3 port map( A => n821, B => n6531, C => n2559, Z => 
                           regfile_o(57));
   U999 : HS65_LH_OAI21X3 port map( A => n2560, B => n2561, C => n6530, Z => 
                           n2559);
   U1000 : HS65_LH_NAND4ABX3 port map( A => n2562, B => n2563, C => n2564, D =>
                           n2565, Z => n2561);
   U1001 : HS65_LH_NAND4ABX3 port map( A => n2567, B => n2568, C => n2569, D =>
                           n2570, Z => n2560);
   U1002 : HS65_LH_OAI21X3 port map( A => n820, B => n6531, C => n2545, Z => 
                           regfile_o(58));
   U1003 : HS65_LH_OAI21X3 port map( A => n2546, B => n2547, C => n6529, Z => 
                           n2545);
   U1004 : HS65_LH_NAND4ABX3 port map( A => n2548, B => n2549, C => n2550, D =>
                           n2551, Z => n2547);
   U1005 : HS65_LH_NAND4ABX3 port map( A => n2553, B => n2554, C => n2555, D =>
                           n2556, Z => n2546);
   U1006 : HS65_LH_OAI21X3 port map( A => n819, B => n6531, C => n2531, Z => 
                           regfile_o(59));
   U1007 : HS65_LH_OAI21X3 port map( A => n2532, B => n2533, C => n6530, Z => 
                           n2531);
   U1008 : HS65_LH_NAND4ABX3 port map( A => n2534, B => n2535, C => n2536, D =>
                           n2537, Z => n2533);
   U1009 : HS65_LH_NAND4ABX3 port map( A => n2539, B => n2540, C => n2541, D =>
                           n2542, Z => n2532);
   U1010 : HS65_LH_OAI21X3 port map( A => n818, B => n6531, C => n2517, Z => 
                           regfile_o(60));
   U1011 : HS65_LH_OAI21X3 port map( A => n2518, B => n2519, C => n6530, Z => 
                           n2517);
   U1012 : HS65_LH_NAND4ABX3 port map( A => n2520, B => n2521, C => n2522, D =>
                           n2523, Z => n2519);
   U1013 : HS65_LH_NAND4ABX3 port map( A => n2525, B => n2526, C => n2527, D =>
                           n2528, Z => n2518);
   U1014 : HS65_LH_OAI21X3 port map( A => n817, B => n6531, C => n2503, Z => 
                           regfile_o(61));
   U1015 : HS65_LH_OAI21X3 port map( A => n2504, B => n2505, C => n6530, Z => 
                           n2503);
   U1016 : HS65_LH_NAND4ABX3 port map( A => n2506, B => n2507, C => n2508, D =>
                           n2509, Z => n2505);
   U1017 : HS65_LH_NAND4ABX3 port map( A => n2511, B => n2512, C => n2513, D =>
                           n2514, Z => n2504);
   U1018 : HS65_LH_OAI21X3 port map( A => n816, B => n6531, C => n2475, Z => 
                           regfile_o(62));
   U1019 : HS65_LH_OAI21X3 port map( A => n2476, B => n2477, C => n6530, Z => 
                           n2475);
   U1020 : HS65_LH_NAND4ABX3 port map( A => n2478, B => n2479, C => n2480, D =>
                           n2481, Z => n2477);
   U1021 : HS65_LH_NAND4ABX3 port map( A => n2483, B => n2484, C => n2485, D =>
                           n2486, Z => n2476);
   U1022 : HS65_LH_OAI21X3 port map( A => n815, B => n6531, C => n2461, Z => 
                           regfile_o(63));
   U1023 : HS65_LH_OAI21X3 port map( A => n2462, B => n2463, C => n6530, Z => 
                           n2461);
   U1024 : HS65_LH_NAND4ABX3 port map( A => n2464, B => n2465, C => n2466, D =>
                           n2467, Z => n2463);
   U1025 : HS65_LH_NAND4ABX3 port map( A => n2469, B => n2470, C => n2471, D =>
                           n2472, Z => n2462);
   U1026 : HS65_LH_OAI21X3 port map( A => n846, B => n6530, C => n2797, Z => 
                           regfile_o(32));
   U1027 : HS65_LH_OAI21X3 port map( A => n2798, B => n2799, C => n6528, Z => 
                           n2797);
   U1028 : HS65_LH_NAND4ABX3 port map( A => n2800, B => n2801, C => n2802, D =>
                           n2803, Z => n2799);
   U1029 : HS65_LH_NAND4ABX3 port map( A => n2814, B => n2815, C => n2816, D =>
                           n2817, Z => n2798);
   U1030 : HS65_LH_OAI21X3 port map( A => n843, B => n6530, C => n2447, Z => 
                           regfile_o(35));
   U1031 : HS65_LH_OAI21X3 port map( A => n2448, B => n2449, C => n6529, Z => 
                           n2447);
   U1032 : HS65_LH_NAND4ABX3 port map( A => n2450, B => n2451, C => n2452, D =>
                           n2453, Z => n2449);
   U1033 : HS65_LH_NAND4ABX3 port map( A => n2455, B => n2456, C => n2457, D =>
                           n2458, Z => n2448);
   U1034 : HS65_LH_OAI21X3 port map( A => n841, B => n6530, C => n1427, Z => 
                           regfile_o(37));
   U1035 : HS65_LH_OAI21X3 port map( A => n1428, B => n1429, C => n6529, Z => 
                           n1427);
   U1036 : HS65_LH_NAND4ABX3 port map( A => n1430, B => n1431, C => n1432, D =>
                           n1433, Z => n1429);
   U1037 : HS65_LH_NAND4ABX3 port map( A => n2427, B => n2428, C => n2429, D =>
                           n2430, Z => n1428);
   U1038 : HS65_LH_OAI21X3 port map( A => n840, B => n6530, C => n1413, Z => 
                           regfile_o(38));
   U1039 : HS65_LH_OAI21X3 port map( A => n1414, B => n1415, C => n6528, Z => 
                           n1413);
   U1040 : HS65_LH_NAND4ABX3 port map( A => n1416, B => n1417, C => n1418, D =>
                           n1419, Z => n1415);
   U1041 : HS65_LH_NAND4ABX3 port map( A => n1421, B => n1422, C => n1423, D =>
                           n1424, Z => n1414);
   U1042 : HS65_LH_OAI21X3 port map( A => n838, B => n6530, C => n1385, Z => 
                           regfile_o(40));
   U1043 : HS65_LH_OAI21X3 port map( A => n1386, B => n1387, C => n6528, Z => 
                           n1385);
   U1044 : HS65_LH_NAND4ABX3 port map( A => n1388, B => n1389, C => n1390, D =>
                           n1391, Z => n1387);
   U1045 : HS65_LH_NAND4ABX3 port map( A => n1393, B => n1394, C => n1395, D =>
                           n1396, Z => n1386);
   U1046 : HS65_LH_OAI21X3 port map( A => n845, B => n6532, C => n2643, Z => 
                           regfile_o(33));
   U1047 : HS65_LH_OAI21X3 port map( A => n2644, B => n2645, C => n6529, Z => 
                           n2643);
   U1048 : HS65_LH_NAND4ABX3 port map( A => n2646, B => n2647, C => n2648, D =>
                           n2649, Z => n2645);
   U1049 : HS65_LH_NAND4ABX3 port map( A => n2651, B => n2652, C => n2653, D =>
                           n2654, Z => n2644);
   U1050 : HS65_LH_OAI21X3 port map( A => n836, B => n6532, C => n2783, Z => 
                           regfile_o(42));
   U1051 : HS65_LH_OAI21X3 port map( A => n2784, B => n2785, C => n6528, Z => 
                           n2783);
   U1052 : HS65_LH_NAND4ABX3 port map( A => n2786, B => n2787, C => n2788, D =>
                           n2789, Z => n2785);
   U1053 : HS65_LH_NAND4ABX3 port map( A => n2791, B => n2792, C => n2793, D =>
                           n2794, Z => n2784);
   U1054 : HS65_LH_OAI21X3 port map( A => n835, B => n6532, C => n2769, Z => 
                           regfile_o(43));
   U1055 : HS65_LH_OAI21X3 port map( A => n2770, B => n2771, C => n6528, Z => 
                           n2769);
   U1056 : HS65_LH_NAND4ABX3 port map( A => n2772, B => n2773, C => n2774, D =>
                           n2775, Z => n2771);
   U1057 : HS65_LH_NAND4ABX3 port map( A => n2777, B => n2778, C => n2779, D =>
                           n2780, Z => n2770);
   U1058 : HS65_LH_OAI21X3 port map( A => n834, B => n6532, C => n2755, Z => 
                           regfile_o(44));
   U1059 : HS65_LH_OAI21X3 port map( A => n2756, B => n2757, C => n6528, Z => 
                           n2755);
   U1060 : HS65_LH_NAND4ABX3 port map( A => n2758, B => n2759, C => n2760, D =>
                           n2761, Z => n2757);
   U1061 : HS65_LH_NAND4ABX3 port map( A => n2763, B => n2764, C => n2765, D =>
                           n2766, Z => n2756);
   U1062 : HS65_LH_OAI21X3 port map( A => n833, B => n6532, C => n2741, Z => 
                           regfile_o(45));
   U1063 : HS65_LH_OAI21X3 port map( A => n2742, B => n2743, C => n6528, Z => 
                           n2741);
   U1064 : HS65_LH_NAND4ABX3 port map( A => n2744, B => n2745, C => n2746, D =>
                           n2747, Z => n2743);
   U1065 : HS65_LH_NAND4ABX3 port map( A => n2749, B => n2750, C => n2751, D =>
                           n2752, Z => n2742);
   U1066 : HS65_LH_OAI21X3 port map( A => n832, B => n6532, C => n2727, Z => 
                           regfile_o(46));
   U1067 : HS65_LH_OAI21X3 port map( A => n2728, B => n2729, C => n6528, Z => 
                           n2727);
   U1068 : HS65_LH_NAND4ABX3 port map( A => n2730, B => n2731, C => n2732, D =>
                           n2733, Z => n2729);
   U1069 : HS65_LH_NAND4ABX3 port map( A => n2735, B => n2736, C => n2737, D =>
                           n2738, Z => n2728);
   U1070 : HS65_LH_OAI21X3 port map( A => n831, B => n6532, C => n2713, Z => 
                           regfile_o(47));
   U1071 : HS65_LH_OAI21X3 port map( A => n2714, B => n2715, C => n6528, Z => 
                           n2713);
   U1072 : HS65_LH_NAND4ABX3 port map( A => n2716, B => n2717, C => n2718, D =>
                           n2719, Z => n2715);
   U1073 : HS65_LH_NAND4ABX3 port map( A => n2721, B => n2722, C => n2723, D =>
                           n2724, Z => n2714);
   U1074 : HS65_LH_OAI21X3 port map( A => n830, B => n6532, C => n2699, Z => 
                           regfile_o(48));
   U1075 : HS65_LH_OAI21X3 port map( A => n2700, B => n2701, C => n6528, Z => 
                           n2699);
   U1076 : HS65_LH_NAND4ABX3 port map( A => n2702, B => n2703, C => n2704, D =>
                           n2705, Z => n2701);
   U1077 : HS65_LH_NAND4ABX3 port map( A => n2707, B => n2708, C => n2709, D =>
                           n2710, Z => n2700);
   U1078 : HS65_LH_OAI21X3 port map( A => n829, B => n6532, C => n2685, Z => 
                           regfile_o(49));
   U1079 : HS65_LH_OAI21X3 port map( A => n2686, B => n2687, C => n6529, Z => 
                           n2685);
   U1080 : HS65_LH_NAND4ABX3 port map( A => n2688, B => n2689, C => n2690, D =>
                           n2691, Z => n2687);
   U1081 : HS65_LH_NAND4ABX3 port map( A => n2693, B => n2694, C => n2695, D =>
                           n2696, Z => n2686);
   U1082 : HS65_LH_OAI21X3 port map( A => n828, B => n6532, C => n2671, Z => 
                           regfile_o(50));
   U1083 : HS65_LH_OAI21X3 port map( A => n2672, B => n2673, C => n6529, Z => 
                           n2671);
   U1084 : HS65_LH_NAND4ABX3 port map( A => n2674, B => n2675, C => n2676, D =>
                           n2677, Z => n2673);
   U1085 : HS65_LH_NAND4ABX3 port map( A => n2679, B => n2680, C => n2681, D =>
                           n2682, Z => n2672);
   U1086 : HS65_LH_OAI21X3 port map( A => n827, B => n6532, C => n2657, Z => 
                           regfile_o(51));
   U1087 : HS65_LH_OAI21X3 port map( A => n2658, B => n2659, C => n6529, Z => 
                           n2657);
   U1088 : HS65_LH_NAND4ABX3 port map( A => n2660, B => n2661, C => n2662, D =>
                           n2663, Z => n2659);
   U1089 : HS65_LH_NAND4ABX3 port map( A => n2665, B => n2666, C => n2667, D =>
                           n2668, Z => n2658);
   U1090 : HS65_LH_OAI21X3 port map( A => n826, B => n6532, C => n2629, Z => 
                           regfile_o(52));
   U1091 : HS65_LH_OAI21X3 port map( A => n2630, B => n2631, C => n6529, Z => 
                           n2629);
   U1092 : HS65_LH_NAND4ABX3 port map( A => n2632, B => n2633, C => n2634, D =>
                           n2635, Z => n2631);
   U1093 : HS65_LH_NAND4ABX3 port map( A => n2637, B => n2638, C => n2639, D =>
                           n2640, Z => n2630);
   U1094 : HS65_LH_OAI21X3 port map( A => n825, B => n6532, C => n2615, Z => 
                           regfile_o(53));
   U1095 : HS65_LH_OAI21X3 port map( A => n2616, B => n2617, C => n6529, Z => 
                           n2615);
   U1096 : HS65_LH_NAND4ABX3 port map( A => n2618, B => n2619, C => n2620, D =>
                           n2621, Z => n2617);
   U1097 : HS65_LH_NAND4ABX3 port map( A => n2623, B => n2624, C => n2625, D =>
                           n2626, Z => n2616);
   U1098 : HS65_LH_BFX9 port map( A => n6536, Z => n6534);
   U1099 : HS65_LH_BFX9 port map( A => n6536, Z => n6533);
   U1100 : HS65_LH_BFX9 port map( A => n6536, Z => n6535);
   U1101 : HS65_LH_OAI22X6 port map( A => n248, B => n6218, C => n838, D => 
                           n6220, Z => n1666);
   U1102 : HS65_LH_OAI22X6 port map( A => n247, B => n6218, C => n837, D => 
                           n6220, Z => n1667);
   U1103 : HS65_LH_OAI22X6 port map( A => n246, B => n6218, C => n836, D => 
                           n6220, Z => n1668);
   U1104 : HS65_LH_OAI22X6 port map( A => n245, B => n6218, C => n835, D => 
                           n6220, Z => n1669);
   U1105 : HS65_LH_OAI22X6 port map( A => n244, B => n6218, C => n834, D => 
                           n6220, Z => n1670);
   U1106 : HS65_LH_OAI22X6 port map( A => n243, B => n6218, C => n833, D => 
                           n6220, Z => n1671);
   U1107 : HS65_LH_OAI22X6 port map( A => n242, B => n6218, C => n832, D => 
                           n6220, Z => n1672);
   U1108 : HS65_LH_OAI22X6 port map( A => n241, B => n6218, C => n831, D => 
                           n6220, Z => n1673);
   U1109 : HS65_LH_OAI22X6 port map( A => n240, B => n6218, C => n830, D => 
                           n6220, Z => n1674);
   U1110 : HS65_LH_OAI22X6 port map( A => n239, B => n6218, C => n829, D => 
                           n6220, Z => n1675);
   U1111 : HS65_LH_OAI22X6 port map( A => n238, B => n6218, C => n828, D => 
                           n6220, Z => n1676);
   U1112 : HS65_LH_OAI22X6 port map( A => n237, B => n6218, C => n827, D => 
                           n6220, Z => n1677);
   U1113 : HS65_LH_OAI22X6 port map( A => n236, B => n6217, C => n826, D => 
                           n6221, Z => n1678);
   U1114 : HS65_LH_OAI22X6 port map( A => n235, B => n6217, C => n825, D => 
                           n6221, Z => n1679);
   U1115 : HS65_LH_OAI22X6 port map( A => n234, B => n6217, C => n824, D => 
                           n6221, Z => n1680);
   U1116 : HS65_LH_OAI22X6 port map( A => n233, B => n6217, C => n823, D => 
                           n6221, Z => n1681);
   U1117 : HS65_LH_OAI22X6 port map( A => n232, B => n6217, C => n822, D => 
                           n6221, Z => n1682);
   U1118 : HS65_LH_OAI22X6 port map( A => n231, B => n6217, C => n821, D => 
                           n6221, Z => n1683);
   U1119 : HS65_LH_OAI22X6 port map( A => n230, B => n6217, C => n820, D => 
                           n6221, Z => n1684);
   U1120 : HS65_LH_OAI22X6 port map( A => n229, B => n6217, C => n819, D => 
                           n6221, Z => n1685);
   U1121 : HS65_LH_OAI22X6 port map( A => n228, B => n6217, C => n818, D => 
                           n6221, Z => n1686);
   U1122 : HS65_LH_OAI22X6 port map( A => n227, B => n6217, C => n817, D => 
                           n6221, Z => n1687);
   U1123 : HS65_LH_OAI22X6 port map( A => n226, B => n6217, C => n816, D => 
                           n6221, Z => n1688);
   U1124 : HS65_LH_OAI22X6 port map( A => n225, B => n6217, C => n815, D => 
                           n6221, Z => n1689);
   U1125 : HS65_LH_OAI22X6 port map( A => n216, B => n6223, C => n838, D => 
                           n6225, Z => n1698);
   U1126 : HS65_LH_OAI22X6 port map( A => n215, B => n6223, C => n837, D => 
                           n6225, Z => n1699);
   U1127 : HS65_LH_OAI22X6 port map( A => n214, B => n6223, C => n836, D => 
                           n6225, Z => n1700);
   U1128 : HS65_LH_OAI22X6 port map( A => n213, B => n6223, C => n835, D => 
                           n6225, Z => n1701);
   U1129 : HS65_LH_OAI22X6 port map( A => n212, B => n6223, C => n834, D => 
                           n6225, Z => n1702);
   U1130 : HS65_LH_OAI22X6 port map( A => n211, B => n6223, C => n833, D => 
                           n6225, Z => n1703);
   U1131 : HS65_LH_OAI22X6 port map( A => n210, B => n6223, C => n832, D => 
                           n6225, Z => n1704);
   U1132 : HS65_LH_OAI22X6 port map( A => n209, B => n6223, C => n831, D => 
                           n6225, Z => n1705);
   U1133 : HS65_LH_OAI22X6 port map( A => n208, B => n6223, C => n830, D => 
                           n6225, Z => n1706);
   U1134 : HS65_LH_OAI22X6 port map( A => n207, B => n6223, C => n829, D => 
                           n6225, Z => n1707);
   U1135 : HS65_LH_OAI22X6 port map( A => n206, B => n6223, C => n828, D => 
                           n6225, Z => n1708);
   U1136 : HS65_LH_OAI22X6 port map( A => n205, B => n6223, C => n827, D => 
                           n6225, Z => n1709);
   U1137 : HS65_LH_OAI22X6 port map( A => n204, B => n6222, C => n826, D => 
                           n6226, Z => n1710);
   U1138 : HS65_LH_OAI22X6 port map( A => n203, B => n6222, C => n825, D => 
                           n6226, Z => n1711);
   U1139 : HS65_LH_OAI22X6 port map( A => n202, B => n6222, C => n824, D => 
                           n6226, Z => n1712);
   U1140 : HS65_LH_OAI22X6 port map( A => n201, B => n6222, C => n823, D => 
                           n6226, Z => n1713);
   U1141 : HS65_LH_OAI22X6 port map( A => n200, B => n6222, C => n822, D => 
                           n6226, Z => n1714);
   U1142 : HS65_LH_OAI22X6 port map( A => n199, B => n6222, C => n821, D => 
                           n6226, Z => n1715);
   U1143 : HS65_LH_OAI22X6 port map( A => n198, B => n6222, C => n820, D => 
                           n6226, Z => n1716);
   U1144 : HS65_LH_OAI22X6 port map( A => n197, B => n6222, C => n819, D => 
                           n6226, Z => n1717);
   U1145 : HS65_LH_OAI22X6 port map( A => n196, B => n6222, C => n818, D => 
                           n6226, Z => n1718);
   U1146 : HS65_LH_OAI22X6 port map( A => n195, B => n6222, C => n817, D => 
                           n6226, Z => n1719);
   U1147 : HS65_LH_OAI22X6 port map( A => n194, B => n6222, C => n816, D => 
                           n6226, Z => n1720);
   U1148 : HS65_LH_OAI22X6 port map( A => n193, B => n6222, C => n815, D => 
                           n6226, Z => n1721);
   U1149 : HS65_LH_OAI22X6 port map( A => n184, B => n6248, C => n838, D => 
                           n6250, Z => n1858);
   U1150 : HS65_LH_OAI22X6 port map( A => n183, B => n6248, C => n837, D => 
                           n6250, Z => n1859);
   U1151 : HS65_LH_OAI22X6 port map( A => n182, B => n6248, C => n836, D => 
                           n6250, Z => n1860);
   U1152 : HS65_LH_OAI22X6 port map( A => n181, B => n6248, C => n835, D => 
                           n6250, Z => n1861);
   U1153 : HS65_LH_OAI22X6 port map( A => n180, B => n6248, C => n834, D => 
                           n6250, Z => n1862);
   U1154 : HS65_LH_OAI22X6 port map( A => n179, B => n6248, C => n833, D => 
                           n6250, Z => n1863);
   U1155 : HS65_LH_OAI22X6 port map( A => n178, B => n6248, C => n832, D => 
                           n6250, Z => n1864);
   U1156 : HS65_LH_OAI22X6 port map( A => n177, B => n6248, C => n831, D => 
                           n6250, Z => n1865);
   U1157 : HS65_LH_OAI22X6 port map( A => n176, B => n6248, C => n830, D => 
                           n6250, Z => n1866);
   U1158 : HS65_LH_OAI22X6 port map( A => n175, B => n6248, C => n829, D => 
                           n6250, Z => n1867);
   U1159 : HS65_LH_OAI22X6 port map( A => n174, B => n6248, C => n828, D => 
                           n6250, Z => n1868);
   U1160 : HS65_LH_OAI22X6 port map( A => n173, B => n6248, C => n827, D => 
                           n6250, Z => n1869);
   U1161 : HS65_LH_OAI22X6 port map( A => n172, B => n6247, C => n826, D => 
                           n6251, Z => n1870);
   U1162 : HS65_LH_OAI22X6 port map( A => n171, B => n6247, C => n825, D => 
                           n6251, Z => n1871);
   U1163 : HS65_LH_OAI22X6 port map( A => n170, B => n6247, C => n824, D => 
                           n6251, Z => n1872);
   U1164 : HS65_LH_OAI22X6 port map( A => n169, B => n6247, C => n823, D => 
                           n6251, Z => n1873);
   U1165 : HS65_LH_OAI22X6 port map( A => n168, B => n6247, C => n822, D => 
                           n6251, Z => n1874);
   U1166 : HS65_LH_OAI22X6 port map( A => n167, B => n6247, C => n821, D => 
                           n6251, Z => n1875);
   U1167 : HS65_LH_OAI22X6 port map( A => n166, B => n6247, C => n820, D => 
                           n6251, Z => n1876);
   U1168 : HS65_LH_OAI22X6 port map( A => n165, B => n6247, C => n819, D => 
                           n6251, Z => n1877);
   U1169 : HS65_LH_OAI22X6 port map( A => n164, B => n6247, C => n818, D => 
                           n6251, Z => n1878);
   U1170 : HS65_LH_OAI22X6 port map( A => n163, B => n6247, C => n817, D => 
                           n6251, Z => n1879);
   U1171 : HS65_LH_OAI22X6 port map( A => n162, B => n6247, C => n816, D => 
                           n6251, Z => n1880);
   U1172 : HS65_LH_OAI22X6 port map( A => n161, B => n6247, C => n815, D => 
                           n6251, Z => n1881);
   U1173 : HS65_LH_OAI22X6 port map( A => n152, B => n6253, C => n838, D => 
                           n6255, Z => n1890);
   U1174 : HS65_LH_OAI22X6 port map( A => n151, B => n6253, C => n837, D => 
                           n6255, Z => n1891);
   U1175 : HS65_LH_OAI22X6 port map( A => n150, B => n6253, C => n836, D => 
                           n6255, Z => n1892);
   U1176 : HS65_LH_OAI22X6 port map( A => n149, B => n6253, C => n835, D => 
                           n6255, Z => n1893);
   U1177 : HS65_LH_OAI22X6 port map( A => n148, B => n6253, C => n834, D => 
                           n6255, Z => n1894);
   U1178 : HS65_LH_OAI22X6 port map( A => n147, B => n6253, C => n833, D => 
                           n6255, Z => n1895);
   U1179 : HS65_LH_OAI22X6 port map( A => n146, B => n6253, C => n832, D => 
                           n6255, Z => n1896);
   U1180 : HS65_LH_OAI22X6 port map( A => n145, B => n6253, C => n831, D => 
                           n6255, Z => n1897);
   U1181 : HS65_LH_OAI22X6 port map( A => n144, B => n6253, C => n830, D => 
                           n6255, Z => n1898);
   U1182 : HS65_LH_OAI22X6 port map( A => n143, B => n6253, C => n829, D => 
                           n6255, Z => n1899);
   U1183 : HS65_LH_OAI22X6 port map( A => n142, B => n6253, C => n828, D => 
                           n6255, Z => n1900);
   U1184 : HS65_LH_OAI22X6 port map( A => n141, B => n6253, C => n827, D => 
                           n6255, Z => n1901);
   U1185 : HS65_LH_OAI22X6 port map( A => n140, B => n6252, C => n826, D => 
                           n6256, Z => n1902);
   U1186 : HS65_LH_OAI22X6 port map( A => n139, B => n6252, C => n825, D => 
                           n6256, Z => n1903);
   U1187 : HS65_LH_OAI22X6 port map( A => n138, B => n6252, C => n824, D => 
                           n6256, Z => n1904);
   U1188 : HS65_LH_OAI22X6 port map( A => n137, B => n6252, C => n823, D => 
                           n6256, Z => n1905);
   U1189 : HS65_LH_OAI22X6 port map( A => n136, B => n6252, C => n822, D => 
                           n6256, Z => n1906);
   U1190 : HS65_LH_OAI22X6 port map( A => n135, B => n6252, C => n821, D => 
                           n6256, Z => n1907);
   U1191 : HS65_LH_OAI22X6 port map( A => n134, B => n6252, C => n820, D => 
                           n6256, Z => n1908);
   U1192 : HS65_LH_OAI22X6 port map( A => n133, B => n6252, C => n819, D => 
                           n6256, Z => n1909);
   U1193 : HS65_LH_OAI22X6 port map( A => n132, B => n6252, C => n818, D => 
                           n6256, Z => n1910);
   U1194 : HS65_LH_OAI22X6 port map( A => n131, B => n6252, C => n817, D => 
                           n6256, Z => n1911);
   U1195 : HS65_LH_OAI22X6 port map( A => n130, B => n6252, C => n816, D => 
                           n6256, Z => n1912);
   U1196 : HS65_LH_OAI22X6 port map( A => n129, B => n6252, C => n815, D => 
                           n6256, Z => n1913);
   U1197 : HS65_LH_OAI22X6 port map( A => n24, B => n6323, C => n838, D => 
                           n6325, Z => n2338);
   U1198 : HS65_LH_OAI22X6 port map( A => n23, B => n6323, C => n837, D => 
                           n6325, Z => n2339);
   U1199 : HS65_LH_OAI22X6 port map( A => n22, B => n6323, C => n836, D => 
                           n6325, Z => n2340);
   U1200 : HS65_LH_OAI22X6 port map( A => n21, B => n6323, C => n835, D => 
                           n6325, Z => n2341);
   U1201 : HS65_LH_OAI22X6 port map( A => n20, B => n6323, C => n834, D => 
                           n6325, Z => n2342);
   U1202 : HS65_LH_OAI22X6 port map( A => n19, B => n6323, C => n833, D => 
                           n6325, Z => n2343);
   U1203 : HS65_LH_OAI22X6 port map( A => n18, B => n6323, C => n832, D => 
                           n6325, Z => n2344);
   U1204 : HS65_LH_OAI22X6 port map( A => n17, B => n6323, C => n831, D => 
                           n6325, Z => n2345);
   U1205 : HS65_LH_OAI22X6 port map( A => n16, B => n6323, C => n830, D => 
                           n6325, Z => n2346);
   U1206 : HS65_LH_OAI22X6 port map( A => n15, B => n6323, C => n829, D => 
                           n6325, Z => n2347);
   U1207 : HS65_LH_OAI22X6 port map( A => n14, B => n6323, C => n828, D => 
                           n6325, Z => n2348);
   U1208 : HS65_LH_OAI22X6 port map( A => n13, B => n6323, C => n827, D => 
                           n6325, Z => n2349);
   U1209 : HS65_LH_OAI22X6 port map( A => n12, B => n6322, C => n826, D => 
                           n6326, Z => n2350);
   U1210 : HS65_LH_OAI22X6 port map( A => n11, B => n6322, C => n825, D => 
                           n6326, Z => n2351);
   U1211 : HS65_LH_OAI22X6 port map( A => n10, B => n6322, C => n824, D => 
                           n6326, Z => n2352);
   U1212 : HS65_LH_OAI22X6 port map( A => n9, B => n6322, C => n823, D => n6326
                           , Z => n2353);
   U1213 : HS65_LH_OAI22X6 port map( A => n8, B => n6322, C => n822, D => n6326
                           , Z => n2354);
   U1214 : HS65_LH_OAI22X6 port map( A => n7, B => n6322, C => n821, D => n6326
                           , Z => n2355);
   U1215 : HS65_LH_OAI22X6 port map( A => n6, B => n6322, C => n820, D => n6326
                           , Z => n2356);
   U1216 : HS65_LH_OAI22X6 port map( A => n5, B => n6322, C => n819, D => n6326
                           , Z => n2357);
   U1217 : HS65_LH_OAI22X6 port map( A => n4, B => n6322, C => n818, D => n6326
                           , Z => n2358);
   U1218 : HS65_LH_OAI22X6 port map( A => n3, B => n6322, C => n817, D => n6326
                           , Z => n2359);
   U1219 : HS65_LH_OAI22X6 port map( A => n2, B => n6322, C => n816, D => n6326
                           , Z => n2360);
   U1220 : HS65_LH_OAI22X6 port map( A => n1, B => n6322, C => n815, D => n6326
                           , Z => n2361);
   U1221 : HS65_LH_OAI22X6 port map( A => n120, B => n6308, C => n838, D => 
                           n6310, Z => n2242);
   U1222 : HS65_LH_OAI22X6 port map( A => n119, B => n6308, C => n837, D => 
                           n6310, Z => n2243);
   U1223 : HS65_LH_OAI22X6 port map( A => n118, B => n6308, C => n836, D => 
                           n6310, Z => n2244);
   U1224 : HS65_LH_OAI22X6 port map( A => n117, B => n6308, C => n835, D => 
                           n6310, Z => n2245);
   U1225 : HS65_LH_OAI22X6 port map( A => n116, B => n6308, C => n834, D => 
                           n6310, Z => n2246);
   U1226 : HS65_LH_OAI22X6 port map( A => n115, B => n6308, C => n833, D => 
                           n6310, Z => n2247);
   U1227 : HS65_LH_OAI22X6 port map( A => n114, B => n6308, C => n832, D => 
                           n6310, Z => n2248);
   U1228 : HS65_LH_OAI22X6 port map( A => n113, B => n6308, C => n831, D => 
                           n6310, Z => n2249);
   U1229 : HS65_LH_OAI22X6 port map( A => n112, B => n6308, C => n830, D => 
                           n6310, Z => n2250);
   U1230 : HS65_LH_OAI22X6 port map( A => n111, B => n6308, C => n829, D => 
                           n6310, Z => n2251);
   U1231 : HS65_LH_OAI22X6 port map( A => n110, B => n6308, C => n828, D => 
                           n6310, Z => n2252);
   U1232 : HS65_LH_OAI22X6 port map( A => n109, B => n6308, C => n827, D => 
                           n6310, Z => n2253);
   U1233 : HS65_LH_OAI22X6 port map( A => n108, B => n6307, C => n826, D => 
                           n6311, Z => n2254);
   U1234 : HS65_LH_OAI22X6 port map( A => n107, B => n6307, C => n825, D => 
                           n6311, Z => n2255);
   U1235 : HS65_LH_OAI22X6 port map( A => n106, B => n6307, C => n824, D => 
                           n6311, Z => n2256);
   U1236 : HS65_LH_OAI22X6 port map( A => n105, B => n6307, C => n823, D => 
                           n6311, Z => n2257);
   U1237 : HS65_LH_OAI22X6 port map( A => n104, B => n6307, C => n822, D => 
                           n6311, Z => n2258);
   U1238 : HS65_LH_OAI22X6 port map( A => n103, B => n6307, C => n821, D => 
                           n6311, Z => n2259);
   U1239 : HS65_LH_OAI22X6 port map( A => n102, B => n6307, C => n820, D => 
                           n6311, Z => n2260);
   U1240 : HS65_LH_OAI22X6 port map( A => n101, B => n6307, C => n819, D => 
                           n6311, Z => n2261);
   U1241 : HS65_LH_OAI22X6 port map( A => n100, B => n6307, C => n818, D => 
                           n6311, Z => n2262);
   U1242 : HS65_LH_OAI22X6 port map( A => n99, B => n6307, C => n817, D => 
                           n6311, Z => n2263);
   U1243 : HS65_LH_OAI22X6 port map( A => n98, B => n6307, C => n816, D => 
                           n6311, Z => n2264);
   U1244 : HS65_LH_OAI22X6 port map( A => n97, B => n6307, C => n815, D => 
                           n6311, Z => n2265);
   U1245 : HS65_LH_OAI22X6 port map( A => n56, B => n6318, C => n838, D => 
                           n6320, Z => n2306);
   U1246 : HS65_LH_OAI22X6 port map( A => n55, B => n6318, C => n837, D => 
                           n6320, Z => n2307);
   U1247 : HS65_LH_OAI22X6 port map( A => n54, B => n6318, C => n836, D => 
                           n6320, Z => n2308);
   U1248 : HS65_LH_OAI22X6 port map( A => n53, B => n6318, C => n835, D => 
                           n6320, Z => n2309);
   U1249 : HS65_LH_OAI22X6 port map( A => n52, B => n6318, C => n834, D => 
                           n6320, Z => n2310);
   U1250 : HS65_LH_OAI22X6 port map( A => n51, B => n6318, C => n833, D => 
                           n6320, Z => n2311);
   U1251 : HS65_LH_OAI22X6 port map( A => n50, B => n6318, C => n832, D => 
                           n6320, Z => n2312);
   U1252 : HS65_LH_OAI22X6 port map( A => n49, B => n6318, C => n831, D => 
                           n6320, Z => n2313);
   U1253 : HS65_LH_OAI22X6 port map( A => n48, B => n6318, C => n830, D => 
                           n6320, Z => n2314);
   U1254 : HS65_LH_OAI22X6 port map( A => n47, B => n6318, C => n829, D => 
                           n6320, Z => n2315);
   U1255 : HS65_LH_OAI22X6 port map( A => n46, B => n6318, C => n828, D => 
                           n6320, Z => n2316);
   U1256 : HS65_LH_OAI22X6 port map( A => n45, B => n6318, C => n827, D => 
                           n6320, Z => n2317);
   U1257 : HS65_LH_OAI22X6 port map( A => n44, B => n6317, C => n826, D => 
                           n6321, Z => n2318);
   U1258 : HS65_LH_OAI22X6 port map( A => n43, B => n6317, C => n825, D => 
                           n6321, Z => n2319);
   U1259 : HS65_LH_OAI22X6 port map( A => n42, B => n6317, C => n824, D => 
                           n6321, Z => n2320);
   U1260 : HS65_LH_OAI22X6 port map( A => n41, B => n6317, C => n823, D => 
                           n6321, Z => n2321);
   U1261 : HS65_LH_OAI22X6 port map( A => n40, B => n6317, C => n822, D => 
                           n6321, Z => n2322);
   U1262 : HS65_LH_OAI22X6 port map( A => n39, B => n6317, C => n821, D => 
                           n6321, Z => n2323);
   U1263 : HS65_LH_OAI22X6 port map( A => n38, B => n6317, C => n820, D => 
                           n6321, Z => n2324);
   U1264 : HS65_LH_OAI22X6 port map( A => n37, B => n6317, C => n819, D => 
                           n6321, Z => n2325);
   U1265 : HS65_LH_OAI22X6 port map( A => n36, B => n6317, C => n818, D => 
                           n6321, Z => n2326);
   U1266 : HS65_LH_OAI22X6 port map( A => n35, B => n6317, C => n817, D => 
                           n6321, Z => n2327);
   U1267 : HS65_LH_OAI22X6 port map( A => n34, B => n6317, C => n816, D => 
                           n6321, Z => n2328);
   U1268 : HS65_LH_OAI22X6 port map( A => n33, B => n6317, C => n815, D => 
                           n6321, Z => n2329);
   U1269 : HS65_LH_OAI22X6 port map( A => n88, B => n6313, C => n838, D => 
                           n6315, Z => n2274);
   U1270 : HS65_LH_OAI22X6 port map( A => n87, B => n6313, C => n837, D => 
                           n6315, Z => n2275);
   U1271 : HS65_LH_OAI22X6 port map( A => n86, B => n6313, C => n836, D => 
                           n6315, Z => n2276);
   U1272 : HS65_LH_OAI22X6 port map( A => n85, B => n6313, C => n835, D => 
                           n6315, Z => n2277);
   U1273 : HS65_LH_OAI22X6 port map( A => n84, B => n6313, C => n834, D => 
                           n6315, Z => n2278);
   U1274 : HS65_LH_OAI22X6 port map( A => n83, B => n6313, C => n833, D => 
                           n6315, Z => n2279);
   U1275 : HS65_LH_OAI22X6 port map( A => n82, B => n6313, C => n832, D => 
                           n6315, Z => n2280);
   U1276 : HS65_LH_OAI22X6 port map( A => n81, B => n6313, C => n831, D => 
                           n6315, Z => n2281);
   U1277 : HS65_LH_OAI22X6 port map( A => n80, B => n6313, C => n830, D => 
                           n6315, Z => n2282);
   U1278 : HS65_LH_OAI22X6 port map( A => n79, B => n6313, C => n829, D => 
                           n6315, Z => n2283);
   U1279 : HS65_LH_OAI22X6 port map( A => n78, B => n6313, C => n828, D => 
                           n6315, Z => n2284);
   U1280 : HS65_LH_OAI22X6 port map( A => n77, B => n6313, C => n827, D => 
                           n6315, Z => n2285);
   U1281 : HS65_LH_OAI22X6 port map( A => n76, B => n6312, C => n826, D => 
                           n6316, Z => n2286);
   U1282 : HS65_LH_OAI22X6 port map( A => n75, B => n6312, C => n825, D => 
                           n6316, Z => n2287);
   U1283 : HS65_LH_OAI22X6 port map( A => n74, B => n6312, C => n824, D => 
                           n6316, Z => n2288);
   U1284 : HS65_LH_OAI22X6 port map( A => n73, B => n6312, C => n823, D => 
                           n6316, Z => n2289);
   U1285 : HS65_LH_OAI22X6 port map( A => n72, B => n6312, C => n822, D => 
                           n6316, Z => n2290);
   U1286 : HS65_LH_OAI22X6 port map( A => n71, B => n6312, C => n821, D => 
                           n6316, Z => n2291);
   U1287 : HS65_LH_OAI22X6 port map( A => n70, B => n6312, C => n820, D => 
                           n6316, Z => n2292);
   U1288 : HS65_LH_OAI22X6 port map( A => n69, B => n6312, C => n819, D => 
                           n6316, Z => n2293);
   U1289 : HS65_LH_OAI22X6 port map( A => n68, B => n6312, C => n818, D => 
                           n6316, Z => n2294);
   U1290 : HS65_LH_OAI22X6 port map( A => n67, B => n6312, C => n817, D => 
                           n6316, Z => n2295);
   U1291 : HS65_LH_OAI22X6 port map( A => n66, B => n6312, C => n816, D => 
                           n6316, Z => n2296);
   U1292 : HS65_LH_OAI22X6 port map( A => n65, B => n6312, C => n815, D => 
                           n6316, Z => n2297);
   U1293 : HS65_LH_OAI22X6 port map( A => n256, B => n6218, C => n846, D => 
                           n6219, Z => n1658);
   U1294 : HS65_LH_OAI22X6 port map( A => n255, B => n6217, C => n845, D => 
                           n6220, Z => n1659);
   U1295 : HS65_LH_OAI22X6 port map( A => n254, B => n6218, C => n844, D => 
                           n6220, Z => n1660);
   U1296 : HS65_LH_OAI22X6 port map( A => n253, B => n6217, C => n843, D => 
                           n6220, Z => n1661);
   U1297 : HS65_LH_OAI22X6 port map( A => n252, B => n6218, C => n842, D => 
                           n6220, Z => n1662);
   U1298 : HS65_LH_OAI22X6 port map( A => n251, B => n6217, C => n841, D => 
                           n6220, Z => n1663);
   U1299 : HS65_LH_OAI22X6 port map( A => n250, B => n6218, C => n840, D => 
                           n6220, Z => n1664);
   U1300 : HS65_LH_OAI22X6 port map( A => n249, B => n6217, C => n839, D => 
                           n6220, Z => n1665);
   U1301 : HS65_LH_OAI22X6 port map( A => n224, B => n6223, C => n846, D => 
                           n6224, Z => n1690);
   U1302 : HS65_LH_OAI22X6 port map( A => n223, B => n6222, C => n845, D => 
                           n6225, Z => n1691);
   U1303 : HS65_LH_OAI22X6 port map( A => n222, B => n6223, C => n844, D => 
                           n6225, Z => n1692);
   U1304 : HS65_LH_OAI22X6 port map( A => n221, B => n6222, C => n843, D => 
                           n6225, Z => n1693);
   U1305 : HS65_LH_OAI22X6 port map( A => n220, B => n6223, C => n842, D => 
                           n6225, Z => n1694);
   U1306 : HS65_LH_OAI22X6 port map( A => n219, B => n6222, C => n841, D => 
                           n6225, Z => n1695);
   U1307 : HS65_LH_OAI22X6 port map( A => n218, B => n6223, C => n840, D => 
                           n6225, Z => n1696);
   U1308 : HS65_LH_OAI22X6 port map( A => n217, B => n6222, C => n839, D => 
                           n6225, Z => n1697);
   U1309 : HS65_LH_OAI22X6 port map( A => n192, B => n6248, C => n846, D => 
                           n6249, Z => n1850);
   U1310 : HS65_LH_OAI22X6 port map( A => n191, B => n6247, C => n845, D => 
                           n6250, Z => n1851);
   U1311 : HS65_LH_OAI22X6 port map( A => n190, B => n6248, C => n844, D => 
                           n6250, Z => n1852);
   U1312 : HS65_LH_OAI22X6 port map( A => n189, B => n6247, C => n843, D => 
                           n6250, Z => n1853);
   U1313 : HS65_LH_OAI22X6 port map( A => n188, B => n6248, C => n842, D => 
                           n6250, Z => n1854);
   U1314 : HS65_LH_OAI22X6 port map( A => n187, B => n6247, C => n841, D => 
                           n6250, Z => n1855);
   U1315 : HS65_LH_OAI22X6 port map( A => n186, B => n6248, C => n840, D => 
                           n6250, Z => n1856);
   U1316 : HS65_LH_OAI22X6 port map( A => n185, B => n6247, C => n839, D => 
                           n6250, Z => n1857);
   U1317 : HS65_LH_OAI22X6 port map( A => n160, B => n6253, C => n846, D => 
                           n6254, Z => n1882);
   U1318 : HS65_LH_OAI22X6 port map( A => n159, B => n6252, C => n845, D => 
                           n6255, Z => n1883);
   U1319 : HS65_LH_OAI22X6 port map( A => n158, B => n6253, C => n844, D => 
                           n6255, Z => n1884);
   U1320 : HS65_LH_OAI22X6 port map( A => n157, B => n6252, C => n843, D => 
                           n6255, Z => n1885);
   U1321 : HS65_LH_OAI22X6 port map( A => n156, B => n6253, C => n842, D => 
                           n6255, Z => n1886);
   U1322 : HS65_LH_OAI22X6 port map( A => n155, B => n6252, C => n841, D => 
                           n6255, Z => n1887);
   U1323 : HS65_LH_OAI22X6 port map( A => n154, B => n6253, C => n840, D => 
                           n6255, Z => n1888);
   U1324 : HS65_LH_OAI22X6 port map( A => n153, B => n6252, C => n839, D => 
                           n6255, Z => n1889);
   U1325 : HS65_LH_OAI22X6 port map( A => n32, B => n6323, C => n846, D => 
                           n6324, Z => n2330);
   U1326 : HS65_LH_OAI22X6 port map( A => n31, B => n6322, C => n845, D => 
                           n6325, Z => n2331);
   U1327 : HS65_LH_OAI22X6 port map( A => n30, B => n6323, C => n844, D => 
                           n6325, Z => n2332);
   U1328 : HS65_LH_OAI22X6 port map( A => n29, B => n6322, C => n843, D => 
                           n6325, Z => n2333);
   U1329 : HS65_LH_OAI22X6 port map( A => n28, B => n6323, C => n842, D => 
                           n6325, Z => n2334);
   U1330 : HS65_LH_OAI22X6 port map( A => n27, B => n6322, C => n841, D => 
                           n6325, Z => n2335);
   U1331 : HS65_LH_OAI22X6 port map( A => n26, B => n6323, C => n840, D => 
                           n6325, Z => n2336);
   U1332 : HS65_LH_OAI22X6 port map( A => n25, B => n6322, C => n839, D => 
                           n6325, Z => n2337);
   U1333 : HS65_LH_OAI22X6 port map( A => n128, B => n6308, C => n846, D => 
                           n6309, Z => n2234);
   U1334 : HS65_LH_OAI22X6 port map( A => n127, B => n6307, C => n845, D => 
                           n6310, Z => n2235);
   U1335 : HS65_LH_OAI22X6 port map( A => n126, B => n6308, C => n844, D => 
                           n6310, Z => n2236);
   U1336 : HS65_LH_OAI22X6 port map( A => n125, B => n6307, C => n843, D => 
                           n6310, Z => n2237);
   U1337 : HS65_LH_OAI22X6 port map( A => n124, B => n6308, C => n842, D => 
                           n6310, Z => n2238);
   U1338 : HS65_LH_OAI22X6 port map( A => n123, B => n6307, C => n841, D => 
                           n6310, Z => n2239);
   U1339 : HS65_LH_OAI22X6 port map( A => n122, B => n6308, C => n840, D => 
                           n6310, Z => n2240);
   U1340 : HS65_LH_OAI22X6 port map( A => n121, B => n6307, C => n839, D => 
                           n6310, Z => n2241);
   U1341 : HS65_LH_OAI22X6 port map( A => n64, B => n6318, C => n846, D => 
                           n6319, Z => n2298);
   U1342 : HS65_LH_OAI22X6 port map( A => n63, B => n6317, C => n845, D => 
                           n6320, Z => n2299);
   U1343 : HS65_LH_OAI22X6 port map( A => n62, B => n6318, C => n844, D => 
                           n6320, Z => n2300);
   U1344 : HS65_LH_OAI22X6 port map( A => n61, B => n6317, C => n843, D => 
                           n6320, Z => n2301);
   U1345 : HS65_LH_OAI22X6 port map( A => n60, B => n6318, C => n842, D => 
                           n6320, Z => n2302);
   U1346 : HS65_LH_OAI22X6 port map( A => n59, B => n6317, C => n841, D => 
                           n6320, Z => n2303);
   U1347 : HS65_LH_OAI22X6 port map( A => n58, B => n6318, C => n840, D => 
                           n6320, Z => n2304);
   U1348 : HS65_LH_OAI22X6 port map( A => n57, B => n6317, C => n839, D => 
                           n6320, Z => n2305);
   U1349 : HS65_LH_OAI22X6 port map( A => n96, B => n6313, C => n846, D => 
                           n6314, Z => n2266);
   U1350 : HS65_LH_OAI22X6 port map( A => n95, B => n6312, C => n845, D => 
                           n6315, Z => n2267);
   U1351 : HS65_LH_OAI22X6 port map( A => n94, B => n6313, C => n844, D => 
                           n6315, Z => n2268);
   U1352 : HS65_LH_OAI22X6 port map( A => n93, B => n6312, C => n843, D => 
                           n6315, Z => n2269);
   U1353 : HS65_LH_OAI22X6 port map( A => n92, B => n6313, C => n842, D => 
                           n6315, Z => n2270);
   U1354 : HS65_LH_OAI22X6 port map( A => n91, B => n6312, C => n841, D => 
                           n6315, Z => n2271);
   U1355 : HS65_LH_OAI22X6 port map( A => n90, B => n6313, C => n840, D => 
                           n6315, Z => n2272);
   U1356 : HS65_LH_OAI22X6 port map( A => n89, B => n6312, C => n839, D => 
                           n6315, Z => n2273);
   U1357 : HS65_LH_IVX9 port map( A => registers_25_0_port, Z => n288);
   U1358 : HS65_LH_IVX9 port map( A => registers_25_1_port, Z => n287);
   U1359 : HS65_LH_IVX9 port map( A => registers_25_2_port, Z => n286);
   U1360 : HS65_LH_IVX9 port map( A => registers_25_3_port, Z => n285);
   U1361 : HS65_LH_IVX9 port map( A => registers_25_4_port, Z => n284);
   U1362 : HS65_LH_IVX9 port map( A => registers_25_5_port, Z => n283);
   U1363 : HS65_LH_IVX9 port map( A => registers_25_6_port, Z => n282);
   U1364 : HS65_LH_IVX9 port map( A => registers_25_7_port, Z => n281);
   U1365 : HS65_LH_IVX9 port map( A => registers_25_8_port, Z => n280);
   U1366 : HS65_LH_IVX9 port map( A => registers_25_9_port, Z => n279);
   U1367 : HS65_LH_IVX9 port map( A => registers_25_10_port, Z => n278);
   U1368 : HS65_LH_IVX9 port map( A => registers_25_11_port, Z => n277);
   U1369 : HS65_LH_IVX9 port map( A => registers_25_12_port, Z => n276);
   U1370 : HS65_LH_IVX9 port map( A => registers_25_13_port, Z => n275);
   U1371 : HS65_LH_IVX9 port map( A => registers_25_14_port, Z => n274);
   U1372 : HS65_LH_IVX9 port map( A => registers_25_15_port, Z => n273);
   U1373 : HS65_LH_IVX9 port map( A => registers_25_16_port, Z => n272);
   U1374 : HS65_LH_IVX9 port map( A => registers_25_17_port, Z => n271);
   U1375 : HS65_LH_IVX9 port map( A => registers_25_18_port, Z => n270);
   U1376 : HS65_LH_IVX9 port map( A => registers_25_19_port, Z => n269);
   U1377 : HS65_LH_IVX9 port map( A => registers_25_20_port, Z => n268);
   U1378 : HS65_LH_IVX9 port map( A => registers_25_21_port, Z => n267);
   U1379 : HS65_LH_IVX9 port map( A => registers_25_22_port, Z => n266);
   U1380 : HS65_LH_IVX9 port map( A => registers_25_23_port, Z => n265);
   U1381 : HS65_LH_IVX9 port map( A => registers_25_24_port, Z => n264);
   U1382 : HS65_LH_IVX9 port map( A => registers_25_25_port, Z => n263);
   U1383 : HS65_LH_IVX9 port map( A => registers_25_26_port, Z => n262);
   U1384 : HS65_LH_IVX9 port map( A => registers_25_27_port, Z => n261);
   U1385 : HS65_LH_IVX9 port map( A => registers_25_28_port, Z => n260);
   U1386 : HS65_LH_IVX9 port map( A => registers_25_29_port, Z => n259);
   U1387 : HS65_LH_IVX9 port map( A => registers_25_30_port, Z => n258);
   U1388 : HS65_LH_IVX9 port map( A => registers_25_31_port, Z => n257);
   U1389 : HS65_LH_IVX9 port map( A => registers_16_0_port, Z => n416);
   U1390 : HS65_LH_IVX9 port map( A => registers_16_1_port, Z => n415);
   U1391 : HS65_LH_IVX9 port map( A => registers_16_2_port, Z => n414);
   U1392 : HS65_LH_IVX9 port map( A => registers_16_3_port, Z => n413);
   U1393 : HS65_LH_IVX9 port map( A => registers_16_4_port, Z => n412);
   U1394 : HS65_LH_IVX9 port map( A => registers_16_5_port, Z => n411);
   U1395 : HS65_LH_IVX9 port map( A => registers_16_6_port, Z => n410);
   U1396 : HS65_LH_IVX9 port map( A => registers_16_7_port, Z => n409);
   U1397 : HS65_LH_IVX9 port map( A => registers_16_8_port, Z => n408);
   U1398 : HS65_LH_IVX9 port map( A => registers_16_9_port, Z => n407);
   U1399 : HS65_LH_IVX9 port map( A => registers_16_10_port, Z => n406);
   U1400 : HS65_LH_IVX9 port map( A => registers_16_11_port, Z => n405);
   U1401 : HS65_LH_IVX9 port map( A => registers_16_12_port, Z => n404);
   U1402 : HS65_LH_IVX9 port map( A => registers_16_13_port, Z => n403);
   U1403 : HS65_LH_IVX9 port map( A => registers_16_14_port, Z => n402);
   U1404 : HS65_LH_IVX9 port map( A => registers_16_15_port, Z => n401);
   U1405 : HS65_LH_IVX9 port map( A => registers_16_16_port, Z => n400);
   U1406 : HS65_LH_IVX9 port map( A => registers_16_17_port, Z => n399);
   U1407 : HS65_LH_IVX9 port map( A => registers_16_18_port, Z => n398);
   U1408 : HS65_LH_IVX9 port map( A => registers_16_19_port, Z => n397);
   U1409 : HS65_LH_IVX9 port map( A => registers_16_20_port, Z => n396);
   U1410 : HS65_LH_IVX9 port map( A => registers_16_21_port, Z => n395);
   U1411 : HS65_LH_IVX9 port map( A => registers_16_22_port, Z => n394);
   U1412 : HS65_LH_IVX9 port map( A => registers_16_23_port, Z => n393);
   U1413 : HS65_LH_IVX9 port map( A => registers_16_24_port, Z => n392);
   U1414 : HS65_LH_IVX9 port map( A => registers_16_25_port, Z => n391);
   U1415 : HS65_LH_IVX9 port map( A => registers_16_26_port, Z => n390);
   U1416 : HS65_LH_IVX9 port map( A => registers_16_27_port, Z => n389);
   U1417 : HS65_LH_IVX9 port map( A => registers_16_28_port, Z => n388);
   U1418 : HS65_LH_IVX9 port map( A => registers_16_29_port, Z => n387);
   U1419 : HS65_LH_IVX9 port map( A => registers_16_30_port, Z => n386);
   U1420 : HS65_LH_IVX9 port map( A => registers_16_31_port, Z => n385);
   U1421 : HS65_LH_IVX9 port map( A => registers_10_0_port, Z => n480);
   U1422 : HS65_LH_IVX9 port map( A => registers_10_1_port, Z => n479);
   U1423 : HS65_LH_IVX9 port map( A => registers_10_2_port, Z => n478);
   U1424 : HS65_LH_IVX9 port map( A => registers_10_3_port, Z => n477);
   U1425 : HS65_LH_IVX9 port map( A => registers_10_4_port, Z => n476);
   U1426 : HS65_LH_IVX9 port map( A => registers_10_5_port, Z => n475);
   U1427 : HS65_LH_IVX9 port map( A => registers_10_6_port, Z => n474);
   U1428 : HS65_LH_IVX9 port map( A => registers_10_7_port, Z => n473);
   U1429 : HS65_LH_IVX9 port map( A => registers_10_8_port, Z => n472);
   U1430 : HS65_LH_IVX9 port map( A => registers_10_9_port, Z => n471);
   U1431 : HS65_LH_IVX9 port map( A => registers_10_10_port, Z => n470);
   U1432 : HS65_LH_IVX9 port map( A => registers_10_11_port, Z => n469);
   U1433 : HS65_LH_IVX9 port map( A => registers_10_12_port, Z => n468);
   U1434 : HS65_LH_IVX9 port map( A => registers_10_13_port, Z => n467);
   U1435 : HS65_LH_IVX9 port map( A => registers_10_14_port, Z => n466);
   U1436 : HS65_LH_IVX9 port map( A => registers_10_15_port, Z => n465);
   U1437 : HS65_LH_IVX9 port map( A => registers_10_16_port, Z => n464);
   U1438 : HS65_LH_IVX9 port map( A => registers_10_17_port, Z => n463);
   U1439 : HS65_LH_IVX9 port map( A => registers_10_18_port, Z => n462);
   U1440 : HS65_LH_IVX9 port map( A => registers_10_19_port, Z => n461);
   U1441 : HS65_LH_IVX9 port map( A => registers_10_20_port, Z => n460);
   U1442 : HS65_LH_IVX9 port map( A => registers_10_21_port, Z => n459);
   U1443 : HS65_LH_IVX9 port map( A => registers_10_22_port, Z => n458);
   U1444 : HS65_LH_IVX9 port map( A => registers_10_23_port, Z => n457);
   U1445 : HS65_LH_IVX9 port map( A => registers_10_24_port, Z => n456);
   U1446 : HS65_LH_IVX9 port map( A => registers_10_25_port, Z => n455);
   U1447 : HS65_LH_IVX9 port map( A => registers_10_26_port, Z => n454);
   U1448 : HS65_LH_IVX9 port map( A => registers_10_27_port, Z => n453);
   U1449 : HS65_LH_IVX9 port map( A => registers_10_28_port, Z => n452);
   U1450 : HS65_LH_IVX9 port map( A => registers_10_29_port, Z => n451);
   U1451 : HS65_LH_IVX9 port map( A => registers_10_30_port, Z => n450);
   U1452 : HS65_LH_IVX9 port map( A => registers_10_31_port, Z => n449);
   U1453 : HS65_LH_IVX9 port map( A => registers_18_0_port, Z => n352);
   U1454 : HS65_LH_IVX9 port map( A => registers_18_1_port, Z => n351);
   U1455 : HS65_LH_IVX9 port map( A => registers_18_2_port, Z => n350);
   U1456 : HS65_LH_IVX9 port map( A => registers_18_3_port, Z => n349);
   U1457 : HS65_LH_IVX9 port map( A => registers_18_4_port, Z => n348);
   U1458 : HS65_LH_IVX9 port map( A => registers_18_5_port, Z => n347);
   U1459 : HS65_LH_IVX9 port map( A => registers_18_6_port, Z => n346);
   U1460 : HS65_LH_IVX9 port map( A => registers_18_7_port, Z => n345);
   U1461 : HS65_LH_IVX9 port map( A => registers_18_8_port, Z => n344);
   U1462 : HS65_LH_IVX9 port map( A => registers_18_9_port, Z => n343);
   U1463 : HS65_LH_IVX9 port map( A => registers_18_10_port, Z => n342);
   U1464 : HS65_LH_IVX9 port map( A => registers_18_11_port, Z => n341);
   U1465 : HS65_LH_IVX9 port map( A => registers_18_12_port, Z => n340);
   U1466 : HS65_LH_IVX9 port map( A => registers_18_13_port, Z => n339);
   U1467 : HS65_LH_IVX9 port map( A => registers_18_14_port, Z => n338);
   U1468 : HS65_LH_IVX9 port map( A => registers_18_15_port, Z => n337);
   U1469 : HS65_LH_IVX9 port map( A => registers_18_16_port, Z => n336);
   U1470 : HS65_LH_IVX9 port map( A => registers_18_17_port, Z => n335);
   U1471 : HS65_LH_IVX9 port map( A => registers_18_18_port, Z => n334);
   U1472 : HS65_LH_IVX9 port map( A => registers_18_19_port, Z => n333);
   U1473 : HS65_LH_IVX9 port map( A => registers_18_20_port, Z => n332);
   U1474 : HS65_LH_IVX9 port map( A => registers_18_21_port, Z => n331);
   U1475 : HS65_LH_IVX9 port map( A => registers_18_22_port, Z => n330);
   U1476 : HS65_LH_IVX9 port map( A => registers_18_23_port, Z => n329);
   U1477 : HS65_LH_IVX9 port map( A => registers_18_24_port, Z => n328);
   U1478 : HS65_LH_IVX9 port map( A => registers_18_25_port, Z => n327);
   U1479 : HS65_LH_IVX9 port map( A => registers_18_26_port, Z => n326);
   U1480 : HS65_LH_IVX9 port map( A => registers_18_27_port, Z => n325);
   U1481 : HS65_LH_IVX9 port map( A => registers_18_28_port, Z => n324);
   U1482 : HS65_LH_IVX9 port map( A => registers_18_29_port, Z => n323);
   U1483 : HS65_LH_IVX9 port map( A => registers_18_30_port, Z => n322);
   U1484 : HS65_LH_IVX9 port map( A => registers_18_31_port, Z => n321);
   U1485 : HS65_LH_IVX9 port map( A => registers_24_0_port, Z => n320);
   U1486 : HS65_LH_IVX9 port map( A => registers_24_1_port, Z => n319);
   U1487 : HS65_LH_IVX9 port map( A => registers_24_2_port, Z => n318);
   U1488 : HS65_LH_IVX9 port map( A => registers_24_3_port, Z => n317);
   U1489 : HS65_LH_IVX9 port map( A => registers_24_4_port, Z => n316);
   U1490 : HS65_LH_IVX9 port map( A => registers_24_5_port, Z => n315);
   U1491 : HS65_LH_IVX9 port map( A => registers_24_6_port, Z => n314);
   U1492 : HS65_LH_IVX9 port map( A => registers_24_7_port, Z => n313);
   U1493 : HS65_LH_IVX9 port map( A => registers_24_8_port, Z => n312);
   U1494 : HS65_LH_IVX9 port map( A => registers_24_9_port, Z => n311);
   U1495 : HS65_LH_IVX9 port map( A => registers_24_10_port, Z => n310);
   U1496 : HS65_LH_IVX9 port map( A => registers_24_11_port, Z => n309);
   U1497 : HS65_LH_IVX9 port map( A => registers_24_12_port, Z => n308);
   U1498 : HS65_LH_IVX9 port map( A => registers_24_13_port, Z => n307);
   U1499 : HS65_LH_IVX9 port map( A => registers_24_14_port, Z => n306);
   U1500 : HS65_LH_IVX9 port map( A => registers_24_15_port, Z => n305);
   U1501 : HS65_LH_IVX9 port map( A => registers_24_16_port, Z => n304);
   U1502 : HS65_LH_IVX9 port map( A => registers_24_17_port, Z => n303);
   U1503 : HS65_LH_IVX9 port map( A => registers_24_18_port, Z => n302);
   U1504 : HS65_LH_IVX9 port map( A => registers_24_19_port, Z => n301);
   U1505 : HS65_LH_IVX9 port map( A => registers_24_20_port, Z => n300);
   U1506 : HS65_LH_IVX9 port map( A => registers_24_21_port, Z => n299);
   U1507 : HS65_LH_IVX9 port map( A => registers_24_22_port, Z => n298);
   U1508 : HS65_LH_IVX9 port map( A => registers_24_23_port, Z => n297);
   U1509 : HS65_LH_IVX9 port map( A => registers_24_24_port, Z => n296);
   U1510 : HS65_LH_IVX9 port map( A => registers_24_25_port, Z => n295);
   U1511 : HS65_LH_IVX9 port map( A => registers_24_26_port, Z => n294);
   U1512 : HS65_LH_IVX9 port map( A => registers_24_27_port, Z => n293);
   U1513 : HS65_LH_IVX9 port map( A => registers_24_28_port, Z => n292);
   U1514 : HS65_LH_IVX9 port map( A => registers_24_29_port, Z => n291);
   U1515 : HS65_LH_IVX9 port map( A => registers_24_30_port, Z => n290);
   U1516 : HS65_LH_IVX9 port map( A => registers_24_31_port, Z => n289);
   U1517 : HS65_LH_IVX9 port map( A => registers_6_0_port, Z => n512);
   U1518 : HS65_LH_IVX9 port map( A => registers_6_1_port, Z => n511);
   U1519 : HS65_LH_IVX9 port map( A => registers_6_2_port, Z => n510);
   U1520 : HS65_LH_IVX9 port map( A => registers_6_3_port, Z => n509);
   U1521 : HS65_LH_IVX9 port map( A => registers_6_4_port, Z => n508);
   U1522 : HS65_LH_IVX9 port map( A => registers_6_5_port, Z => n507);
   U1523 : HS65_LH_IVX9 port map( A => registers_6_6_port, Z => n506);
   U1524 : HS65_LH_IVX9 port map( A => registers_6_7_port, Z => n505);
   U1525 : HS65_LH_IVX9 port map( A => registers_6_8_port, Z => n504);
   U1526 : HS65_LH_IVX9 port map( A => registers_6_9_port, Z => n503);
   U1527 : HS65_LH_IVX9 port map( A => registers_6_10_port, Z => n502);
   U1528 : HS65_LH_IVX9 port map( A => registers_6_11_port, Z => n501);
   U1529 : HS65_LH_IVX9 port map( A => registers_6_12_port, Z => n500);
   U1530 : HS65_LH_IVX9 port map( A => registers_6_13_port, Z => n499);
   U1531 : HS65_LH_IVX9 port map( A => registers_6_14_port, Z => n498);
   U1532 : HS65_LH_IVX9 port map( A => registers_6_15_port, Z => n497);
   U1533 : HS65_LH_IVX9 port map( A => registers_6_16_port, Z => n496);
   U1534 : HS65_LH_IVX9 port map( A => registers_6_17_port, Z => n495);
   U1535 : HS65_LH_IVX9 port map( A => registers_6_18_port, Z => n494);
   U1536 : HS65_LH_IVX9 port map( A => registers_6_19_port, Z => n493);
   U1537 : HS65_LH_IVX9 port map( A => registers_6_20_port, Z => n492);
   U1538 : HS65_LH_IVX9 port map( A => registers_6_21_port, Z => n491);
   U1539 : HS65_LH_IVX9 port map( A => registers_6_22_port, Z => n490);
   U1540 : HS65_LH_IVX9 port map( A => registers_6_23_port, Z => n489);
   U1541 : HS65_LH_IVX9 port map( A => registers_6_24_port, Z => n488);
   U1542 : HS65_LH_IVX9 port map( A => registers_6_25_port, Z => n487);
   U1543 : HS65_LH_IVX9 port map( A => registers_6_26_port, Z => n486);
   U1544 : HS65_LH_IVX9 port map( A => registers_6_27_port, Z => n485);
   U1545 : HS65_LH_IVX9 port map( A => registers_6_28_port, Z => n484);
   U1546 : HS65_LH_IVX9 port map( A => registers_6_29_port, Z => n483);
   U1547 : HS65_LH_IVX9 port map( A => registers_6_30_port, Z => n482);
   U1548 : HS65_LH_IVX9 port map( A => registers_6_31_port, Z => n481);
   U1549 : HS65_LH_IVX9 port map( A => registers_17_0_port, Z => n384);
   U1550 : HS65_LH_IVX9 port map( A => registers_17_1_port, Z => n383);
   U1551 : HS65_LH_IVX9 port map( A => registers_17_2_port, Z => n382);
   U1552 : HS65_LH_IVX9 port map( A => registers_17_3_port, Z => n381);
   U1553 : HS65_LH_IVX9 port map( A => registers_17_4_port, Z => n380);
   U1554 : HS65_LH_IVX9 port map( A => registers_17_5_port, Z => n379);
   U1555 : HS65_LH_IVX9 port map( A => registers_17_6_port, Z => n378);
   U1556 : HS65_LH_IVX9 port map( A => registers_17_7_port, Z => n377);
   U1557 : HS65_LH_IVX9 port map( A => registers_17_8_port, Z => n376);
   U1558 : HS65_LH_IVX9 port map( A => registers_17_9_port, Z => n375);
   U1559 : HS65_LH_IVX9 port map( A => registers_17_10_port, Z => n374);
   U1560 : HS65_LH_IVX9 port map( A => registers_17_11_port, Z => n373);
   U1561 : HS65_LH_IVX9 port map( A => registers_17_12_port, Z => n372);
   U1562 : HS65_LH_IVX9 port map( A => registers_17_13_port, Z => n371);
   U1563 : HS65_LH_IVX9 port map( A => registers_17_14_port, Z => n370);
   U1564 : HS65_LH_IVX9 port map( A => registers_17_15_port, Z => n369);
   U1565 : HS65_LH_IVX9 port map( A => registers_17_16_port, Z => n368);
   U1566 : HS65_LH_IVX9 port map( A => registers_17_17_port, Z => n367);
   U1567 : HS65_LH_IVX9 port map( A => registers_17_18_port, Z => n366);
   U1568 : HS65_LH_IVX9 port map( A => registers_17_19_port, Z => n365);
   U1569 : HS65_LH_IVX9 port map( A => registers_17_20_port, Z => n364);
   U1570 : HS65_LH_IVX9 port map( A => registers_17_21_port, Z => n363);
   U1571 : HS65_LH_IVX9 port map( A => registers_17_22_port, Z => n362);
   U1572 : HS65_LH_IVX9 port map( A => registers_17_23_port, Z => n361);
   U1573 : HS65_LH_IVX9 port map( A => registers_17_24_port, Z => n360);
   U1574 : HS65_LH_IVX9 port map( A => registers_17_25_port, Z => n359);
   U1575 : HS65_LH_IVX9 port map( A => registers_17_26_port, Z => n358);
   U1576 : HS65_LH_IVX9 port map( A => registers_17_27_port, Z => n357);
   U1577 : HS65_LH_IVX9 port map( A => registers_17_28_port, Z => n356);
   U1578 : HS65_LH_IVX9 port map( A => registers_17_29_port, Z => n355);
   U1579 : HS65_LH_IVX9 port map( A => registers_17_30_port, Z => n354);
   U1580 : HS65_LH_IVX9 port map( A => registers_17_31_port, Z => n353);
   U1581 : HS65_LH_IVX9 port map( A => registers_12_0_port, Z => n448);
   U1582 : HS65_LH_IVX9 port map( A => registers_12_1_port, Z => n447);
   U1583 : HS65_LH_IVX9 port map( A => registers_12_2_port, Z => n446);
   U1584 : HS65_LH_IVX9 port map( A => registers_12_3_port, Z => n445);
   U1585 : HS65_LH_IVX9 port map( A => registers_12_4_port, Z => n444);
   U1586 : HS65_LH_IVX9 port map( A => registers_12_5_port, Z => n443);
   U1587 : HS65_LH_IVX9 port map( A => registers_12_6_port, Z => n442);
   U1588 : HS65_LH_IVX9 port map( A => registers_12_7_port, Z => n441);
   U1589 : HS65_LH_IVX9 port map( A => registers_12_8_port, Z => n440);
   U1590 : HS65_LH_IVX9 port map( A => registers_12_9_port, Z => n439);
   U1591 : HS65_LH_IVX9 port map( A => registers_12_10_port, Z => n438);
   U1592 : HS65_LH_IVX9 port map( A => registers_12_11_port, Z => n437);
   U1593 : HS65_LH_IVX9 port map( A => registers_12_12_port, Z => n436);
   U1594 : HS65_LH_IVX9 port map( A => registers_12_13_port, Z => n435);
   U1595 : HS65_LH_IVX9 port map( A => registers_12_14_port, Z => n434);
   U1596 : HS65_LH_IVX9 port map( A => registers_12_15_port, Z => n433);
   U1597 : HS65_LH_IVX9 port map( A => registers_12_16_port, Z => n432);
   U1598 : HS65_LH_IVX9 port map( A => registers_12_17_port, Z => n431);
   U1599 : HS65_LH_IVX9 port map( A => registers_12_18_port, Z => n430);
   U1600 : HS65_LH_IVX9 port map( A => registers_12_19_port, Z => n429);
   U1601 : HS65_LH_IVX9 port map( A => registers_12_20_port, Z => n428);
   U1602 : HS65_LH_IVX9 port map( A => registers_12_21_port, Z => n427);
   U1603 : HS65_LH_IVX9 port map( A => registers_12_22_port, Z => n426);
   U1604 : HS65_LH_IVX9 port map( A => registers_12_23_port, Z => n425);
   U1605 : HS65_LH_IVX9 port map( A => registers_12_24_port, Z => n424);
   U1606 : HS65_LH_IVX9 port map( A => registers_12_25_port, Z => n423);
   U1607 : HS65_LH_IVX9 port map( A => registers_12_26_port, Z => n422);
   U1608 : HS65_LH_IVX9 port map( A => registers_12_27_port, Z => n421);
   U1609 : HS65_LH_IVX9 port map( A => registers_12_28_port, Z => n420);
   U1610 : HS65_LH_IVX9 port map( A => registers_12_29_port, Z => n419);
   U1611 : HS65_LH_IVX9 port map( A => registers_12_30_port, Z => n418);
   U1612 : HS65_LH_IVX9 port map( A => registers_12_31_port, Z => n417);
   U1613 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6246, C => n6242, 
                           D => registers_13_0_port, Z => n1818);
   U1614 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6246, C => n6242, 
                           D => registers_13_1_port, Z => n1819);
   U1615 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6246, C => n6242, 
                           D => registers_13_2_port, Z => n1820);
   U1616 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6246, C => n6242, 
                           D => registers_13_3_port, Z => n1821);
   U1617 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6246, C => n6242, 
                           D => registers_13_4_port, Z => n1822);
   U1618 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6246, C => n6242, 
                           D => registers_13_5_port, Z => n1823);
   U1619 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6246, C => n6242, 
                           D => registers_13_6_port, Z => n1824);
   U1620 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6246, C => n6242,
                           D => registers_13_7_port, Z => n1825);
   U1621 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6246, C => n6242,
                           D => registers_13_8_port, Z => n1826);
   U1622 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6246, C => n6242,
                           D => registers_13_9_port, Z => n1827);
   U1623 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6246, C => n6242,
                           D => registers_13_10_port, Z => n1828);
   U1624 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6245, C => n6242,
                           D => registers_13_11_port, Z => n1829);
   U1625 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6245, C => n6242,
                           D => registers_13_12_port, Z => n1830);
   U1626 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6245, C => n6243,
                           D => registers_13_13_port, Z => n1831);
   U1627 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6245, C => n6243,
                           D => registers_13_14_port, Z => n1832);
   U1628 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6245, C => n6243,
                           D => registers_13_15_port, Z => n1833);
   U1629 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6245, C => n6243,
                           D => registers_13_16_port, Z => n1834);
   U1630 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6245, C => n6243,
                           D => registers_13_17_port, Z => n1835);
   U1631 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6245, C => n6243,
                           D => registers_13_18_port, Z => n1836);
   U1632 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6245, C => n6243,
                           D => registers_13_19_port, Z => n1837);
   U1633 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6245, C => n6243,
                           D => registers_13_20_port, Z => n1838);
   U1634 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6245, C => n6243,
                           D => registers_13_21_port, Z => n1839);
   U1635 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6245, C => n6243,
                           D => registers_13_22_port, Z => n1840);
   U1636 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6245, C => n6243,
                           D => registers_13_23_port, Z => n1841);
   U1637 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6245, C => n6243,
                           D => registers_13_24_port, Z => n1842);
   U1638 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6245, C => n6243,
                           D => registers_13_25_port, Z => n1843);
   U1639 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6245, C => n6242,
                           D => registers_13_26_port, Z => n1844);
   U1640 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6245, C => n6243,
                           D => registers_13_27_port, Z => n1845);
   U1641 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6245, C => n6242,
                           D => registers_13_28_port, Z => n1846);
   U1642 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6245, C => n6243,
                           D => registers_13_29_port, Z => n1847);
   U1643 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6245, C => n6242,
                           D => registers_13_30_port, Z => n1848);
   U1644 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6244, C => n6243,
                           D => registers_13_31_port, Z => n1849);
   U1645 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6201, C => n6197, 
                           D => registers_4_0_port, Z => n1530);
   U1646 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6201, C => n6197, 
                           D => registers_4_1_port, Z => n1531);
   U1647 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6201, C => n6197, 
                           D => registers_4_2_port, Z => n1532);
   U1648 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6201, C => n6197, 
                           D => registers_4_3_port, Z => n1533);
   U1649 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6201, C => n6197, 
                           D => registers_4_4_port, Z => n1534);
   U1650 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6201, C => n6197, 
                           D => registers_4_5_port, Z => n1535);
   U1651 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6201, C => n6197, 
                           D => registers_4_6_port, Z => n1536);
   U1652 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6201, C => n6197,
                           D => registers_4_7_port, Z => n1537);
   U1653 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6201, C => n6197,
                           D => registers_4_8_port, Z => n1538);
   U1654 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6201, C => n6197,
                           D => registers_4_9_port, Z => n1539);
   U1655 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6201, C => n6197,
                           D => registers_4_10_port, Z => n1540);
   U1656 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6200, C => n6197,
                           D => registers_4_11_port, Z => n1541);
   U1657 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6200, C => n6197,
                           D => registers_4_12_port, Z => n1542);
   U1658 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6200, C => n6198,
                           D => registers_4_13_port, Z => n1543);
   U1659 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6200, C => n6198,
                           D => registers_4_14_port, Z => n1544);
   U1660 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6200, C => n6198,
                           D => registers_4_15_port, Z => n1545);
   U1661 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6200, C => n6198,
                           D => registers_4_16_port, Z => n1546);
   U1662 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6200, C => n6198,
                           D => registers_4_17_port, Z => n1547);
   U1663 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6200, C => n6198,
                           D => registers_4_18_port, Z => n1548);
   U1664 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6200, C => n6198,
                           D => registers_4_19_port, Z => n1549);
   U1665 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6200, C => n6198,
                           D => registers_4_20_port, Z => n1550);
   U1666 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6200, C => n6198,
                           D => registers_4_21_port, Z => n1551);
   U1667 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6200, C => n6198,
                           D => registers_4_22_port, Z => n1552);
   U1668 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6200, C => n6198,
                           D => registers_4_23_port, Z => n1553);
   U1669 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6200, C => n6198,
                           D => registers_4_24_port, Z => n1554);
   U1670 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6200, C => n6198,
                           D => registers_4_25_port, Z => n1555);
   U1671 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6200, C => n6197,
                           D => registers_4_26_port, Z => n1556);
   U1672 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6200, C => n6198,
                           D => registers_4_27_port, Z => n1557);
   U1673 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6200, C => n6197,
                           D => registers_4_28_port, Z => n1558);
   U1674 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6200, C => n6198,
                           D => registers_4_29_port, Z => n1559);
   U1675 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6200, C => n6197,
                           D => registers_4_30_port, Z => n1560);
   U1676 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6199, C => n6198,
                           D => registers_4_31_port, Z => n1561);
   U1677 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6236, C => n6232, 
                           D => registers_11_0_port, Z => n1754);
   U1678 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6236, C => n6232, 
                           D => registers_11_1_port, Z => n1755);
   U1679 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6236, C => n6232, 
                           D => registers_11_2_port, Z => n1756);
   U1680 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6236, C => n6232, 
                           D => registers_11_3_port, Z => n1757);
   U1681 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6236, C => n6232, 
                           D => registers_11_4_port, Z => n1758);
   U1682 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6236, C => n6232, 
                           D => registers_11_5_port, Z => n1759);
   U1683 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6236, C => n6232, 
                           D => registers_11_6_port, Z => n1760);
   U1684 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6236, C => n6232,
                           D => registers_11_7_port, Z => n1761);
   U1685 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6236, C => n6232,
                           D => registers_11_8_port, Z => n1762);
   U1686 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6236, C => n6232,
                           D => registers_11_9_port, Z => n1763);
   U1687 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6236, C => n6232,
                           D => registers_11_10_port, Z => n1764);
   U1688 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6235, C => n6232,
                           D => registers_11_11_port, Z => n1765);
   U1689 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6235, C => n6232,
                           D => registers_11_12_port, Z => n1766);
   U1690 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6235, C => n6233,
                           D => registers_11_13_port, Z => n1767);
   U1691 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6235, C => n6233,
                           D => registers_11_14_port, Z => n1768);
   U1692 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6235, C => n6233,
                           D => registers_11_15_port, Z => n1769);
   U1693 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6235, C => n6233,
                           D => registers_11_16_port, Z => n1770);
   U1694 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6235, C => n6233,
                           D => registers_11_17_port, Z => n1771);
   U1695 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6235, C => n6233,
                           D => registers_11_18_port, Z => n1772);
   U1696 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6235, C => n6233,
                           D => registers_11_19_port, Z => n1773);
   U1697 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6235, C => n6233,
                           D => registers_11_20_port, Z => n1774);
   U1698 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6235, C => n6233,
                           D => registers_11_21_port, Z => n1775);
   U1699 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6235, C => n6233,
                           D => registers_11_22_port, Z => n1776);
   U1700 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6235, C => n6233,
                           D => registers_11_23_port, Z => n1777);
   U1701 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6235, C => n6233,
                           D => registers_11_24_port, Z => n1778);
   U1702 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6235, C => n6233,
                           D => registers_11_25_port, Z => n1779);
   U1703 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6235, C => n6232,
                           D => registers_11_26_port, Z => n1780);
   U1704 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6235, C => n6233,
                           D => registers_11_27_port, Z => n1781);
   U1705 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6235, C => n6232,
                           D => registers_11_28_port, Z => n1782);
   U1706 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6235, C => n6233,
                           D => registers_11_29_port, Z => n1783);
   U1707 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6235, C => n6232,
                           D => registers_11_30_port, Z => n1784);
   U1708 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6234, C => n6233,
                           D => registers_11_31_port, Z => n1785);
   U1709 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6196, C => n6192, 
                           D => registers_3_0_port, Z => n1498);
   U1710 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6196, C => n6192, 
                           D => registers_3_1_port, Z => n1499);
   U1711 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6196, C => n6192, 
                           D => registers_3_2_port, Z => n1500);
   U1712 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6196, C => n6192, 
                           D => registers_3_3_port, Z => n1501);
   U1713 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6196, C => n6192, 
                           D => registers_3_4_port, Z => n1502);
   U1714 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6196, C => n6192, 
                           D => registers_3_5_port, Z => n1503);
   U1715 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6196, C => n6192, 
                           D => registers_3_6_port, Z => n1504);
   U1716 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6196, C => n6192,
                           D => registers_3_7_port, Z => n1505);
   U1717 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6196, C => n6192,
                           D => registers_3_8_port, Z => n1506);
   U1718 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6196, C => n6192,
                           D => registers_3_9_port, Z => n1507);
   U1719 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6196, C => n6192,
                           D => registers_3_10_port, Z => n1508);
   U1720 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6195, C => n6192,
                           D => registers_3_11_port, Z => n1509);
   U1721 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6195, C => n6192,
                           D => registers_3_12_port, Z => n1510);
   U1722 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6195, C => n6193,
                           D => registers_3_13_port, Z => n1511);
   U1723 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6195, C => n6193,
                           D => registers_3_14_port, Z => n1512);
   U1724 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6195, C => n6193,
                           D => registers_3_15_port, Z => n1513);
   U1725 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6195, C => n6193,
                           D => registers_3_16_port, Z => n1514);
   U1726 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6195, C => n6193,
                           D => registers_3_17_port, Z => n1515);
   U1727 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6195, C => n6193,
                           D => registers_3_18_port, Z => n1516);
   U1728 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6195, C => n6193,
                           D => registers_3_19_port, Z => n1517);
   U1729 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6195, C => n6193,
                           D => registers_3_20_port, Z => n1518);
   U1730 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6195, C => n6193,
                           D => registers_3_21_port, Z => n1519);
   U1731 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6195, C => n6193,
                           D => registers_3_22_port, Z => n1520);
   U1732 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6195, C => n6193,
                           D => registers_3_23_port, Z => n1521);
   U1733 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6195, C => n6193,
                           D => registers_3_24_port, Z => n1522);
   U1734 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6195, C => n6193,
                           D => registers_3_25_port, Z => n1523);
   U1735 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6195, C => n6192,
                           D => registers_3_26_port, Z => n1524);
   U1736 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6195, C => n6193,
                           D => registers_3_27_port, Z => n1525);
   U1737 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6195, C => n6192,
                           D => registers_3_28_port, Z => n1526);
   U1738 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6195, C => n6193,
                           D => registers_3_29_port, Z => n1527);
   U1739 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6195, C => n6192,
                           D => registers_3_30_port, Z => n1528);
   U1740 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6194, C => n6193,
                           D => registers_3_31_port, Z => n1529);
   U1741 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6191, C => n6187, 
                           D => registers_2_0_port, Z => n1466);
   U1742 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6191, C => n6187, 
                           D => registers_2_1_port, Z => n1467);
   U1743 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6191, C => n6187, 
                           D => registers_2_2_port, Z => n1468);
   U1744 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6191, C => n6187, 
                           D => registers_2_3_port, Z => n1469);
   U1745 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6191, C => n6187, 
                           D => registers_2_4_port, Z => n1470);
   U1746 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6191, C => n6187, 
                           D => registers_2_5_port, Z => n1471);
   U1747 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6191, C => n6187, 
                           D => registers_2_6_port, Z => n1472);
   U1748 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6191, C => n6187,
                           D => registers_2_7_port, Z => n1473);
   U1749 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6191, C => n6187,
                           D => registers_2_8_port, Z => n1474);
   U1750 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6191, C => n6187,
                           D => registers_2_9_port, Z => n1475);
   U1751 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6191, C => n6187,
                           D => registers_2_10_port, Z => n1476);
   U1752 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6190, C => n6187,
                           D => registers_2_11_port, Z => n1477);
   U1753 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6190, C => n6187,
                           D => registers_2_12_port, Z => n1478);
   U1754 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6190, C => n6188,
                           D => registers_2_13_port, Z => n1479);
   U1755 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6190, C => n6188,
                           D => registers_2_14_port, Z => n1480);
   U1756 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6190, C => n6188,
                           D => registers_2_15_port, Z => n1481);
   U1757 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6190, C => n6188,
                           D => registers_2_16_port, Z => n1482);
   U1758 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6190, C => n6188,
                           D => registers_2_17_port, Z => n1483);
   U1759 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6190, C => n6188,
                           D => registers_2_18_port, Z => n1484);
   U1760 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6190, C => n6188,
                           D => registers_2_19_port, Z => n1485);
   U1761 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6190, C => n6188,
                           D => registers_2_20_port, Z => n1486);
   U1762 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6190, C => n6188,
                           D => registers_2_21_port, Z => n1487);
   U1763 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6190, C => n6188,
                           D => registers_2_22_port, Z => n1488);
   U1764 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6190, C => n6188,
                           D => registers_2_23_port, Z => n1489);
   U1765 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6190, C => n6188,
                           D => registers_2_24_port, Z => n1490);
   U1766 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6190, C => n6188,
                           D => registers_2_25_port, Z => n1491);
   U1767 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6190, C => n6187,
                           D => registers_2_26_port, Z => n1492);
   U1768 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6190, C => n6188,
                           D => registers_2_27_port, Z => n1493);
   U1769 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6190, C => n6187,
                           D => registers_2_28_port, Z => n1494);
   U1770 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6190, C => n6188,
                           D => registers_2_29_port, Z => n1495);
   U1771 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6190, C => n6187,
                           D => registers_2_30_port, Z => n1496);
   U1772 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6189, C => n6188,
                           D => registers_2_31_port, Z => n1497);
   U1773 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n6206, C => n6202, 
                           D => registers_5_0_port, Z => n1562);
   U1774 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n6206, C => n6202, 
                           D => registers_5_1_port, Z => n1563);
   U1775 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n6206, C => n6202, 
                           D => registers_5_2_port, Z => n1564);
   U1776 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n6206, C => n6202, 
                           D => registers_5_3_port, Z => n1565);
   U1777 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n6206, C => n6202, 
                           D => registers_5_4_port, Z => n1566);
   U1778 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n6206, C => n6202, 
                           D => registers_5_5_port, Z => n1567);
   U1779 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n6206, C => n6202, 
                           D => registers_5_6_port, Z => n1568);
   U1780 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n6206, C => n6202,
                           D => registers_5_7_port, Z => n1569);
   U1781 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n6206, C => n6202,
                           D => registers_5_8_port, Z => n1570);
   U1782 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n6206, C => n6202,
                           D => registers_5_9_port, Z => n1571);
   U1783 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n6206, C => n6202,
                           D => registers_5_10_port, Z => n1572);
   U1784 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n6205, C => n6202,
                           D => registers_5_11_port, Z => n1573);
   U1785 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n6205, C => n6202,
                           D => registers_5_12_port, Z => n1574);
   U1786 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n6205, C => n6203,
                           D => registers_5_13_port, Z => n1575);
   U1787 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n6205, C => n6203,
                           D => registers_5_14_port, Z => n1576);
   U1788 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n6205, C => n6203,
                           D => registers_5_15_port, Z => n1577);
   U1789 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n6205, C => n6203,
                           D => registers_5_16_port, Z => n1578);
   U1790 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n6205, C => n6203,
                           D => registers_5_17_port, Z => n1579);
   U1791 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n6205, C => n6203,
                           D => registers_5_18_port, Z => n1580);
   U1792 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n6205, C => n6203,
                           D => registers_5_19_port, Z => n1581);
   U1793 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n6205, C => n6203,
                           D => registers_5_20_port, Z => n1582);
   U1794 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n6205, C => n6203,
                           D => registers_5_21_port, Z => n1583);
   U1795 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n6205, C => n6203,
                           D => registers_5_22_port, Z => n1584);
   U1796 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n6205, C => n6203,
                           D => registers_5_23_port, Z => n1585);
   U1797 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n6205, C => n6203,
                           D => registers_5_24_port, Z => n1586);
   U1798 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n6205, C => n6203,
                           D => registers_5_25_port, Z => n1587);
   U1799 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n6205, C => n6202,
                           D => registers_5_26_port, Z => n1588);
   U1800 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n6205, C => n6203,
                           D => registers_5_27_port, Z => n1589);
   U1801 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n6205, C => n6202,
                           D => registers_5_28_port, Z => n1590);
   U1802 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n6205, C => n6203,
                           D => registers_5_29_port, Z => n1591);
   U1803 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n6205, C => n6202,
                           D => registers_5_30_port, Z => n1592);
   U1804 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n6204, C => n6203,
                           D => registers_5_31_port, Z => n1593);
   U1805 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_0_port, C => 
                           regfile_i(3), D => n6186, Z => n1434);
   U1806 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_1_port, C => 
                           regfile_i(4), D => n6186, Z => n1435);
   U1807 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_2_port, C => 
                           regfile_i(5), D => n6186, Z => n1436);
   U1808 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_3_port, C => 
                           regfile_i(6), D => n6186, Z => n1437);
   U1809 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_4_port, C => 
                           regfile_i(7), D => n6186, Z => n1438);
   U1810 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_5_port, C => 
                           regfile_i(8), D => n6186, Z => n1439);
   U1811 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_6_port, C => 
                           regfile_i(9), D => n6186, Z => n1440);
   U1812 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_7_port, C => 
                           regfile_i(10), D => n6186, Z => n1441);
   U1813 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_8_port, C => 
                           regfile_i(11), D => n6186, Z => n1442);
   U1814 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_9_port, C => 
                           regfile_i(12), D => n6186, Z => n1443);
   U1815 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_10_port, C => 
                           regfile_i(13), D => n6186, Z => n1444);
   U1816 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_11_port, C => 
                           regfile_i(14), D => n6185, Z => n1445);
   U1817 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_12_port, C => 
                           regfile_i(15), D => n6185, Z => n1446);
   U1818 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_13_port, C => 
                           regfile_i(16), D => n6185, Z => n1447);
   U1819 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_14_port, C => 
                           regfile_i(17), D => n6185, Z => n1448);
   U1820 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_15_port, C => 
                           regfile_i(18), D => n6185, Z => n1449);
   U1821 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_16_port, C => 
                           regfile_i(19), D => n6185, Z => n1450);
   U1822 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_17_port, C => 
                           regfile_i(20), D => n6185, Z => n1451);
   U1823 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_18_port, C => 
                           regfile_i(21), D => n6185, Z => n1452);
   U1824 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_19_port, C => 
                           regfile_i(22), D => n6185, Z => n1453);
   U1825 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_20_port, C => 
                           regfile_i(23), D => n6185, Z => n1454);
   U1826 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_21_port, C => 
                           regfile_i(24), D => n6185, Z => n1455);
   U1827 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_22_port, C => 
                           regfile_i(25), D => n6185, Z => n1456);
   U1828 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_23_port, C => 
                           regfile_i(26), D => n6185, Z => n1457);
   U1829 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_24_port, C => 
                           regfile_i(27), D => n6185, Z => n1458);
   U1830 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_25_port, C => 
                           regfile_i(28), D => n6185, Z => n1459);
   U1831 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_26_port, C => 
                           regfile_i(29), D => n6185, Z => n1460);
   U1832 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_27_port, C => 
                           regfile_i(30), D => n6185, Z => n1461);
   U1833 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_28_port, C => 
                           regfile_i(31), D => n6185, Z => n1462);
   U1834 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_29_port, C => 
                           regfile_i(32), D => n6185, Z => n1463);
   U1835 : HS65_LH_AO22X9 port map( A => n6182, B => registers_1_30_port, C => 
                           regfile_i(33), D => n6185, Z => n1464);
   U1836 : HS65_LH_AO22X9 port map( A => n6183, B => registers_1_31_port, C => 
                           regfile_i(34), D => n6184, Z => n1465);
   U1837 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_0_port, C => 
                           regfile_i(3), D => n6336, Z => n2394);
   U1838 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_1_port, C => 
                           regfile_i(4), D => n6336, Z => n2395);
   U1839 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_2_port, C => 
                           regfile_i(5), D => n6336, Z => n2396);
   U1840 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_3_port, C => 
                           regfile_i(6), D => n6336, Z => n2397);
   U1841 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_4_port, C => 
                           regfile_i(7), D => n6336, Z => n2398);
   U1842 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_5_port, C => 
                           regfile_i(8), D => n6336, Z => n2399);
   U1843 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_6_port, C => 
                           regfile_i(9), D => n6336, Z => n2400);
   U1844 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_7_port, C => 
                           regfile_i(10), D => n6336, Z => n2401);
   U1845 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_8_port, C => 
                           regfile_i(11), D => n6336, Z => n2402);
   U1846 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_9_port, C => 
                           regfile_i(12), D => n6336, Z => n2403);
   U1847 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_10_port, C =>
                           regfile_i(13), D => n6336, Z => n2404);
   U1848 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_11_port, C =>
                           regfile_i(14), D => n6335, Z => n2405);
   U1849 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_12_port, C =>
                           regfile_i(15), D => n6335, Z => n2406);
   U1850 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_13_port, C =>
                           regfile_i(16), D => n6335, Z => n2407);
   U1851 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_14_port, C =>
                           regfile_i(17), D => n6335, Z => n2408);
   U1852 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_15_port, C =>
                           regfile_i(18), D => n6335, Z => n2409);
   U1853 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_16_port, C =>
                           regfile_i(19), D => n6335, Z => n2410);
   U1854 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_17_port, C =>
                           regfile_i(20), D => n6335, Z => n2411);
   U1855 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_18_port, C =>
                           regfile_i(21), D => n6335, Z => n2412);
   U1856 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_19_port, C =>
                           regfile_i(22), D => n6335, Z => n2413);
   U1857 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_20_port, C =>
                           regfile_i(23), D => n6335, Z => n2414);
   U1858 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_21_port, C =>
                           regfile_i(24), D => n6335, Z => n2415);
   U1859 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_22_port, C =>
                           regfile_i(25), D => n6335, Z => n2416);
   U1860 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_23_port, C =>
                           regfile_i(26), D => n6335, Z => n2417);
   U1861 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_24_port, C =>
                           regfile_i(27), D => n6335, Z => n2418);
   U1862 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_25_port, C =>
                           regfile_i(28), D => n6335, Z => n2419);
   U1863 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_26_port, C =>
                           regfile_i(29), D => n6335, Z => n2420);
   U1864 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_27_port, C =>
                           regfile_i(30), D => n6335, Z => n2421);
   U1865 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_28_port, C =>
                           regfile_i(31), D => n6335, Z => n2422);
   U1866 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_29_port, C =>
                           regfile_i(32), D => n6335, Z => n2423);
   U1867 : HS65_LH_AO22X9 port map( A => n6332, B => registers_31_30_port, C =>
                           regfile_i(33), D => n6335, Z => n2424);
   U1868 : HS65_LH_AO22X9 port map( A => n6333, B => registers_31_31_port, C =>
                           regfile_i(34), D => n6334, Z => n2425);
   U1869 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_0_port, C => 
                           regfile_i(3), D => n6276, Z => n2010);
   U1870 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_1_port, C => 
                           regfile_i(4), D => n6276, Z => n2011);
   U1871 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_2_port, C => 
                           regfile_i(5), D => n6276, Z => n2012);
   U1872 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_3_port, C => 
                           regfile_i(6), D => n6276, Z => n2013);
   U1873 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_4_port, C => 
                           regfile_i(7), D => n6276, Z => n2014);
   U1874 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_5_port, C => 
                           regfile_i(8), D => n6276, Z => n2015);
   U1875 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_6_port, C => 
                           regfile_i(9), D => n6276, Z => n2016);
   U1876 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_7_port, C => 
                           regfile_i(10), D => n6276, Z => n2017);
   U1877 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_8_port, C => 
                           regfile_i(11), D => n6276, Z => n2018);
   U1878 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_9_port, C => 
                           regfile_i(12), D => n6276, Z => n2019);
   U1879 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_10_port, C =>
                           regfile_i(13), D => n6276, Z => n2020);
   U1880 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_11_port, C =>
                           regfile_i(14), D => n6275, Z => n2021);
   U1881 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_12_port, C =>
                           regfile_i(15), D => n6275, Z => n2022);
   U1882 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_13_port, C =>
                           regfile_i(16), D => n6275, Z => n2023);
   U1883 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_14_port, C =>
                           regfile_i(17), D => n6275, Z => n2024);
   U1884 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_15_port, C =>
                           regfile_i(18), D => n6275, Z => n2025);
   U1885 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_16_port, C =>
                           regfile_i(19), D => n6275, Z => n2026);
   U1886 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_17_port, C =>
                           regfile_i(20), D => n6275, Z => n2027);
   U1887 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_18_port, C =>
                           regfile_i(21), D => n6275, Z => n2028);
   U1888 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_19_port, C =>
                           regfile_i(22), D => n6275, Z => n2029);
   U1889 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_20_port, C =>
                           regfile_i(23), D => n6275, Z => n2030);
   U1890 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_21_port, C =>
                           regfile_i(24), D => n6275, Z => n2031);
   U1891 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_22_port, C =>
                           regfile_i(25), D => n6275, Z => n2032);
   U1892 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_23_port, C =>
                           regfile_i(26), D => n6275, Z => n2033);
   U1893 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_24_port, C =>
                           regfile_i(27), D => n6275, Z => n2034);
   U1894 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_25_port, C =>
                           regfile_i(28), D => n6275, Z => n2035);
   U1895 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_26_port, C =>
                           regfile_i(29), D => n6275, Z => n2036);
   U1896 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_27_port, C =>
                           regfile_i(30), D => n6275, Z => n2037);
   U1897 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_28_port, C =>
                           regfile_i(31), D => n6275, Z => n2038);
   U1898 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_29_port, C =>
                           regfile_i(32), D => n6275, Z => n2039);
   U1899 : HS65_LH_AO22X9 port map( A => n6272, B => registers_19_30_port, C =>
                           regfile_i(33), D => n6275, Z => n2040);
   U1900 : HS65_LH_AO22X9 port map( A => n6273, B => registers_19_31_port, C =>
                           regfile_i(34), D => n6274, Z => n2041);
   U1901 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_0_port, C => 
                           regfile_i(3), D => n6216, Z => n1626);
   U1902 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_1_port, C => 
                           regfile_i(4), D => n6216, Z => n1627);
   U1903 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_2_port, C => 
                           regfile_i(5), D => n6216, Z => n1628);
   U1904 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_3_port, C => 
                           regfile_i(6), D => n6216, Z => n1629);
   U1905 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_4_port, C => 
                           regfile_i(7), D => n6216, Z => n1630);
   U1906 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_5_port, C => 
                           regfile_i(8), D => n6216, Z => n1631);
   U1907 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_6_port, C => 
                           regfile_i(9), D => n6216, Z => n1632);
   U1908 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_7_port, C => 
                           regfile_i(10), D => n6216, Z => n1633);
   U1909 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_8_port, C => 
                           regfile_i(11), D => n6216, Z => n1634);
   U1910 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_9_port, C => 
                           regfile_i(12), D => n6216, Z => n1635);
   U1911 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_10_port, C => 
                           regfile_i(13), D => n6216, Z => n1636);
   U1912 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_11_port, C => 
                           regfile_i(14), D => n6215, Z => n1637);
   U1913 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_12_port, C => 
                           regfile_i(15), D => n6215, Z => n1638);
   U1914 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_13_port, C => 
                           regfile_i(16), D => n6215, Z => n1639);
   U1915 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_14_port, C => 
                           regfile_i(17), D => n6215, Z => n1640);
   U1916 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_15_port, C => 
                           regfile_i(18), D => n6215, Z => n1641);
   U1917 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_16_port, C => 
                           regfile_i(19), D => n6215, Z => n1642);
   U1918 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_17_port, C => 
                           regfile_i(20), D => n6215, Z => n1643);
   U1919 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_18_port, C => 
                           regfile_i(21), D => n6215, Z => n1644);
   U1920 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_19_port, C => 
                           regfile_i(22), D => n6215, Z => n1645);
   U1921 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_20_port, C => 
                           regfile_i(23), D => n6215, Z => n1646);
   U1922 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_21_port, C => 
                           regfile_i(24), D => n6215, Z => n1647);
   U1923 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_22_port, C => 
                           regfile_i(25), D => n6215, Z => n1648);
   U1924 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_23_port, C => 
                           regfile_i(26), D => n6215, Z => n1649);
   U1925 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_24_port, C => 
                           regfile_i(27), D => n6215, Z => n1650);
   U1926 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_25_port, C => 
                           regfile_i(28), D => n6215, Z => n1651);
   U1927 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_26_port, C => 
                           regfile_i(29), D => n6215, Z => n1652);
   U1928 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_27_port, C => 
                           regfile_i(30), D => n6215, Z => n1653);
   U1929 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_28_port, C => 
                           regfile_i(31), D => n6215, Z => n1654);
   U1930 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_29_port, C => 
                           regfile_i(32), D => n6215, Z => n1655);
   U1931 : HS65_LH_AO22X9 port map( A => n6212, B => registers_7_30_port, C => 
                           regfile_i(33), D => n6215, Z => n1656);
   U1932 : HS65_LH_AO22X9 port map( A => n6213, B => registers_7_31_port, C => 
                           regfile_i(34), D => n6214, Z => n1657);
   U1933 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_0_port, C => 
                           regfile_i(3), D => n6281, Z => n2042);
   U1934 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_1_port, C => 
                           regfile_i(4), D => n6281, Z => n2043);
   U1935 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_2_port, C => 
                           regfile_i(5), D => n6281, Z => n2044);
   U1936 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_3_port, C => 
                           regfile_i(6), D => n6281, Z => n2045);
   U1937 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_4_port, C => 
                           regfile_i(7), D => n6281, Z => n2046);
   U1938 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_5_port, C => 
                           regfile_i(8), D => n6281, Z => n2047);
   U1939 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_6_port, C => 
                           regfile_i(9), D => n6281, Z => n2048);
   U1940 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_7_port, C => 
                           regfile_i(10), D => n6281, Z => n2049);
   U1941 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_8_port, C => 
                           regfile_i(11), D => n6281, Z => n2050);
   U1942 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_9_port, C => 
                           regfile_i(12), D => n6281, Z => n2051);
   U1943 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_10_port, C =>
                           regfile_i(13), D => n6281, Z => n2052);
   U1944 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_11_port, C =>
                           regfile_i(14), D => n6280, Z => n2053);
   U1945 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_12_port, C =>
                           regfile_i(15), D => n6280, Z => n2054);
   U1946 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_13_port, C =>
                           regfile_i(16), D => n6280, Z => n2055);
   U1947 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_14_port, C =>
                           regfile_i(17), D => n6280, Z => n2056);
   U1948 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_15_port, C =>
                           regfile_i(18), D => n6280, Z => n2057);
   U1949 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_16_port, C =>
                           regfile_i(19), D => n6280, Z => n2058);
   U1950 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_17_port, C =>
                           regfile_i(20), D => n6280, Z => n2059);
   U1951 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_18_port, C =>
                           regfile_i(21), D => n6280, Z => n2060);
   U1952 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_19_port, C =>
                           regfile_i(22), D => n6280, Z => n2061);
   U1953 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_20_port, C =>
                           regfile_i(23), D => n6280, Z => n2062);
   U1954 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_21_port, C =>
                           regfile_i(24), D => n6280, Z => n2063);
   U1955 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_22_port, C =>
                           regfile_i(25), D => n6280, Z => n2064);
   U1956 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_23_port, C =>
                           regfile_i(26), D => n6280, Z => n2065);
   U1957 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_24_port, C =>
                           regfile_i(27), D => n6280, Z => n2066);
   U1958 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_25_port, C =>
                           regfile_i(28), D => n6280, Z => n2067);
   U1959 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_26_port, C =>
                           regfile_i(29), D => n6280, Z => n2068);
   U1960 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_27_port, C =>
                           regfile_i(30), D => n6280, Z => n2069);
   U1961 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_28_port, C =>
                           regfile_i(31), D => n6280, Z => n2070);
   U1962 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_29_port, C =>
                           regfile_i(32), D => n6280, Z => n2071);
   U1963 : HS65_LH_AO22X9 port map( A => n6277, B => registers_20_30_port, C =>
                           regfile_i(33), D => n6280, Z => n2072);
   U1964 : HS65_LH_AO22X9 port map( A => n6278, B => registers_20_31_port, C =>
                           regfile_i(34), D => n6279, Z => n2073);
   U1965 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_0_port, C => 
                           regfile_i(3), D => n6286, Z => n2074);
   U1966 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_1_port, C => 
                           regfile_i(4), D => n6286, Z => n2075);
   U1967 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_2_port, C => 
                           regfile_i(5), D => n6286, Z => n2076);
   U1968 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_3_port, C => 
                           regfile_i(6), D => n6286, Z => n2077);
   U1969 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_4_port, C => 
                           regfile_i(7), D => n6286, Z => n2078);
   U1970 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_5_port, C => 
                           regfile_i(8), D => n6286, Z => n2079);
   U1971 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_6_port, C => 
                           regfile_i(9), D => n6286, Z => n2080);
   U1972 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_7_port, C => 
                           regfile_i(10), D => n6286, Z => n2081);
   U1973 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_8_port, C => 
                           regfile_i(11), D => n6286, Z => n2082);
   U1974 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_9_port, C => 
                           regfile_i(12), D => n6286, Z => n2083);
   U1975 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_10_port, C =>
                           regfile_i(13), D => n6286, Z => n2084);
   U1976 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_11_port, C =>
                           regfile_i(14), D => n6285, Z => n2085);
   U1977 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_12_port, C =>
                           regfile_i(15), D => n6285, Z => n2086);
   U1978 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_13_port, C =>
                           regfile_i(16), D => n6285, Z => n2087);
   U1979 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_14_port, C =>
                           regfile_i(17), D => n6285, Z => n2088);
   U1980 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_15_port, C =>
                           regfile_i(18), D => n6285, Z => n2089);
   U1981 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_16_port, C =>
                           regfile_i(19), D => n6285, Z => n2090);
   U1982 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_17_port, C =>
                           regfile_i(20), D => n6285, Z => n2091);
   U1983 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_18_port, C =>
                           regfile_i(21), D => n6285, Z => n2092);
   U1984 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_19_port, C =>
                           regfile_i(22), D => n6285, Z => n2093);
   U1985 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_20_port, C =>
                           regfile_i(23), D => n6285, Z => n2094);
   U1986 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_21_port, C =>
                           regfile_i(24), D => n6285, Z => n2095);
   U1987 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_22_port, C =>
                           regfile_i(25), D => n6285, Z => n2096);
   U1988 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_23_port, C =>
                           regfile_i(26), D => n6285, Z => n2097);
   U1989 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_24_port, C =>
                           regfile_i(27), D => n6285, Z => n2098);
   U1990 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_25_port, C =>
                           regfile_i(28), D => n6285, Z => n2099);
   U1991 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_26_port, C =>
                           regfile_i(29), D => n6285, Z => n2100);
   U1992 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_27_port, C =>
                           regfile_i(30), D => n6285, Z => n2101);
   U1993 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_28_port, C =>
                           regfile_i(31), D => n6285, Z => n2102);
   U1994 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_29_port, C =>
                           regfile_i(32), D => n6285, Z => n2103);
   U1995 : HS65_LH_AO22X9 port map( A => n6282, B => registers_21_30_port, C =>
                           regfile_i(33), D => n6285, Z => n2104);
   U1996 : HS65_LH_AO22X9 port map( A => n6283, B => registers_21_31_port, C =>
                           regfile_i(34), D => n6284, Z => n2105);
   U1997 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_0_port, C => 
                           regfile_i(3), D => n6331, Z => n2362);
   U1998 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_1_port, C => 
                           regfile_i(4), D => n6331, Z => n2363);
   U1999 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_2_port, C => 
                           regfile_i(5), D => n6331, Z => n2364);
   U2000 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_3_port, C => 
                           regfile_i(6), D => n6331, Z => n2365);
   U2001 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_4_port, C => 
                           regfile_i(7), D => n6331, Z => n2366);
   U2002 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_5_port, C => 
                           regfile_i(8), D => n6331, Z => n2367);
   U2003 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_6_port, C => 
                           regfile_i(9), D => n6331, Z => n2368);
   U2004 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_7_port, C => 
                           regfile_i(10), D => n6331, Z => n2369);
   U2005 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_8_port, C => 
                           regfile_i(11), D => n6331, Z => n2370);
   U2006 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_9_port, C => 
                           regfile_i(12), D => n6331, Z => n2371);
   U2007 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_10_port, C =>
                           regfile_i(13), D => n6331, Z => n2372);
   U2008 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_11_port, C =>
                           regfile_i(14), D => n6330, Z => n2373);
   U2009 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_12_port, C =>
                           regfile_i(15), D => n6330, Z => n2374);
   U2010 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_13_port, C =>
                           regfile_i(16), D => n6330, Z => n2375);
   U2011 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_14_port, C =>
                           regfile_i(17), D => n6330, Z => n2376);
   U2012 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_15_port, C =>
                           regfile_i(18), D => n6330, Z => n2377);
   U2013 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_16_port, C =>
                           regfile_i(19), D => n6330, Z => n2378);
   U2014 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_17_port, C =>
                           regfile_i(20), D => n6330, Z => n2379);
   U2015 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_18_port, C =>
                           regfile_i(21), D => n6330, Z => n2380);
   U2016 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_19_port, C =>
                           regfile_i(22), D => n6330, Z => n2381);
   U2017 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_20_port, C =>
                           regfile_i(23), D => n6330, Z => n2382);
   U2018 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_21_port, C =>
                           regfile_i(24), D => n6330, Z => n2383);
   U2019 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_22_port, C =>
                           regfile_i(25), D => n6330, Z => n2384);
   U2020 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_23_port, C =>
                           regfile_i(26), D => n6330, Z => n2385);
   U2021 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_24_port, C =>
                           regfile_i(27), D => n6330, Z => n2386);
   U2022 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_25_port, C =>
                           regfile_i(28), D => n6330, Z => n2387);
   U2023 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_26_port, C =>
                           regfile_i(29), D => n6330, Z => n2388);
   U2024 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_27_port, C =>
                           regfile_i(30), D => n6330, Z => n2389);
   U2025 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_28_port, C =>
                           regfile_i(31), D => n6330, Z => n2390);
   U2026 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_29_port, C =>
                           regfile_i(32), D => n6330, Z => n2391);
   U2027 : HS65_LH_AO22X9 port map( A => n6327, B => registers_30_30_port, C =>
                           regfile_i(33), D => n6330, Z => n2392);
   U2028 : HS65_LH_AO22X9 port map( A => n6328, B => registers_30_31_port, C =>
                           regfile_i(34), D => n6329, Z => n2393);
   U2029 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_0_port, C => 
                           regfile_i(3), D => n6296, Z => n2138);
   U2030 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_1_port, C => 
                           regfile_i(4), D => n6296, Z => n2139);
   U2031 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_2_port, C => 
                           regfile_i(5), D => n6296, Z => n2140);
   U2032 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_3_port, C => 
                           regfile_i(6), D => n6296, Z => n2141);
   U2033 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_4_port, C => 
                           regfile_i(7), D => n6296, Z => n2142);
   U2034 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_5_port, C => 
                           regfile_i(8), D => n6296, Z => n2143);
   U2035 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_6_port, C => 
                           regfile_i(9), D => n6296, Z => n2144);
   U2036 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_7_port, C => 
                           regfile_i(10), D => n6296, Z => n2145);
   U2037 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_8_port, C => 
                           regfile_i(11), D => n6296, Z => n2146);
   U2038 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_9_port, C => 
                           regfile_i(12), D => n6296, Z => n2147);
   U2039 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_10_port, C =>
                           regfile_i(13), D => n6296, Z => n2148);
   U2040 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_11_port, C =>
                           regfile_i(14), D => n6295, Z => n2149);
   U2041 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_12_port, C =>
                           regfile_i(15), D => n6295, Z => n2150);
   U2042 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_13_port, C =>
                           regfile_i(16), D => n6295, Z => n2151);
   U2043 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_14_port, C =>
                           regfile_i(17), D => n6295, Z => n2152);
   U2044 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_15_port, C =>
                           regfile_i(18), D => n6295, Z => n2153);
   U2045 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_16_port, C =>
                           regfile_i(19), D => n6295, Z => n2154);
   U2046 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_17_port, C =>
                           regfile_i(20), D => n6295, Z => n2155);
   U2047 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_18_port, C =>
                           regfile_i(21), D => n6295, Z => n2156);
   U2048 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_19_port, C =>
                           regfile_i(22), D => n6295, Z => n2157);
   U2049 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_20_port, C =>
                           regfile_i(23), D => n6295, Z => n2158);
   U2050 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_21_port, C =>
                           regfile_i(24), D => n6295, Z => n2159);
   U2051 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_22_port, C =>
                           regfile_i(25), D => n6295, Z => n2160);
   U2052 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_23_port, C =>
                           regfile_i(26), D => n6295, Z => n2161);
   U2053 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_24_port, C =>
                           regfile_i(27), D => n6295, Z => n2162);
   U2054 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_25_port, C =>
                           regfile_i(28), D => n6295, Z => n2163);
   U2055 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_26_port, C =>
                           regfile_i(29), D => n6295, Z => n2164);
   U2056 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_27_port, C =>
                           regfile_i(30), D => n6295, Z => n2165);
   U2057 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_28_port, C =>
                           regfile_i(31), D => n6295, Z => n2166);
   U2058 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_29_port, C =>
                           regfile_i(32), D => n6295, Z => n2167);
   U2059 : HS65_LH_AO22X9 port map( A => n6292, B => registers_23_30_port, C =>
                           regfile_i(33), D => n6295, Z => n2168);
   U2060 : HS65_LH_AO22X9 port map( A => n6293, B => registers_23_31_port, C =>
                           regfile_i(34), D => n6294, Z => n2169);
   U2061 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_0_port, C => 
                           regfile_i(3), D => n6291, Z => n2106);
   U2062 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_1_port, C => 
                           regfile_i(4), D => n6291, Z => n2107);
   U2063 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_2_port, C => 
                           regfile_i(5), D => n6291, Z => n2108);
   U2064 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_3_port, C => 
                           regfile_i(6), D => n6291, Z => n2109);
   U2065 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_4_port, C => 
                           regfile_i(7), D => n6291, Z => n2110);
   U2066 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_5_port, C => 
                           regfile_i(8), D => n6291, Z => n2111);
   U2067 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_6_port, C => 
                           regfile_i(9), D => n6291, Z => n2112);
   U2068 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_7_port, C => 
                           regfile_i(10), D => n6291, Z => n2113);
   U2069 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_8_port, C => 
                           regfile_i(11), D => n6291, Z => n2114);
   U2070 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_9_port, C => 
                           regfile_i(12), D => n6291, Z => n2115);
   U2071 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_10_port, C =>
                           regfile_i(13), D => n6291, Z => n2116);
   U2072 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_11_port, C =>
                           regfile_i(14), D => n6290, Z => n2117);
   U2073 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_12_port, C =>
                           regfile_i(15), D => n6290, Z => n2118);
   U2074 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_13_port, C =>
                           regfile_i(16), D => n6290, Z => n2119);
   U2075 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_14_port, C =>
                           regfile_i(17), D => n6290, Z => n2120);
   U2076 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_15_port, C =>
                           regfile_i(18), D => n6290, Z => n2121);
   U2077 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_16_port, C =>
                           regfile_i(19), D => n6290, Z => n2122);
   U2078 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_17_port, C =>
                           regfile_i(20), D => n6290, Z => n2123);
   U2079 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_18_port, C =>
                           regfile_i(21), D => n6290, Z => n2124);
   U2080 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_19_port, C =>
                           regfile_i(22), D => n6290, Z => n2125);
   U2081 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_20_port, C =>
                           regfile_i(23), D => n6290, Z => n2126);
   U2082 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_21_port, C =>
                           regfile_i(24), D => n6290, Z => n2127);
   U2083 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_22_port, C =>
                           regfile_i(25), D => n6290, Z => n2128);
   U2084 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_23_port, C =>
                           regfile_i(26), D => n6290, Z => n2129);
   U2085 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_24_port, C =>
                           regfile_i(27), D => n6290, Z => n2130);
   U2086 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_25_port, C =>
                           regfile_i(28), D => n6290, Z => n2131);
   U2087 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_26_port, C =>
                           regfile_i(29), D => n6290, Z => n2132);
   U2088 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_27_port, C =>
                           regfile_i(30), D => n6290, Z => n2133);
   U2089 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_28_port, C =>
                           regfile_i(31), D => n6290, Z => n2134);
   U2090 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_29_port, C =>
                           regfile_i(32), D => n6290, Z => n2135);
   U2091 : HS65_LH_AO22X9 port map( A => n6287, B => registers_22_30_port, C =>
                           regfile_i(33), D => n6290, Z => n2136);
   U2092 : HS65_LH_AO22X9 port map( A => n6288, B => registers_22_31_port, C =>
                           regfile_i(34), D => n6289, Z => n2137);
   U2093 : HS65_LH_NOR3X4 port map( A => regfile_i(36), B => regfile_i(37), C 
                           => n814, Z => n2837);
   U2094 : HS65_LH_NOR3X4 port map( A => regfile_i(35), B => regfile_i(37), C 
                           => n813, Z => n2835);
   U2095 : HS65_LH_NOR3X4 port map( A => n814, B => regfile_i(37), C => n813, Z
                           => n2833);
   U2096 : HS65_LH_NOR3X4 port map( A => regfile_i(35), B => regfile_i(36), C 
                           => n812, Z => n2831);
   U2097 : HS65_LH_NOR3X4 port map( A => n814, B => regfile_i(36), C => n812, Z
                           => n2829);
   U2098 : HS65_LH_NOR3X4 port map( A => n813, B => regfile_i(35), C => n812, Z
                           => n2827);
   U2099 : HS65_LH_NOR3X4 port map( A => n770, B => regfile_i(49), C => n773, Z
                           => n2805);
   U2100 : HS65_LH_NOR3X4 port map( A => regfile_i(45), B => regfile_i(48), C 
                           => n769, Z => n2822);
   U2101 : HS65_LH_NOR3X4 port map( A => regfile_i(40), B => regfile_i(44), C 
                           => n775, Z => n1324);
   U2102 : HS65_LH_NOR3X4 port map( A => n774, B => regfile_i(43), C => n778, Z
                           => n1331);
   U2103 : HS65_LH_NOR3X4 port map( A => n770, B => regfile_i(45), C => n769, Z
                           => n2809);
   U2104 : HS65_LH_NOR3X4 port map( A => regfile_i(36), B => regfile_i(37), C 
                           => regfile_i(35), Z => n2839);
   U2105 : HS65_LH_NOR3X4 port map( A => regfile_i(40), B => regfile_i(43), C 
                           => n774, Z => n1337);
   U2106 : HS65_LH_NOR3X4 port map( A => regfile_i(43), B => regfile_i(44), C 
                           => n778, Z => n1329);
   U2107 : HS65_LH_NOR3X4 port map( A => n775, B => regfile_i(44), C => n778, Z
                           => n1326);
   U2108 : HS65_LH_NOR3X4 port map( A => regfile_i(48), B => regfile_i(49), C 
                           => n773, Z => n2813);
   U2109 : HS65_LH_NOR3X4 port map( A => regfile_i(45), B => regfile_i(49), C 
                           => n770, Z => n2811);
   U2110 : HS65_LH_NOR3X4 port map( A => n774, B => regfile_i(40), C => n775, Z
                           => n1338);
   U2111 : HS65_LH_NOR3X4 port map( A => n769, B => regfile_i(48), C => n773, Z
                           => n2820);
   U2112 : HS65_LH_NOR2X6 port map( A => regfile_i(46), B => regfile_i(47), Z 
                           => n2807);
   U2113 : HS65_LH_AOI222X2 port map( A => n6508, B => n704, C => 
                           registers_4_0_port, D => n6505, E => 
                           registers_1_0_port, F => n6502, Z => n1319);
   U2114 : HS65_LH_AOI222X2 port map( A => n6508, B => n703, C => 
                           registers_4_1_port, D => n6505, E => 
                           registers_1_1_port, F => n6502, Z => n1165);
   U2115 : HS65_LH_AOI222X2 port map( A => n6509, B => n702, C => 
                           registers_4_2_port, D => n6506, E => 
                           registers_1_2_port, F => n6503, Z => n1011);
   U2116 : HS65_LH_AOI222X2 port map( A => n6510, B => n701, C => 
                           registers_4_3_port, D => n6507, E => 
                           registers_1_3_port, F => n6504, Z => n969);
   U2117 : HS65_LH_AOI222X2 port map( A => n6510, B => n700, C => 
                           registers_4_4_port, D => n6507, E => 
                           registers_1_4_port, F => n6504, Z => n955);
   U2118 : HS65_LH_AOI222X2 port map( A => n6510, B => n699, C => 
                           registers_4_5_port, D => n6507, E => 
                           registers_1_5_port, F => n6504, Z => n941);
   U2119 : HS65_LH_AOI222X2 port map( A => n6510, B => n698, C => 
                           registers_4_6_port, D => n6507, E => 
                           registers_1_6_port, F => n6504, Z => n927);
   U2120 : HS65_LH_AOI222X2 port map( A => n6510, B => n697, C => 
                           registers_4_7_port, D => n6507, E => 
                           registers_1_7_port, F => n6504, Z => n913);
   U2121 : HS65_LH_AOI222X2 port map( A => n6510, B => n696, C => 
                           registers_4_8_port, D => n6507, E => 
                           registers_1_8_port, F => n6504, Z => n899);
   U2122 : HS65_LH_AOI222X2 port map( A => n6510, B => n695, C => 
                           registers_4_9_port, D => n6507, E => 
                           registers_1_9_port, F => n6504, Z => n854);
   U2123 : HS65_LH_AOI222X2 port map( A => n6508, B => n694, C => 
                           registers_4_10_port, D => n6505, E => 
                           registers_1_10_port, F => n6502, Z => n1305);
   U2124 : HS65_LH_AOI222X2 port map( A => n6508, B => n693, C => 
                           registers_4_11_port, D => n6505, E => 
                           registers_1_11_port, F => n6502, Z => n1291);
   U2125 : HS65_LH_AOI222X2 port map( A => n6508, B => n692, C => 
                           registers_4_12_port, D => n6505, E => 
                           registers_1_12_port, F => n6502, Z => n1277);
   U2126 : HS65_LH_AOI222X2 port map( A => n6508, B => n691, C => 
                           registers_4_13_port, D => n6505, E => 
                           registers_1_13_port, F => n6502, Z => n1263);
   U2127 : HS65_LH_AOI222X2 port map( A => n6508, B => n690, C => 
                           registers_4_14_port, D => n6505, E => 
                           registers_1_14_port, F => n6502, Z => n1249);
   U2128 : HS65_LH_AOI222X2 port map( A => n6508, B => n689, C => 
                           registers_4_15_port, D => n6505, E => 
                           registers_1_15_port, F => n6502, Z => n1235);
   U2129 : HS65_LH_AOI222X2 port map( A => n6508, B => n688, C => 
                           registers_4_16_port, D => n6505, E => 
                           registers_1_16_port, F => n6502, Z => n1221);
   U2130 : HS65_LH_AOI222X2 port map( A => n6508, B => n687, C => 
                           registers_4_17_port, D => n6505, E => 
                           registers_1_17_port, F => n6502, Z => n1207);
   U2131 : HS65_LH_AOI222X2 port map( A => n6508, B => n686, C => 
                           registers_4_18_port, D => n6505, E => 
                           registers_1_18_port, F => n6502, Z => n1193);
   U2132 : HS65_LH_AOI222X2 port map( A => n6508, B => n685, C => 
                           registers_4_19_port, D => n6505, E => 
                           registers_1_19_port, F => n6502, Z => n1179);
   U2133 : HS65_LH_AOI222X2 port map( A => n6509, B => n684, C => 
                           registers_4_20_port, D => n6506, E => 
                           registers_1_20_port, F => n6503, Z => n1151);
   U2134 : HS65_LH_AOI222X2 port map( A => n6509, B => n683, C => 
                           registers_4_21_port, D => n6506, E => 
                           registers_1_21_port, F => n6503, Z => n1137);
   U2135 : HS65_LH_AOI222X2 port map( A => n6509, B => n682, C => 
                           registers_4_22_port, D => n6506, E => 
                           registers_1_22_port, F => n6503, Z => n1123);
   U2136 : HS65_LH_AOI222X2 port map( A => n6509, B => n681, C => 
                           registers_4_23_port, D => n6506, E => 
                           registers_1_23_port, F => n6503, Z => n1109);
   U2137 : HS65_LH_AOI222X2 port map( A => n6509, B => n680, C => 
                           registers_4_24_port, D => n6506, E => 
                           registers_1_24_port, F => n6503, Z => n1095);
   U2138 : HS65_LH_AOI222X2 port map( A => n6509, B => n679, C => 
                           registers_4_25_port, D => n6506, E => 
                           registers_1_25_port, F => n6503, Z => n1081);
   U2139 : HS65_LH_AOI222X2 port map( A => n6509, B => n678, C => 
                           registers_4_26_port, D => n6506, E => 
                           registers_1_26_port, F => n6503, Z => n1067);
   U2140 : HS65_LH_AOI222X2 port map( A => n6509, B => n677, C => 
                           registers_4_27_port, D => n6506, E => 
                           registers_1_27_port, F => n6503, Z => n1053);
   U2141 : HS65_LH_AOI222X2 port map( A => n6509, B => n676, C => 
                           registers_4_28_port, D => n6506, E => 
                           registers_1_28_port, F => n6503, Z => n1039);
   U2142 : HS65_LH_AOI222X2 port map( A => n6509, B => n675, C => 
                           registers_4_29_port, D => n6506, E => 
                           registers_1_29_port, F => n6503, Z => n1025);
   U2143 : HS65_LH_AOI222X2 port map( A => n6509, B => n674, C => 
                           registers_4_30_port, D => n6506, E => 
                           registers_1_30_port, F => n6503, Z => n997);
   U2144 : HS65_LH_AOI222X2 port map( A => n6510, B => n673, C => 
                           registers_4_31_port, D => n6507, E => 
                           registers_1_31_port, F => n6504, Z => n983);
   U2145 : HS65_LH_NOR2X6 port map( A => n776, B => regfile_i(41), Z => n1327);
   U2146 : HS65_LH_NOR2X6 port map( A => n772, B => regfile_i(47), Z => n2808);
   U2147 : HS65_LH_NOR2X6 port map( A => regfile_i(41), B => regfile_i(42), Z 
                           => n1328);
   U2148 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_0_port, C 
                           => n6412, D => registers_10_0_port, E => n6409, F =>
                           registers_6_0_port, Z => n2802);
   U2149 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_1_port, C 
                           => n6412, D => registers_10_1_port, E => n6409, F =>
                           registers_6_1_port, Z => n2648);
   U2150 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_2_port, C 
                           => n6413, D => registers_10_2_port, E => n6410, F =>
                           registers_6_2_port, Z => n2494);
   U2151 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_3_port, C 
                           => n6414, D => registers_10_3_port, E => n6410, F =>
                           registers_6_3_port, Z => n2452);
   U2152 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_10_port, C 
                           => n6412, D => registers_10_10_port, E => n6409, F 
                           => registers_6_10_port, Z => n2788);
   U2153 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_11_port, C 
                           => n6412, D => registers_10_11_port, E => n6409, F 
                           => registers_6_11_port, Z => n2774);
   U2154 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_12_port, C 
                           => n6412, D => registers_10_12_port, E => n6409, F 
                           => registers_6_12_port, Z => n2760);
   U2155 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_13_port, C 
                           => n6412, D => registers_10_13_port, E => n6409, F 
                           => registers_6_13_port, Z => n2746);
   U2156 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_14_port, C 
                           => n6412, D => registers_10_14_port, E => n6409, F 
                           => registers_6_14_port, Z => n2732);
   U2157 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_15_port, C 
                           => n6412, D => registers_10_15_port, E => n6409, F 
                           => registers_6_15_port, Z => n2718);
   U2158 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_16_port, C 
                           => n6412, D => registers_10_16_port, E => n6409, F 
                           => registers_6_16_port, Z => n2704);
   U2159 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_17_port, C 
                           => n6412, D => registers_10_17_port, E => n6409, F 
                           => registers_6_17_port, Z => n2690);
   U2160 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_18_port, C 
                           => n6412, D => registers_10_18_port, E => n6409, F 
                           => registers_6_18_port, Z => n2676);
   U2161 : HS65_LH_AOI222X2 port map( A => n6415, B => registers_13_19_port, C 
                           => n6412, D => registers_10_19_port, E => n6409, F 
                           => registers_6_19_port, Z => n2662);
   U2162 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_20_port, C 
                           => n6413, D => registers_10_20_port, E => n6409, F 
                           => registers_6_20_port, Z => n2634);
   U2163 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_21_port, C 
                           => n6413, D => registers_10_21_port, E => n6410, F 
                           => registers_6_21_port, Z => n2620);
   U2164 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_22_port, C 
                           => n6413, D => registers_10_22_port, E => n6410, F 
                           => registers_6_22_port, Z => n2606);
   U2165 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_23_port, C 
                           => n6413, D => registers_10_23_port, E => n6410, F 
                           => registers_6_23_port, Z => n2592);
   U2166 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_24_port, C 
                           => n6413, D => registers_10_24_port, E => n6410, F 
                           => registers_6_24_port, Z => n2578);
   U2167 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_25_port, C 
                           => n6413, D => registers_10_25_port, E => n6410, F 
                           => registers_6_25_port, Z => n2564);
   U2168 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_26_port, C 
                           => n6413, D => registers_10_26_port, E => n6410, F 
                           => registers_6_26_port, Z => n2550);
   U2169 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_27_port, C 
                           => n6413, D => registers_10_27_port, E => n6410, F 
                           => registers_6_27_port, Z => n2536);
   U2170 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_28_port, C 
                           => n6413, D => registers_10_28_port, E => n6410, F 
                           => registers_6_28_port, Z => n2522);
   U2171 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_29_port, C 
                           => n6413, D => registers_10_29_port, E => n6410, F 
                           => registers_6_29_port, Z => n2508);
   U2172 : HS65_LH_AOI222X2 port map( A => n6416, B => registers_13_30_port, C 
                           => n6413, D => registers_10_30_port, E => n6410, F 
                           => registers_6_30_port, Z => n2480);
   U2173 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_31_port, C 
                           => n6414, D => registers_10_31_port, E => n6410, F 
                           => registers_6_31_port, Z => n2466);
   U2174 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_4_port, C 
                           => n6414, D => registers_10_4_port, E => n6411, F =>
                           registers_6_4_port, Z => n2438);
   U2175 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_5_port, C 
                           => n6414, D => registers_10_5_port, E => n6411, F =>
                           registers_6_5_port, Z => n1432);
   U2176 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_6_port, C 
                           => n6414, D => registers_10_6_port, E => n6411, F =>
                           registers_6_6_port, Z => n1418);
   U2177 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_7_port, C 
                           => n6414, D => registers_10_7_port, E => n6411, F =>
                           registers_6_7_port, Z => n1404);
   U2178 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_8_port, C 
                           => n6414, D => registers_10_8_port, E => n6411, F =>
                           registers_6_8_port, Z => n1390);
   U2179 : HS65_LH_AOI222X2 port map( A => n6417, B => registers_13_9_port, C 
                           => n6414, D => registers_10_9_port, E => n6411, F =>
                           registers_6_9_port, Z => n1345);
   U2180 : HS65_LH_NOR2X6 port map( A => n777, B => regfile_i(42), Z => n1325);
   U2181 : HS65_LH_AOI212X4 port map( A => n6463, B => n544, C => 
                           registers_31_0_port, D => n6460, E => n1339, Z => 
                           n1334);
   U2182 : HS65_LH_OAI22X6 port map( A => n6457, B => n288, C => n6454, D => 
                           n448, Z => n1339);
   U2183 : HS65_LH_AOI212X4 port map( A => n6463, B => n543, C => 
                           registers_31_1_port, D => n6460, E => n1173, Z => 
                           n1170);
   U2184 : HS65_LH_OAI22X6 port map( A => n6457, B => n287, C => n6454, D => 
                           n447, Z => n1173);
   U2185 : HS65_LH_AOI212X4 port map( A => n6464, B => n542, C => 
                           registers_31_2_port, D => n6461, E => n1019, Z => 
                           n1016);
   U2186 : HS65_LH_OAI22X6 port map( A => n6458, B => n286, C => n6455, D => 
                           n446, Z => n1019);
   U2187 : HS65_LH_AOI212X4 port map( A => n6464, B => n541, C => 
                           registers_31_3_port, D => n6461, E => n977, Z => 
                           n974);
   U2188 : HS65_LH_OAI22X6 port map( A => n6459, B => n285, C => n6455, D => 
                           n445, Z => n977);
   U2189 : HS65_LH_AOI212X4 port map( A => n6465, B => n540, C => 
                           registers_31_4_port, D => n6462, E => n963, Z => 
                           n960);
   U2190 : HS65_LH_OAI22X6 port map( A => n6459, B => n284, C => n6456, D => 
                           n444, Z => n963);
   U2191 : HS65_LH_AOI212X4 port map( A => n6465, B => n539, C => 
                           registers_31_5_port, D => n6462, E => n949, Z => 
                           n946);
   U2192 : HS65_LH_OAI22X6 port map( A => n6459, B => n283, C => n6456, D => 
                           n443, Z => n949);
   U2193 : HS65_LH_AOI212X4 port map( A => n6465, B => n538, C => 
                           registers_31_6_port, D => n6462, E => n935, Z => 
                           n932);
   U2194 : HS65_LH_OAI22X6 port map( A => n6459, B => n282, C => n6456, D => 
                           n442, Z => n935);
   U2195 : HS65_LH_AOI212X4 port map( A => n6465, B => n537, C => 
                           registers_31_7_port, D => n6462, E => n921, Z => 
                           n918);
   U2196 : HS65_LH_OAI22X6 port map( A => n6459, B => n281, C => n6456, D => 
                           n441, Z => n921);
   U2197 : HS65_LH_AOI212X4 port map( A => n6465, B => n536, C => 
                           registers_31_8_port, D => n6462, E => n907, Z => 
                           n904);
   U2198 : HS65_LH_OAI22X6 port map( A => n6459, B => n280, C => n6456, D => 
                           n440, Z => n907);
   U2199 : HS65_LH_AOI212X4 port map( A => n6465, B => n535, C => 
                           registers_31_9_port, D => n6462, E => n883, Z => 
                           n874);
   U2200 : HS65_LH_OAI22X6 port map( A => n6459, B => n279, C => n6456, D => 
                           n439, Z => n883);
   U2201 : HS65_LH_AOI212X4 port map( A => n6463, B => n534, C => 
                           registers_31_10_port, D => n6460, E => n1313, Z => 
                           n1310);
   U2202 : HS65_LH_OAI22X6 port map( A => n6457, B => n278, C => n6454, D => 
                           n438, Z => n1313);
   U2203 : HS65_LH_AOI212X4 port map( A => n6463, B => n533, C => 
                           registers_31_11_port, D => n6460, E => n1299, Z => 
                           n1296);
   U2204 : HS65_LH_OAI22X6 port map( A => n6457, B => n277, C => n6454, D => 
                           n437, Z => n1299);
   U2205 : HS65_LH_AOI212X4 port map( A => n6463, B => n532, C => 
                           registers_31_12_port, D => n6460, E => n1285, Z => 
                           n1282);
   U2206 : HS65_LH_OAI22X6 port map( A => n6457, B => n276, C => n6454, D => 
                           n436, Z => n1285);
   U2207 : HS65_LH_AOI212X4 port map( A => n6463, B => n531, C => 
                           registers_31_13_port, D => n6460, E => n1271, Z => 
                           n1268);
   U2208 : HS65_LH_OAI22X6 port map( A => n6457, B => n275, C => n6454, D => 
                           n435, Z => n1271);
   U2209 : HS65_LH_AOI212X4 port map( A => n6463, B => n530, C => 
                           registers_31_14_port, D => n6460, E => n1257, Z => 
                           n1254);
   U2210 : HS65_LH_OAI22X6 port map( A => n6457, B => n274, C => n6454, D => 
                           n434, Z => n1257);
   U2211 : HS65_LH_AOI212X4 port map( A => n6463, B => n529, C => 
                           registers_31_15_port, D => n6460, E => n1243, Z => 
                           n1240);
   U2212 : HS65_LH_OAI22X6 port map( A => n6457, B => n273, C => n6454, D => 
                           n433, Z => n1243);
   U2213 : HS65_LH_AOI212X4 port map( A => n6463, B => n528, C => 
                           registers_31_16_port, D => n6460, E => n1229, Z => 
                           n1226);
   U2214 : HS65_LH_OAI22X6 port map( A => n6457, B => n272, C => n6454, D => 
                           n432, Z => n1229);
   U2215 : HS65_LH_AOI212X4 port map( A => n6463, B => n527, C => 
                           registers_31_17_port, D => n6460, E => n1215, Z => 
                           n1212);
   U2216 : HS65_LH_OAI22X6 port map( A => n6457, B => n271, C => n6454, D => 
                           n431, Z => n1215);
   U2217 : HS65_LH_AOI212X4 port map( A => n6463, B => n526, C => 
                           registers_31_18_port, D => n6460, E => n1201, Z => 
                           n1198);
   U2218 : HS65_LH_OAI22X6 port map( A => n6457, B => n270, C => n6454, D => 
                           n430, Z => n1201);
   U2219 : HS65_LH_AOI212X4 port map( A => n6463, B => n525, C => 
                           registers_31_19_port, D => n6460, E => n1187, Z => 
                           n1184);
   U2220 : HS65_LH_OAI22X6 port map( A => n6457, B => n269, C => n6454, D => 
                           n429, Z => n1187);
   U2221 : HS65_LH_AOI212X4 port map( A => n6463, B => n524, C => 
                           registers_31_20_port, D => n6460, E => n1159, Z => 
                           n1156);
   U2222 : HS65_LH_OAI22X6 port map( A => n6458, B => n268, C => n6454, D => 
                           n428, Z => n1159);
   U2223 : HS65_LH_AOI212X4 port map( A => n6464, B => n523, C => 
                           registers_31_21_port, D => n6461, E => n1145, Z => 
                           n1142);
   U2224 : HS65_LH_OAI22X6 port map( A => n6458, B => n267, C => n6455, D => 
                           n427, Z => n1145);
   U2225 : HS65_LH_AOI212X4 port map( A => n6464, B => n522, C => 
                           registers_31_22_port, D => n6461, E => n1131, Z => 
                           n1128);
   U2226 : HS65_LH_OAI22X6 port map( A => n6458, B => n266, C => n6455, D => 
                           n426, Z => n1131);
   U2227 : HS65_LH_AOI212X4 port map( A => n6464, B => n521, C => 
                           registers_31_23_port, D => n6461, E => n1117, Z => 
                           n1114);
   U2228 : HS65_LH_OAI22X6 port map( A => n6458, B => n265, C => n6455, D => 
                           n425, Z => n1117);
   U2229 : HS65_LH_AOI212X4 port map( A => n6464, B => n520, C => 
                           registers_31_24_port, D => n6461, E => n1103, Z => 
                           n1100);
   U2230 : HS65_LH_OAI22X6 port map( A => n6458, B => n264, C => n6455, D => 
                           n424, Z => n1103);
   U2231 : HS65_LH_AOI212X4 port map( A => n6464, B => n519, C => 
                           registers_31_25_port, D => n6461, E => n1089, Z => 
                           n1086);
   U2232 : HS65_LH_OAI22X6 port map( A => n6458, B => n263, C => n6455, D => 
                           n423, Z => n1089);
   U2233 : HS65_LH_AOI212X4 port map( A => n6464, B => n518, C => 
                           registers_31_26_port, D => n6461, E => n1075, Z => 
                           n1072);
   U2234 : HS65_LH_OAI22X6 port map( A => n6458, B => n262, C => n6455, D => 
                           n422, Z => n1075);
   U2235 : HS65_LH_AOI212X4 port map( A => n6464, B => n517, C => 
                           registers_31_27_port, D => n6461, E => n1061, Z => 
                           n1058);
   U2236 : HS65_LH_OAI22X6 port map( A => n6458, B => n261, C => n6455, D => 
                           n421, Z => n1061);
   U2237 : HS65_LH_AOI212X4 port map( A => n6464, B => n516, C => 
                           registers_31_28_port, D => n6461, E => n1047, Z => 
                           n1044);
   U2238 : HS65_LH_OAI22X6 port map( A => n6458, B => n260, C => n6455, D => 
                           n420, Z => n1047);
   U2239 : HS65_LH_AOI212X4 port map( A => n6464, B => n515, C => 
                           registers_31_29_port, D => n6461, E => n1033, Z => 
                           n1030);
   U2240 : HS65_LH_OAI22X6 port map( A => n6458, B => n259, C => n6455, D => 
                           n419, Z => n1033);
   U2241 : HS65_LH_AOI212X4 port map( A => n6464, B => n514, C => 
                           registers_31_30_port, D => n6461, E => n1005, Z => 
                           n1002);
   U2242 : HS65_LH_OAI22X6 port map( A => n6458, B => n258, C => n6455, D => 
                           n418, Z => n1005);
   U2243 : HS65_LH_AOI212X4 port map( A => n6464, B => n513, C => 
                           registers_31_31_port, D => n6461, E => n991, Z => 
                           n988);
   U2244 : HS65_LH_OAI22X6 port map( A => n6459, B => n257, C => n6455, D => 
                           n417, Z => n991);
   U2245 : HS65_LH_AOI212X4 port map( A => n6520, B => n736, C => 
                           registers_13_0_port, D => n6517, E => n1321, Z => 
                           n1320);
   U2246 : HS65_LH_IVX9 port map( A => n224, Z => n736);
   U2247 : HS65_LH_OAI22X6 port map( A => n6514, B => n480, C => n6511, D => 
                           n512, Z => n1321);
   U2248 : HS65_LH_AOI212X4 port map( A => n6520, B => n735, C => 
                           registers_13_1_port, D => n6517, E => n1167, Z => 
                           n1166);
   U2249 : HS65_LH_IVX9 port map( A => n223, Z => n735);
   U2250 : HS65_LH_OAI22X6 port map( A => n6514, B => n479, C => n6511, D => 
                           n511, Z => n1167);
   U2251 : HS65_LH_AOI212X4 port map( A => n6521, B => n734, C => 
                           registers_13_2_port, D => n6518, E => n1013, Z => 
                           n1012);
   U2252 : HS65_LH_IVX9 port map( A => n222, Z => n734);
   U2253 : HS65_LH_OAI22X6 port map( A => n6515, B => n478, C => n6512, D => 
                           n510, Z => n1013);
   U2254 : HS65_LH_AOI212X4 port map( A => n6521, B => n733, C => 
                           registers_13_3_port, D => n6518, E => n971, Z => 
                           n970);
   U2255 : HS65_LH_IVX9 port map( A => n221, Z => n733);
   U2256 : HS65_LH_OAI22X6 port map( A => n6516, B => n477, C => n6512, D => 
                           n509, Z => n971);
   U2257 : HS65_LH_AOI212X4 port map( A => n6522, B => n732, C => 
                           registers_13_4_port, D => n6519, E => n957, Z => 
                           n956);
   U2258 : HS65_LH_IVX9 port map( A => n220, Z => n732);
   U2259 : HS65_LH_OAI22X6 port map( A => n6516, B => n476, C => n6513, D => 
                           n508, Z => n957);
   U2260 : HS65_LH_AOI212X4 port map( A => n6522, B => n731, C => 
                           registers_13_5_port, D => n6519, E => n943, Z => 
                           n942);
   U2261 : HS65_LH_IVX9 port map( A => n219, Z => n731);
   U2262 : HS65_LH_OAI22X6 port map( A => n6516, B => n475, C => n6513, D => 
                           n507, Z => n943);
   U2263 : HS65_LH_AOI212X4 port map( A => n6522, B => n730, C => 
                           registers_13_6_port, D => n6519, E => n929, Z => 
                           n928);
   U2264 : HS65_LH_IVX9 port map( A => n218, Z => n730);
   U2265 : HS65_LH_OAI22X6 port map( A => n6516, B => n474, C => n6513, D => 
                           n506, Z => n929);
   U2266 : HS65_LH_AOI212X4 port map( A => n6522, B => n729, C => 
                           registers_13_7_port, D => n6519, E => n915, Z => 
                           n914);
   U2267 : HS65_LH_IVX9 port map( A => n217, Z => n729);
   U2268 : HS65_LH_OAI22X6 port map( A => n6516, B => n473, C => n6513, D => 
                           n505, Z => n915);
   U2269 : HS65_LH_AOI212X4 port map( A => n6522, B => n728, C => 
                           registers_13_8_port, D => n6519, E => n901, Z => 
                           n900);
   U2270 : HS65_LH_IVX9 port map( A => n216, Z => n728);
   U2271 : HS65_LH_OAI22X6 port map( A => n6516, B => n472, C => n6513, D => 
                           n504, Z => n901);
   U2272 : HS65_LH_AOI212X4 port map( A => n6522, B => n727, C => 
                           registers_13_9_port, D => n6519, E => n858, Z => 
                           n855);
   U2273 : HS65_LH_IVX9 port map( A => n215, Z => n727);
   U2274 : HS65_LH_OAI22X6 port map( A => n6516, B => n471, C => n6513, D => 
                           n503, Z => n858);
   U2275 : HS65_LH_AOI212X4 port map( A => n6520, B => n726, C => 
                           registers_13_10_port, D => n6517, E => n1307, Z => 
                           n1306);
   U2276 : HS65_LH_IVX9 port map( A => n214, Z => n726);
   U2277 : HS65_LH_OAI22X6 port map( A => n6514, B => n470, C => n6511, D => 
                           n502, Z => n1307);
   U2278 : HS65_LH_AOI212X4 port map( A => n6520, B => n725, C => 
                           registers_13_11_port, D => n6517, E => n1293, Z => 
                           n1292);
   U2279 : HS65_LH_IVX9 port map( A => n213, Z => n725);
   U2280 : HS65_LH_OAI22X6 port map( A => n6514, B => n469, C => n6511, D => 
                           n501, Z => n1293);
   U2281 : HS65_LH_AOI212X4 port map( A => n6520, B => n724, C => 
                           registers_13_12_port, D => n6517, E => n1279, Z => 
                           n1278);
   U2282 : HS65_LH_IVX9 port map( A => n212, Z => n724);
   U2283 : HS65_LH_OAI22X6 port map( A => n6514, B => n468, C => n6511, D => 
                           n500, Z => n1279);
   U2284 : HS65_LH_AOI212X4 port map( A => n6520, B => n723, C => 
                           registers_13_13_port, D => n6517, E => n1265, Z => 
                           n1264);
   U2285 : HS65_LH_IVX9 port map( A => n211, Z => n723);
   U2286 : HS65_LH_OAI22X6 port map( A => n6514, B => n467, C => n6511, D => 
                           n499, Z => n1265);
   U2287 : HS65_LH_AOI212X4 port map( A => n6520, B => n722, C => 
                           registers_13_14_port, D => n6517, E => n1251, Z => 
                           n1250);
   U2288 : HS65_LH_IVX9 port map( A => n210, Z => n722);
   U2289 : HS65_LH_OAI22X6 port map( A => n6514, B => n466, C => n6511, D => 
                           n498, Z => n1251);
   U2290 : HS65_LH_AOI212X4 port map( A => n6520, B => n721, C => 
                           registers_13_15_port, D => n6517, E => n1237, Z => 
                           n1236);
   U2291 : HS65_LH_IVX9 port map( A => n209, Z => n721);
   U2292 : HS65_LH_OAI22X6 port map( A => n6514, B => n465, C => n6511, D => 
                           n497, Z => n1237);
   U2293 : HS65_LH_AOI212X4 port map( A => n6520, B => n720, C => 
                           registers_13_16_port, D => n6517, E => n1223, Z => 
                           n1222);
   U2294 : HS65_LH_IVX9 port map( A => n208, Z => n720);
   U2295 : HS65_LH_OAI22X6 port map( A => n6514, B => n464, C => n6511, D => 
                           n496, Z => n1223);
   U2296 : HS65_LH_AOI212X4 port map( A => n6520, B => n719, C => 
                           registers_13_17_port, D => n6517, E => n1209, Z => 
                           n1208);
   U2297 : HS65_LH_IVX9 port map( A => n207, Z => n719);
   U2298 : HS65_LH_OAI22X6 port map( A => n6514, B => n463, C => n6511, D => 
                           n495, Z => n1209);
   U2299 : HS65_LH_AOI212X4 port map( A => n6520, B => n718, C => 
                           registers_13_18_port, D => n6517, E => n1195, Z => 
                           n1194);
   U2300 : HS65_LH_IVX9 port map( A => n206, Z => n718);
   U2301 : HS65_LH_OAI22X6 port map( A => n6514, B => n462, C => n6511, D => 
                           n494, Z => n1195);
   U2302 : HS65_LH_AOI212X4 port map( A => n6520, B => n717, C => 
                           registers_13_19_port, D => n6517, E => n1181, Z => 
                           n1180);
   U2303 : HS65_LH_IVX9 port map( A => n205, Z => n717);
   U2304 : HS65_LH_OAI22X6 port map( A => n6514, B => n461, C => n6511, D => 
                           n493, Z => n1181);
   U2305 : HS65_LH_AOI212X4 port map( A => n6520, B => n716, C => 
                           registers_13_20_port, D => n6517, E => n1153, Z => 
                           n1152);
   U2306 : HS65_LH_IVX9 port map( A => n204, Z => n716);
   U2307 : HS65_LH_OAI22X6 port map( A => n6515, B => n460, C => n6511, D => 
                           n492, Z => n1153);
   U2308 : HS65_LH_AOI212X4 port map( A => n6521, B => n715, C => 
                           registers_13_21_port, D => n6518, E => n1139, Z => 
                           n1138);
   U2309 : HS65_LH_IVX9 port map( A => n203, Z => n715);
   U2310 : HS65_LH_OAI22X6 port map( A => n6515, B => n459, C => n6512, D => 
                           n491, Z => n1139);
   U2311 : HS65_LH_AOI212X4 port map( A => n6521, B => n714, C => 
                           registers_13_22_port, D => n6518, E => n1125, Z => 
                           n1124);
   U2312 : HS65_LH_IVX9 port map( A => n202, Z => n714);
   U2313 : HS65_LH_OAI22X6 port map( A => n6515, B => n458, C => n6512, D => 
                           n490, Z => n1125);
   U2314 : HS65_LH_AOI212X4 port map( A => n6521, B => n713, C => 
                           registers_13_23_port, D => n6518, E => n1111, Z => 
                           n1110);
   U2315 : HS65_LH_IVX9 port map( A => n201, Z => n713);
   U2316 : HS65_LH_OAI22X6 port map( A => n6515, B => n457, C => n6512, D => 
                           n489, Z => n1111);
   U2317 : HS65_LH_AOI212X4 port map( A => n6521, B => n712, C => 
                           registers_13_24_port, D => n6518, E => n1097, Z => 
                           n1096);
   U2318 : HS65_LH_IVX9 port map( A => n200, Z => n712);
   U2319 : HS65_LH_OAI22X6 port map( A => n6515, B => n456, C => n6512, D => 
                           n488, Z => n1097);
   U2320 : HS65_LH_AOI212X4 port map( A => n6521, B => n711, C => 
                           registers_13_25_port, D => n6518, E => n1083, Z => 
                           n1082);
   U2321 : HS65_LH_IVX9 port map( A => n199, Z => n711);
   U2322 : HS65_LH_OAI22X6 port map( A => n6515, B => n455, C => n6512, D => 
                           n487, Z => n1083);
   U2323 : HS65_LH_AOI212X4 port map( A => n6521, B => n710, C => 
                           registers_13_26_port, D => n6518, E => n1069, Z => 
                           n1068);
   U2324 : HS65_LH_IVX9 port map( A => n198, Z => n710);
   U2325 : HS65_LH_OAI22X6 port map( A => n6515, B => n454, C => n6512, D => 
                           n486, Z => n1069);
   U2326 : HS65_LH_AOI212X4 port map( A => n6521, B => n709, C => 
                           registers_13_27_port, D => n6518, E => n1055, Z => 
                           n1054);
   U2327 : HS65_LH_IVX9 port map( A => n197, Z => n709);
   U2328 : HS65_LH_OAI22X6 port map( A => n6515, B => n453, C => n6512, D => 
                           n485, Z => n1055);
   U2329 : HS65_LH_AOI212X4 port map( A => n6521, B => n708, C => 
                           registers_13_28_port, D => n6518, E => n1041, Z => 
                           n1040);
   U2330 : HS65_LH_IVX9 port map( A => n196, Z => n708);
   U2331 : HS65_LH_OAI22X6 port map( A => n6515, B => n452, C => n6512, D => 
                           n484, Z => n1041);
   U2332 : HS65_LH_AOI212X4 port map( A => n6521, B => n707, C => 
                           registers_13_29_port, D => n6518, E => n1027, Z => 
                           n1026);
   U2333 : HS65_LH_IVX9 port map( A => n195, Z => n707);
   U2334 : HS65_LH_OAI22X6 port map( A => n6515, B => n451, C => n6512, D => 
                           n483, Z => n1027);
   U2335 : HS65_LH_AOI212X4 port map( A => n6521, B => n706, C => 
                           registers_13_30_port, D => n6518, E => n999, Z => 
                           n998);
   U2336 : HS65_LH_IVX9 port map( A => n194, Z => n706);
   U2337 : HS65_LH_OAI22X6 port map( A => n6515, B => n450, C => n6512, D => 
                           n482, Z => n999);
   U2338 : HS65_LH_AOI212X4 port map( A => n6521, B => n705, C => 
                           registers_13_31_port, D => n6518, E => n985, Z => 
                           n984);
   U2339 : HS65_LH_IVX9 port map( A => n193, Z => n705);
   U2340 : HS65_LH_OAI22X6 port map( A => n6516, B => n449, C => n6512, D => 
                           n481, Z => n985);
   U2341 : HS65_LH_NOR3X4 port map( A => regfile_i(43), B => regfile_i(44), C 
                           => regfile_i(40), Z => n1322);
   U2342 : HS65_LH_AOI212X4 port map( A => registers_18_0_port, B => n6475, C 
                           => registers_24_0_port, D => n6472, E => n1336, Z =>
                           n1335);
   U2343 : HS65_LH_OAI22X6 port map( A => n6469, B => n416, C => n6466, D => 
                           n384, Z => n1336);
   U2344 : HS65_LH_AOI212X4 port map( A => registers_18_1_port, B => n6475, C 
                           => registers_24_1_port, D => n6472, E => n1172, Z =>
                           n1171);
   U2345 : HS65_LH_OAI22X6 port map( A => n6469, B => n415, C => n6466, D => 
                           n383, Z => n1172);
   U2346 : HS65_LH_AOI212X4 port map( A => registers_18_2_port, B => n6476, C 
                           => registers_24_2_port, D => n6473, E => n1018, Z =>
                           n1017);
   U2347 : HS65_LH_OAI22X6 port map( A => n6470, B => n414, C => n6467, D => 
                           n382, Z => n1018);
   U2348 : HS65_LH_AOI212X4 port map( A => registers_18_3_port, B => n6477, C 
                           => registers_24_3_port, D => n6473, E => n976, Z => 
                           n975);
   U2349 : HS65_LH_OAI22X6 port map( A => n6471, B => n413, C => n6467, D => 
                           n381, Z => n976);
   U2350 : HS65_LH_AOI212X4 port map( A => registers_18_4_port, B => n6477, C 
                           => registers_24_4_port, D => n6474, E => n962, Z => 
                           n961);
   U2351 : HS65_LH_OAI22X6 port map( A => n6471, B => n412, C => n6468, D => 
                           n380, Z => n962);
   U2352 : HS65_LH_AOI212X4 port map( A => registers_18_5_port, B => n6477, C 
                           => registers_24_5_port, D => n6474, E => n948, Z => 
                           n947);
   U2353 : HS65_LH_OAI22X6 port map( A => n6471, B => n411, C => n6468, D => 
                           n379, Z => n948);
   U2354 : HS65_LH_AOI212X4 port map( A => registers_18_6_port, B => n6477, C 
                           => registers_24_6_port, D => n6474, E => n934, Z => 
                           n933);
   U2355 : HS65_LH_OAI22X6 port map( A => n6471, B => n410, C => n6468, D => 
                           n378, Z => n934);
   U2356 : HS65_LH_AOI212X4 port map( A => registers_18_7_port, B => n6477, C 
                           => registers_24_7_port, D => n6474, E => n920, Z => 
                           n919);
   U2357 : HS65_LH_OAI22X6 port map( A => n6471, B => n409, C => n6468, D => 
                           n377, Z => n920);
   U2358 : HS65_LH_AOI212X4 port map( A => registers_18_8_port, B => n6477, C 
                           => registers_24_8_port, D => n6474, E => n906, Z => 
                           n905);
   U2359 : HS65_LH_OAI22X6 port map( A => n6471, B => n408, C => n6468, D => 
                           n376, Z => n906);
   U2360 : HS65_LH_AOI212X4 port map( A => registers_18_9_port, B => n6477, C 
                           => registers_24_9_port, D => n6474, E => n878, Z => 
                           n875);
   U2361 : HS65_LH_OAI22X6 port map( A => n6471, B => n407, C => n6468, D => 
                           n375, Z => n878);
   U2362 : HS65_LH_AOI212X4 port map( A => registers_18_11_port, B => n6475, C 
                           => registers_24_11_port, D => n6472, E => n1298, Z 
                           => n1297);
   U2363 : HS65_LH_OAI22X6 port map( A => n6469, B => n405, C => n6466, D => 
                           n373, Z => n1298);
   U2364 : HS65_LH_AOI212X4 port map( A => registers_18_12_port, B => n6475, C 
                           => registers_24_12_port, D => n6472, E => n1284, Z 
                           => n1283);
   U2365 : HS65_LH_OAI22X6 port map( A => n6469, B => n404, C => n6466, D => 
                           n372, Z => n1284);
   U2366 : HS65_LH_AOI212X4 port map( A => registers_18_13_port, B => n6475, C 
                           => registers_24_13_port, D => n6472, E => n1270, Z 
                           => n1269);
   U2367 : HS65_LH_OAI22X6 port map( A => n6469, B => n403, C => n6466, D => 
                           n371, Z => n1270);
   U2368 : HS65_LH_AOI212X4 port map( A => registers_18_14_port, B => n6475, C 
                           => registers_24_14_port, D => n6472, E => n1256, Z 
                           => n1255);
   U2369 : HS65_LH_OAI22X6 port map( A => n6469, B => n402, C => n6466, D => 
                           n370, Z => n1256);
   U2370 : HS65_LH_AOI212X4 port map( A => registers_18_15_port, B => n6475, C 
                           => registers_24_15_port, D => n6472, E => n1242, Z 
                           => n1241);
   U2371 : HS65_LH_OAI22X6 port map( A => n6469, B => n401, C => n6466, D => 
                           n369, Z => n1242);
   U2372 : HS65_LH_AOI212X4 port map( A => registers_18_16_port, B => n6475, C 
                           => registers_24_16_port, D => n6472, E => n1228, Z 
                           => n1227);
   U2373 : HS65_LH_OAI22X6 port map( A => n6469, B => n400, C => n6466, D => 
                           n368, Z => n1228);
   U2374 : HS65_LH_AOI212X4 port map( A => registers_18_17_port, B => n6475, C 
                           => registers_24_17_port, D => n6472, E => n1214, Z 
                           => n1213);
   U2375 : HS65_LH_OAI22X6 port map( A => n6469, B => n399, C => n6466, D => 
                           n367, Z => n1214);
   U2376 : HS65_LH_AOI212X4 port map( A => registers_18_18_port, B => n6475, C 
                           => registers_24_18_port, D => n6472, E => n1200, Z 
                           => n1199);
   U2377 : HS65_LH_OAI22X6 port map( A => n6469, B => n398, C => n6466, D => 
                           n366, Z => n1200);
   U2378 : HS65_LH_AOI212X4 port map( A => registers_18_19_port, B => n6475, C 
                           => registers_24_19_port, D => n6472, E => n1186, Z 
                           => n1185);
   U2379 : HS65_LH_OAI22X6 port map( A => n6469, B => n397, C => n6466, D => 
                           n365, Z => n1186);
   U2380 : HS65_LH_AOI212X4 port map( A => registers_18_20_port, B => n6476, C 
                           => registers_24_20_port, D => n6472, E => n1158, Z 
                           => n1157);
   U2381 : HS65_LH_OAI22X6 port map( A => n6470, B => n396, C => n6466, D => 
                           n364, Z => n1158);
   U2382 : HS65_LH_AOI212X4 port map( A => registers_18_21_port, B => n6476, C 
                           => registers_24_21_port, D => n6473, E => n1144, Z 
                           => n1143);
   U2383 : HS65_LH_OAI22X6 port map( A => n6470, B => n395, C => n6467, D => 
                           n363, Z => n1144);
   U2384 : HS65_LH_AOI212X4 port map( A => registers_18_22_port, B => n6476, C 
                           => registers_24_22_port, D => n6473, E => n1130, Z 
                           => n1129);
   U2385 : HS65_LH_OAI22X6 port map( A => n6470, B => n394, C => n6467, D => 
                           n362, Z => n1130);
   U2386 : HS65_LH_AOI212X4 port map( A => registers_18_23_port, B => n6476, C 
                           => registers_24_23_port, D => n6473, E => n1116, Z 
                           => n1115);
   U2387 : HS65_LH_OAI22X6 port map( A => n6470, B => n393, C => n6467, D => 
                           n361, Z => n1116);
   U2388 : HS65_LH_AOI212X4 port map( A => registers_18_24_port, B => n6476, C 
                           => registers_24_24_port, D => n6473, E => n1102, Z 
                           => n1101);
   U2389 : HS65_LH_OAI22X6 port map( A => n6470, B => n392, C => n6467, D => 
                           n360, Z => n1102);
   U2390 : HS65_LH_AOI212X4 port map( A => registers_18_25_port, B => n6476, C 
                           => registers_24_25_port, D => n6473, E => n1088, Z 
                           => n1087);
   U2391 : HS65_LH_OAI22X6 port map( A => n6470, B => n391, C => n6467, D => 
                           n359, Z => n1088);
   U2392 : HS65_LH_AOI212X4 port map( A => registers_18_26_port, B => n6476, C 
                           => registers_24_26_port, D => n6473, E => n1074, Z 
                           => n1073);
   U2393 : HS65_LH_OAI22X6 port map( A => n6470, B => n390, C => n6467, D => 
                           n358, Z => n1074);
   U2394 : HS65_LH_AOI212X4 port map( A => registers_18_27_port, B => n6476, C 
                           => registers_24_27_port, D => n6473, E => n1060, Z 
                           => n1059);
   U2395 : HS65_LH_OAI22X6 port map( A => n6470, B => n389, C => n6467, D => 
                           n357, Z => n1060);
   U2396 : HS65_LH_AOI212X4 port map( A => registers_18_28_port, B => n6476, C 
                           => registers_24_28_port, D => n6473, E => n1046, Z 
                           => n1045);
   U2397 : HS65_LH_OAI22X6 port map( A => n6470, B => n388, C => n6467, D => 
                           n356, Z => n1046);
   U2398 : HS65_LH_AOI212X4 port map( A => registers_18_29_port, B => n6476, C 
                           => registers_24_29_port, D => n6473, E => n1032, Z 
                           => n1031);
   U2399 : HS65_LH_OAI22X6 port map( A => n6470, B => n387, C => n6467, D => 
                           n355, Z => n1032);
   U2400 : HS65_LH_AOI212X4 port map( A => registers_18_30_port, B => n6476, C 
                           => registers_24_30_port, D => n6473, E => n1004, Z 
                           => n1003);
   U2401 : HS65_LH_OAI22X6 port map( A => n6470, B => n386, C => n6467, D => 
                           n354, Z => n1004);
   U2402 : HS65_LH_AOI212X4 port map( A => registers_18_31_port, B => n6477, C 
                           => registers_24_31_port, D => n6473, E => n990, Z =>
                           n989);
   U2403 : HS65_LH_OAI22X6 port map( A => n6471, B => n385, C => n6467, D => 
                           n353, Z => n990);
   U2404 : HS65_LH_NOR2X6 port map( A => n771, B => regfile_i(46), Z => n2812);
   U2405 : HS65_LH_AOI212X4 port map( A => n6370, B => n544, C => n6367, D => 
                           registers_31_0_port, E => n2821, Z => n2816);
   U2406 : HS65_LH_OAI22X6 port map( A => n416, B => n6364, C => n352, D => 
                           n6361, Z => n2821);
   U2407 : HS65_LH_AOI212X4 port map( A => n6370, B => n543, C => n6367, D => 
                           registers_31_1_port, E => n2656, Z => n2653);
   U2408 : HS65_LH_OAI22X6 port map( A => n415, B => n6364, C => n351, D => 
                           n6361, Z => n2656);
   U2409 : HS65_LH_AOI212X4 port map( A => n6371, B => n542, C => n6368, D => 
                           registers_31_2_port, E => n2502, Z => n2499);
   U2410 : HS65_LH_OAI22X6 port map( A => n414, B => n6365, C => n350, D => 
                           n6362, Z => n2502);
   U2411 : HS65_LH_AOI212X4 port map( A => n6371, B => n541, C => n6368, D => 
                           registers_31_3_port, E => n2460, Z => n2457);
   U2412 : HS65_LH_OAI22X6 port map( A => n413, B => n6366, C => n349, D => 
                           n6362, Z => n2460);
   U2413 : HS65_LH_AOI212X4 port map( A => n6370, B => n534, C => n6367, D => 
                           registers_31_10_port, E => n2796, Z => n2793);
   U2414 : HS65_LH_OAI22X6 port map( A => n406, B => n6364, C => n342, D => 
                           n6361, Z => n2796);
   U2415 : HS65_LH_AOI212X4 port map( A => n6370, B => n533, C => n6367, D => 
                           registers_31_11_port, E => n2782, Z => n2779);
   U2416 : HS65_LH_OAI22X6 port map( A => n405, B => n6364, C => n341, D => 
                           n6361, Z => n2782);
   U2417 : HS65_LH_AOI212X4 port map( A => n6370, B => n532, C => n6367, D => 
                           registers_31_12_port, E => n2768, Z => n2765);
   U2418 : HS65_LH_OAI22X6 port map( A => n404, B => n6364, C => n340, D => 
                           n6361, Z => n2768);
   U2419 : HS65_LH_AOI212X4 port map( A => n6370, B => n531, C => n6367, D => 
                           registers_31_13_port, E => n2754, Z => n2751);
   U2420 : HS65_LH_OAI22X6 port map( A => n403, B => n6364, C => n339, D => 
                           n6361, Z => n2754);
   U2421 : HS65_LH_AOI212X4 port map( A => n6370, B => n530, C => n6367, D => 
                           registers_31_14_port, E => n2740, Z => n2737);
   U2422 : HS65_LH_OAI22X6 port map( A => n402, B => n6364, C => n338, D => 
                           n6361, Z => n2740);
   U2423 : HS65_LH_AOI212X4 port map( A => n6370, B => n529, C => n6367, D => 
                           registers_31_15_port, E => n2726, Z => n2723);
   U2424 : HS65_LH_OAI22X6 port map( A => n401, B => n6364, C => n337, D => 
                           n6361, Z => n2726);
   U2425 : HS65_LH_AOI212X4 port map( A => n6370, B => n528, C => n6367, D => 
                           registers_31_16_port, E => n2712, Z => n2709);
   U2426 : HS65_LH_OAI22X6 port map( A => n400, B => n6364, C => n336, D => 
                           n6361, Z => n2712);
   U2427 : HS65_LH_AOI212X4 port map( A => n6370, B => n527, C => n6367, D => 
                           registers_31_17_port, E => n2698, Z => n2695);
   U2428 : HS65_LH_OAI22X6 port map( A => n399, B => n6364, C => n335, D => 
                           n6361, Z => n2698);
   U2429 : HS65_LH_AOI212X4 port map( A => n6370, B => n526, C => n6367, D => 
                           registers_31_18_port, E => n2684, Z => n2681);
   U2430 : HS65_LH_OAI22X6 port map( A => n398, B => n6364, C => n334, D => 
                           n6361, Z => n2684);
   U2431 : HS65_LH_AOI212X4 port map( A => n6370, B => n525, C => n6367, D => 
                           registers_31_19_port, E => n2670, Z => n2667);
   U2432 : HS65_LH_OAI22X6 port map( A => n397, B => n6364, C => n333, D => 
                           n6361, Z => n2670);
   U2433 : HS65_LH_AOI212X4 port map( A => n6370, B => n524, C => n6367, D => 
                           registers_31_20_port, E => n2642, Z => n2639);
   U2434 : HS65_LH_OAI22X6 port map( A => n396, B => n6365, C => n332, D => 
                           n6361, Z => n2642);
   U2435 : HS65_LH_AOI212X4 port map( A => n6371, B => n523, C => n6368, D => 
                           registers_31_21_port, E => n2628, Z => n2625);
   U2436 : HS65_LH_OAI22X6 port map( A => n395, B => n6365, C => n331, D => 
                           n6362, Z => n2628);
   U2437 : HS65_LH_AOI212X4 port map( A => n6371, B => n522, C => n6368, D => 
                           registers_31_22_port, E => n2614, Z => n2611);
   U2438 : HS65_LH_OAI22X6 port map( A => n394, B => n6365, C => n330, D => 
                           n6362, Z => n2614);
   U2439 : HS65_LH_AOI212X4 port map( A => n6371, B => n521, C => n6368, D => 
                           registers_31_23_port, E => n2600, Z => n2597);
   U2440 : HS65_LH_OAI22X6 port map( A => n393, B => n6365, C => n329, D => 
                           n6362, Z => n2600);
   U2441 : HS65_LH_AOI212X4 port map( A => n6371, B => n520, C => n6368, D => 
                           registers_31_24_port, E => n2586, Z => n2583);
   U2442 : HS65_LH_OAI22X6 port map( A => n392, B => n6365, C => n328, D => 
                           n6362, Z => n2586);
   U2443 : HS65_LH_AOI212X4 port map( A => n6371, B => n519, C => n6368, D => 
                           registers_31_25_port, E => n2572, Z => n2569);
   U2444 : HS65_LH_OAI22X6 port map( A => n391, B => n6365, C => n327, D => 
                           n6362, Z => n2572);
   U2445 : HS65_LH_AOI212X4 port map( A => n6371, B => n518, C => n6368, D => 
                           registers_31_26_port, E => n2558, Z => n2555);
   U2446 : HS65_LH_OAI22X6 port map( A => n390, B => n6365, C => n326, D => 
                           n6362, Z => n2558);
   U2447 : HS65_LH_AOI212X4 port map( A => n6371, B => n517, C => n6368, D => 
                           registers_31_27_port, E => n2544, Z => n2541);
   U2448 : HS65_LH_OAI22X6 port map( A => n389, B => n6365, C => n325, D => 
                           n6362, Z => n2544);
   U2449 : HS65_LH_AOI212X4 port map( A => n6371, B => n516, C => n6368, D => 
                           registers_31_28_port, E => n2530, Z => n2527);
   U2450 : HS65_LH_OAI22X6 port map( A => n388, B => n6365, C => n324, D => 
                           n6362, Z => n2530);
   U2451 : HS65_LH_AOI212X4 port map( A => n6371, B => n515, C => n6368, D => 
                           registers_31_29_port, E => n2516, Z => n2513);
   U2452 : HS65_LH_OAI22X6 port map( A => n387, B => n6365, C => n323, D => 
                           n6362, Z => n2516);
   U2453 : HS65_LH_AOI212X4 port map( A => n6371, B => n514, C => n6368, D => 
                           registers_31_30_port, E => n2488, Z => n2485);
   U2454 : HS65_LH_OAI22X6 port map( A => n386, B => n6365, C => n322, D => 
                           n6362, Z => n2488);
   U2455 : HS65_LH_AOI212X4 port map( A => n6371, B => n513, C => n6368, D => 
                           registers_31_31_port, E => n2474, Z => n2471);
   U2456 : HS65_LH_OAI22X6 port map( A => n385, B => n6366, C => n321, D => 
                           n6362, Z => n2474);
   U2457 : HS65_LH_AOI212X4 port map( A => n6372, B => n540, C => n6369, D => 
                           registers_31_4_port, E => n2446, Z => n2443);
   U2458 : HS65_LH_OAI22X6 port map( A => n412, B => n6366, C => n348, D => 
                           n6363, Z => n2446);
   U2459 : HS65_LH_AOI212X4 port map( A => n6372, B => n539, C => n6369, D => 
                           registers_31_5_port, E => n2432, Z => n2429);
   U2460 : HS65_LH_OAI22X6 port map( A => n411, B => n6366, C => n347, D => 
                           n6363, Z => n2432);
   U2461 : HS65_LH_AOI212X4 port map( A => n6372, B => n538, C => n6369, D => 
                           registers_31_6_port, E => n1426, Z => n1423);
   U2462 : HS65_LH_OAI22X6 port map( A => n410, B => n6366, C => n346, D => 
                           n6363, Z => n1426);
   U2463 : HS65_LH_AOI212X4 port map( A => n6372, B => n537, C => n6369, D => 
                           registers_31_7_port, E => n1412, Z => n1409);
   U2464 : HS65_LH_OAI22X6 port map( A => n409, B => n6366, C => n345, D => 
                           n6363, Z => n1412);
   U2465 : HS65_LH_AOI212X4 port map( A => n6372, B => n536, C => n6369, D => 
                           registers_31_8_port, E => n1398, Z => n1395);
   U2466 : HS65_LH_OAI22X6 port map( A => n408, B => n6366, C => n344, D => 
                           n6363, Z => n1398);
   U2467 : HS65_LH_AOI212X4 port map( A => n6372, B => n535, C => n6369, D => 
                           registers_31_9_port, E => n1374, Z => n1365);
   U2468 : HS65_LH_OAI22X6 port map( A => n407, B => n6366, C => n343, D => 
                           n6363, Z => n1374);
   U2469 : HS65_LH_AOI212X4 port map( A => n6427, B => n672, C => n6424, D => 
                           registers_11_0_port, E => n2804, Z => n2803);
   U2470 : HS65_LH_OAI22X6 port map( A => n224, B => n6421, C => n160, D => 
                           n6418, Z => n2804);
   U2471 : HS65_LH_AOI212X4 port map( A => n6427, B => n671, C => n6424, D => 
                           registers_11_1_port, E => n2650, Z => n2649);
   U2472 : HS65_LH_OAI22X6 port map( A => n223, B => n6421, C => n159, D => 
                           n6418, Z => n2650);
   U2473 : HS65_LH_AOI212X4 port map( A => n6428, B => n670, C => n6425, D => 
                           registers_11_2_port, E => n2496, Z => n2495);
   U2474 : HS65_LH_OAI22X6 port map( A => n222, B => n6422, C => n158, D => 
                           n6419, Z => n2496);
   U2475 : HS65_LH_AOI212X4 port map( A => n6428, B => n669, C => n6425, D => 
                           registers_11_3_port, E => n2454, Z => n2453);
   U2476 : HS65_LH_OAI22X6 port map( A => n221, B => n6423, C => n157, D => 
                           n6419, Z => n2454);
   U2477 : HS65_LH_AOI212X4 port map( A => n6429, B => n668, C => n6426, D => 
                           registers_11_4_port, E => n2440, Z => n2439);
   U2478 : HS65_LH_OAI22X6 port map( A => n220, B => n6423, C => n156, D => 
                           n6420, Z => n2440);
   U2479 : HS65_LH_AOI212X4 port map( A => n6429, B => n667, C => n6426, D => 
                           registers_11_5_port, E => n2426, Z => n1433);
   U2480 : HS65_LH_OAI22X6 port map( A => n219, B => n6423, C => n155, D => 
                           n6420, Z => n2426);
   U2481 : HS65_LH_AOI212X4 port map( A => n6429, B => n666, C => n6426, D => 
                           registers_11_6_port, E => n1420, Z => n1419);
   U2482 : HS65_LH_OAI22X6 port map( A => n218, B => n6423, C => n154, D => 
                           n6420, Z => n1420);
   U2483 : HS65_LH_AOI212X4 port map( A => n6429, B => n665, C => n6426, D => 
                           registers_11_7_port, E => n1406, Z => n1405);
   U2484 : HS65_LH_OAI22X6 port map( A => n217, B => n6423, C => n153, D => 
                           n6420, Z => n1406);
   U2485 : HS65_LH_AOI212X4 port map( A => n6429, B => n664, C => n6426, D => 
                           registers_11_8_port, E => n1392, Z => n1391);
   U2486 : HS65_LH_OAI22X6 port map( A => n216, B => n6423, C => n152, D => 
                           n6420, Z => n1392);
   U2487 : HS65_LH_AOI212X4 port map( A => n6429, B => n663, C => n6426, D => 
                           registers_11_9_port, E => n1349, Z => n1346);
   U2488 : HS65_LH_OAI22X6 port map( A => n215, B => n6423, C => n151, D => 
                           n6420, Z => n1349);
   U2489 : HS65_LH_AOI212X4 port map( A => n6427, B => n662, C => n6424, D => 
                           registers_11_10_port, E => n2790, Z => n2789);
   U2490 : HS65_LH_OAI22X6 port map( A => n214, B => n6421, C => n150, D => 
                           n6418, Z => n2790);
   U2491 : HS65_LH_AOI212X4 port map( A => n6427, B => n661, C => n6424, D => 
                           registers_11_11_port, E => n2776, Z => n2775);
   U2492 : HS65_LH_OAI22X6 port map( A => n213, B => n6421, C => n149, D => 
                           n6418, Z => n2776);
   U2493 : HS65_LH_AOI212X4 port map( A => n6427, B => n660, C => n6424, D => 
                           registers_11_12_port, E => n2762, Z => n2761);
   U2494 : HS65_LH_OAI22X6 port map( A => n212, B => n6421, C => n148, D => 
                           n6418, Z => n2762);
   U2495 : HS65_LH_AOI212X4 port map( A => n6427, B => n659, C => n6424, D => 
                           registers_11_13_port, E => n2748, Z => n2747);
   U2496 : HS65_LH_OAI22X6 port map( A => n211, B => n6421, C => n147, D => 
                           n6418, Z => n2748);
   U2497 : HS65_LH_AOI212X4 port map( A => n6427, B => n658, C => n6424, D => 
                           registers_11_14_port, E => n2734, Z => n2733);
   U2498 : HS65_LH_OAI22X6 port map( A => n210, B => n6421, C => n146, D => 
                           n6418, Z => n2734);
   U2499 : HS65_LH_AOI212X4 port map( A => n6427, B => n657, C => n6424, D => 
                           registers_11_15_port, E => n2720, Z => n2719);
   U2500 : HS65_LH_OAI22X6 port map( A => n209, B => n6421, C => n145, D => 
                           n6418, Z => n2720);
   U2501 : HS65_LH_AOI212X4 port map( A => n6427, B => n656, C => n6424, D => 
                           registers_11_16_port, E => n2706, Z => n2705);
   U2502 : HS65_LH_OAI22X6 port map( A => n208, B => n6421, C => n144, D => 
                           n6418, Z => n2706);
   U2503 : HS65_LH_AOI212X4 port map( A => n6427, B => n655, C => n6424, D => 
                           registers_11_17_port, E => n2692, Z => n2691);
   U2504 : HS65_LH_OAI22X6 port map( A => n207, B => n6421, C => n143, D => 
                           n6418, Z => n2692);
   U2505 : HS65_LH_AOI212X4 port map( A => n6427, B => n654, C => n6424, D => 
                           registers_11_18_port, E => n2678, Z => n2677);
   U2506 : HS65_LH_OAI22X6 port map( A => n206, B => n6421, C => n142, D => 
                           n6418, Z => n2678);
   U2507 : HS65_LH_AOI212X4 port map( A => n6427, B => n653, C => n6424, D => 
                           registers_11_19_port, E => n2664, Z => n2663);
   U2508 : HS65_LH_OAI22X6 port map( A => n205, B => n6421, C => n141, D => 
                           n6418, Z => n2664);
   U2509 : HS65_LH_AOI212X4 port map( A => n6427, B => n652, C => n6424, D => 
                           registers_11_20_port, E => n2636, Z => n2635);
   U2510 : HS65_LH_OAI22X6 port map( A => n204, B => n6422, C => n140, D => 
                           n6418, Z => n2636);
   U2511 : HS65_LH_AOI212X4 port map( A => n6428, B => n651, C => n6425, D => 
                           registers_11_21_port, E => n2622, Z => n2621);
   U2512 : HS65_LH_OAI22X6 port map( A => n203, B => n6422, C => n139, D => 
                           n6419, Z => n2622);
   U2513 : HS65_LH_AOI212X4 port map( A => n6428, B => n650, C => n6425, D => 
                           registers_11_22_port, E => n2608, Z => n2607);
   U2514 : HS65_LH_OAI22X6 port map( A => n202, B => n6422, C => n138, D => 
                           n6419, Z => n2608);
   U2515 : HS65_LH_AOI212X4 port map( A => n6428, B => n649, C => n6425, D => 
                           registers_11_23_port, E => n2594, Z => n2593);
   U2516 : HS65_LH_OAI22X6 port map( A => n201, B => n6422, C => n137, D => 
                           n6419, Z => n2594);
   U2517 : HS65_LH_AOI212X4 port map( A => n6428, B => n648, C => n6425, D => 
                           registers_11_24_port, E => n2580, Z => n2579);
   U2518 : HS65_LH_OAI22X6 port map( A => n200, B => n6422, C => n136, D => 
                           n6419, Z => n2580);
   U2519 : HS65_LH_AOI212X4 port map( A => n6428, B => n647, C => n6425, D => 
                           registers_11_25_port, E => n2566, Z => n2565);
   U2520 : HS65_LH_OAI22X6 port map( A => n199, B => n6422, C => n135, D => 
                           n6419, Z => n2566);
   U2521 : HS65_LH_AOI212X4 port map( A => n6428, B => n646, C => n6425, D => 
                           registers_11_26_port, E => n2552, Z => n2551);
   U2522 : HS65_LH_OAI22X6 port map( A => n198, B => n6422, C => n134, D => 
                           n6419, Z => n2552);
   U2523 : HS65_LH_AOI212X4 port map( A => n6428, B => n645, C => n6425, D => 
                           registers_11_27_port, E => n2538, Z => n2537);
   U2524 : HS65_LH_OAI22X6 port map( A => n197, B => n6422, C => n133, D => 
                           n6419, Z => n2538);
   U2525 : HS65_LH_AOI212X4 port map( A => n6428, B => n644, C => n6425, D => 
                           registers_11_28_port, E => n2524, Z => n2523);
   U2526 : HS65_LH_OAI22X6 port map( A => n196, B => n6422, C => n132, D => 
                           n6419, Z => n2524);
   U2527 : HS65_LH_AOI212X4 port map( A => n6428, B => n643, C => n6425, D => 
                           registers_11_29_port, E => n2510, Z => n2509);
   U2528 : HS65_LH_OAI22X6 port map( A => n195, B => n6422, C => n131, D => 
                           n6419, Z => n2510);
   U2529 : HS65_LH_AOI212X4 port map( A => n6428, B => n642, C => n6425, D => 
                           registers_11_30_port, E => n2482, Z => n2481);
   U2530 : HS65_LH_OAI22X6 port map( A => n194, B => n6422, C => n130, D => 
                           n6419, Z => n2482);
   U2531 : HS65_LH_AOI212X4 port map( A => n6428, B => n641, C => n6425, D => 
                           registers_11_31_port, E => n2468, Z => n2467);
   U2532 : HS65_LH_OAI22X6 port map( A => n193, B => n6423, C => n129, D => 
                           n6419, Z => n2468);
   U2533 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_0_port, C 
                           => n6379, D => registers_19_0_port, E => n2818, Z =>
                           n2817);
   U2534 : HS65_LH_OAI22X6 port map( A => n288, B => n6376, C => n320, D => 
                           n6373, Z => n2818);
   U2535 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_1_port, C 
                           => n6379, D => registers_19_1_port, E => n2655, Z =>
                           n2654);
   U2536 : HS65_LH_OAI22X6 port map( A => n287, B => n6376, C => n319, D => 
                           n6373, Z => n2655);
   U2537 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_2_port, C 
                           => n6380, D => registers_19_2_port, E => n2501, Z =>
                           n2500);
   U2538 : HS65_LH_OAI22X6 port map( A => n286, B => n6377, C => n318, D => 
                           n6374, Z => n2501);
   U2539 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_3_port, C 
                           => n6380, D => registers_19_3_port, E => n2459, Z =>
                           n2458);
   U2540 : HS65_LH_OAI22X6 port map( A => n285, B => n6378, C => n317, D => 
                           n6374, Z => n2459);
   U2541 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_10_port, C 
                           => n6379, D => registers_19_10_port, E => n2795, Z 
                           => n2794);
   U2542 : HS65_LH_OAI22X6 port map( A => n278, B => n6376, C => n310, D => 
                           n6373, Z => n2795);
   U2543 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_11_port, C 
                           => n6379, D => registers_19_11_port, E => n2781, Z 
                           => n2780);
   U2544 : HS65_LH_OAI22X6 port map( A => n277, B => n6376, C => n309, D => 
                           n6373, Z => n2781);
   U2545 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_12_port, C 
                           => n6379, D => registers_19_12_port, E => n2767, Z 
                           => n2766);
   U2546 : HS65_LH_OAI22X6 port map( A => n276, B => n6376, C => n308, D => 
                           n6373, Z => n2767);
   U2547 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_13_port, C 
                           => n6379, D => registers_19_13_port, E => n2753, Z 
                           => n2752);
   U2548 : HS65_LH_OAI22X6 port map( A => n275, B => n6376, C => n307, D => 
                           n6373, Z => n2753);
   U2549 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_14_port, C 
                           => n6379, D => registers_19_14_port, E => n2739, Z 
                           => n2738);
   U2550 : HS65_LH_OAI22X6 port map( A => n274, B => n6376, C => n306, D => 
                           n6373, Z => n2739);
   U2551 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_15_port, C 
                           => n6379, D => registers_19_15_port, E => n2725, Z 
                           => n2724);
   U2552 : HS65_LH_OAI22X6 port map( A => n273, B => n6376, C => n305, D => 
                           n6373, Z => n2725);
   U2553 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_16_port, C 
                           => n6379, D => registers_19_16_port, E => n2711, Z 
                           => n2710);
   U2554 : HS65_LH_OAI22X6 port map( A => n272, B => n6376, C => n304, D => 
                           n6373, Z => n2711);
   U2555 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_17_port, C 
                           => n6379, D => registers_19_17_port, E => n2697, Z 
                           => n2696);
   U2556 : HS65_LH_OAI22X6 port map( A => n271, B => n6376, C => n303, D => 
                           n6373, Z => n2697);
   U2557 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_18_port, C 
                           => n6379, D => registers_19_18_port, E => n2683, Z 
                           => n2682);
   U2558 : HS65_LH_OAI22X6 port map( A => n270, B => n6376, C => n302, D => 
                           n6373, Z => n2683);
   U2559 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_19_port, C 
                           => n6379, D => registers_19_19_port, E => n2669, Z 
                           => n2668);
   U2560 : HS65_LH_OAI22X6 port map( A => n269, B => n6376, C => n301, D => 
                           n6373, Z => n2669);
   U2561 : HS65_LH_AOI212X4 port map( A => n6382, B => registers_17_20_port, C 
                           => n6379, D => registers_19_20_port, E => n2641, Z 
                           => n2640);
   U2562 : HS65_LH_OAI22X6 port map( A => n268, B => n6377, C => n300, D => 
                           n6373, Z => n2641);
   U2563 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_21_port, C 
                           => n6380, D => registers_19_21_port, E => n2627, Z 
                           => n2626);
   U2564 : HS65_LH_OAI22X6 port map( A => n267, B => n6377, C => n299, D => 
                           n6374, Z => n2627);
   U2565 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_22_port, C 
                           => n6380, D => registers_19_22_port, E => n2613, Z 
                           => n2612);
   U2566 : HS65_LH_OAI22X6 port map( A => n266, B => n6377, C => n298, D => 
                           n6374, Z => n2613);
   U2567 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_23_port, C 
                           => n6380, D => registers_19_23_port, E => n2599, Z 
                           => n2598);
   U2568 : HS65_LH_OAI22X6 port map( A => n265, B => n6377, C => n297, D => 
                           n6374, Z => n2599);
   U2569 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_24_port, C 
                           => n6380, D => registers_19_24_port, E => n2585, Z 
                           => n2584);
   U2570 : HS65_LH_OAI22X6 port map( A => n264, B => n6377, C => n296, D => 
                           n6374, Z => n2585);
   U2571 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_25_port, C 
                           => n6380, D => registers_19_25_port, E => n2571, Z 
                           => n2570);
   U2572 : HS65_LH_OAI22X6 port map( A => n263, B => n6377, C => n295, D => 
                           n6374, Z => n2571);
   U2573 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_26_port, C 
                           => n6380, D => registers_19_26_port, E => n2557, Z 
                           => n2556);
   U2574 : HS65_LH_OAI22X6 port map( A => n262, B => n6377, C => n294, D => 
                           n6374, Z => n2557);
   U2575 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_27_port, C 
                           => n6380, D => registers_19_27_port, E => n2543, Z 
                           => n2542);
   U2576 : HS65_LH_OAI22X6 port map( A => n261, B => n6377, C => n293, D => 
                           n6374, Z => n2543);
   U2577 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_28_port, C 
                           => n6380, D => registers_19_28_port, E => n2529, Z 
                           => n2528);
   U2578 : HS65_LH_OAI22X6 port map( A => n260, B => n6377, C => n292, D => 
                           n6374, Z => n2529);
   U2579 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_29_port, C 
                           => n6380, D => registers_19_29_port, E => n2515, Z 
                           => n2514);
   U2580 : HS65_LH_OAI22X6 port map( A => n259, B => n6377, C => n291, D => 
                           n6374, Z => n2515);
   U2581 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_30_port, C 
                           => n6380, D => registers_19_30_port, E => n2487, Z 
                           => n2486);
   U2582 : HS65_LH_OAI22X6 port map( A => n258, B => n6377, C => n290, D => 
                           n6374, Z => n2487);
   U2583 : HS65_LH_AOI212X4 port map( A => n6383, B => registers_17_31_port, C 
                           => n6380, D => registers_19_31_port, E => n2473, Z 
                           => n2472);
   U2584 : HS65_LH_OAI22X6 port map( A => n257, B => n6378, C => n289, D => 
                           n6374, Z => n2473);
   U2585 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_4_port, C 
                           => n6381, D => registers_19_4_port, E => n2445, Z =>
                           n2444);
   U2586 : HS65_LH_OAI22X6 port map( A => n284, B => n6378, C => n316, D => 
                           n6375, Z => n2445);
   U2587 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_5_port, C 
                           => n6381, D => registers_19_5_port, E => n2431, Z =>
                           n2430);
   U2588 : HS65_LH_OAI22X6 port map( A => n283, B => n6378, C => n315, D => 
                           n6375, Z => n2431);
   U2589 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_6_port, C 
                           => n6381, D => registers_19_6_port, E => n1425, Z =>
                           n1424);
   U2590 : HS65_LH_OAI22X6 port map( A => n282, B => n6378, C => n314, D => 
                           n6375, Z => n1425);
   U2591 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_7_port, C 
                           => n6381, D => registers_19_7_port, E => n1411, Z =>
                           n1410);
   U2592 : HS65_LH_OAI22X6 port map( A => n281, B => n6378, C => n313, D => 
                           n6375, Z => n1411);
   U2593 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_8_port, C 
                           => n6381, D => registers_19_8_port, E => n1397, Z =>
                           n1396);
   U2594 : HS65_LH_OAI22X6 port map( A => n280, B => n6378, C => n312, D => 
                           n6375, Z => n1397);
   U2595 : HS65_LH_AOI212X4 port map( A => n6384, B => registers_17_9_port, C 
                           => n6381, D => registers_19_9_port, E => n1369, Z =>
                           n1366);
   U2596 : HS65_LH_OAI22X6 port map( A => n279, B => n6378, C => n311, D => 
                           n6375, Z => n1369);
   U2597 : HS65_LH_NOR3X4 port map( A => regfile_i(48), B => regfile_i(49), C 
                           => regfile_i(45), Z => n2810);
   U2598 : HS65_LH_NAND4ABX3 port map( A => n1308, B => n1309, C => n1310, D =>
                           n1311, Z => n1301);
   U2599 : HS65_LH_MX41X7 port map( D0 => registers_22_10_port, S0 => n6439, D1
                           => registers_21_10_port, S1 => n6436, D2 => 
                           registers_19_10_port, S2 => n6433, D3 => n6430, S3 
                           => n598, Z => n1308);
   U2600 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n758, D1 => 
                           registers_30_10_port, S1 => n6448, D2 => n6445, S2 
                           => n662, D3 => registers_20_10_port, S3 => n6442, Z 
                           => n1309);
   U2601 : HS65_LH_AOI212X4 port map( A => registers_18_10_port, B => n6475, C 
                           => registers_24_10_port, D => n6472, E => n1312, Z 
                           => n1311);
   U2602 : HS65_LH_IVX9 port map( A => regfile_i(44), Z => n774);
   U2603 : HS65_LH_IVX9 port map( A => regfile_i(48), Z => n770);
   U2604 : HS65_LH_IVX9 port map( A => regfile_i(35), Z => n814);
   U2605 : HS65_LH_IVX9 port map( A => regfile_i(43), Z => n775);
   U2606 : HS65_LH_IVX9 port map( A => regfile_i(49), Z => n769);
   U2607 : HS65_LH_IVX9 port map( A => regfile_i(36), Z => n813);
   U2608 : HS65_LH_MX41X7 port map( D0 => registers_5_0_port, S0 => n6487, D1 
                           => registers_11_0_port, S1 => n6484, D2 => 
                           registers_7_0_port, S2 => n6481, D3 => 
                           registers_3_0_port, S3 => n6478, Z => n1317);
   U2609 : HS65_LH_MX41X7 port map( D0 => registers_5_1_port, S0 => n6487, D1 
                           => registers_11_1_port, S1 => n6484, D2 => 
                           registers_7_1_port, S2 => n6481, D3 => 
                           registers_3_1_port, S3 => n6478, Z => n1163);
   U2610 : HS65_LH_MX41X7 port map( D0 => registers_5_2_port, S0 => n6488, D1 
                           => registers_11_2_port, S1 => n6485, D2 => 
                           registers_7_2_port, S2 => n6482, D3 => 
                           registers_3_2_port, S3 => n6479, Z => n1009);
   U2611 : HS65_LH_MX41X7 port map( D0 => registers_5_3_port, S0 => n6489, D1 
                           => registers_11_3_port, S1 => n6486, D2 => 
                           registers_7_3_port, S2 => n6483, D3 => 
                           registers_3_3_port, S3 => n6480, Z => n967);
   U2612 : HS65_LH_MX41X7 port map( D0 => registers_5_4_port, S0 => n6489, D1 
                           => registers_11_4_port, S1 => n6486, D2 => 
                           registers_7_4_port, S2 => n6483, D3 => 
                           registers_3_4_port, S3 => n6480, Z => n953);
   U2613 : HS65_LH_MX41X7 port map( D0 => registers_5_5_port, S0 => n6489, D1 
                           => registers_11_5_port, S1 => n6486, D2 => 
                           registers_7_5_port, S2 => n6483, D3 => 
                           registers_3_5_port, S3 => n6480, Z => n939);
   U2614 : HS65_LH_MX41X7 port map( D0 => registers_5_6_port, S0 => n6489, D1 
                           => registers_11_6_port, S1 => n6486, D2 => 
                           registers_7_6_port, S2 => n6483, D3 => 
                           registers_3_6_port, S3 => n6480, Z => n925);
   U2615 : HS65_LH_MX41X7 port map( D0 => registers_5_7_port, S0 => n6489, D1 
                           => registers_11_7_port, S1 => n6486, D2 => 
                           registers_7_7_port, S2 => n6483, D3 => 
                           registers_3_7_port, S3 => n6480, Z => n911);
   U2616 : HS65_LH_MX41X7 port map( D0 => registers_5_8_port, S0 => n6489, D1 
                           => registers_11_8_port, S1 => n6486, D2 => 
                           registers_7_8_port, S2 => n6483, D3 => 
                           registers_3_8_port, S3 => n6480, Z => n897);
   U2617 : HS65_LH_MX41X7 port map( D0 => registers_5_9_port, S0 => n6489, D1 
                           => registers_11_9_port, S1 => n6486, D2 => 
                           registers_7_9_port, S2 => n6483, D3 => 
                           registers_3_9_port, S3 => n6480, Z => n852);
   U2618 : HS65_LH_MX41X7 port map( D0 => registers_5_10_port, S0 => n6487, D1 
                           => registers_11_10_port, S1 => n6484, D2 => 
                           registers_7_10_port, S2 => n6481, D3 => 
                           registers_3_10_port, S3 => n6478, Z => n1303);
   U2619 : HS65_LH_MX41X7 port map( D0 => registers_5_11_port, S0 => n6487, D1 
                           => registers_11_11_port, S1 => n6484, D2 => 
                           registers_7_11_port, S2 => n6481, D3 => 
                           registers_3_11_port, S3 => n6478, Z => n1289);
   U2620 : HS65_LH_MX41X7 port map( D0 => registers_5_12_port, S0 => n6487, D1 
                           => registers_11_12_port, S1 => n6484, D2 => 
                           registers_7_12_port, S2 => n6481, D3 => 
                           registers_3_12_port, S3 => n6478, Z => n1275);
   U2621 : HS65_LH_MX41X7 port map( D0 => registers_5_13_port, S0 => n6487, D1 
                           => registers_11_13_port, S1 => n6484, D2 => 
                           registers_7_13_port, S2 => n6481, D3 => 
                           registers_3_13_port, S3 => n6478, Z => n1261);
   U2622 : HS65_LH_MX41X7 port map( D0 => registers_5_14_port, S0 => n6487, D1 
                           => registers_11_14_port, S1 => n6484, D2 => 
                           registers_7_14_port, S2 => n6481, D3 => 
                           registers_3_14_port, S3 => n6478, Z => n1247);
   U2623 : HS65_LH_MX41X7 port map( D0 => registers_5_15_port, S0 => n6487, D1 
                           => registers_11_15_port, S1 => n6484, D2 => 
                           registers_7_15_port, S2 => n6481, D3 => 
                           registers_3_15_port, S3 => n6478, Z => n1233);
   U2624 : HS65_LH_MX41X7 port map( D0 => registers_5_16_port, S0 => n6487, D1 
                           => registers_11_16_port, S1 => n6484, D2 => 
                           registers_7_16_port, S2 => n6481, D3 => 
                           registers_3_16_port, S3 => n6478, Z => n1219);
   U2625 : HS65_LH_MX41X7 port map( D0 => registers_5_17_port, S0 => n6487, D1 
                           => registers_11_17_port, S1 => n6484, D2 => 
                           registers_7_17_port, S2 => n6481, D3 => 
                           registers_3_17_port, S3 => n6478, Z => n1205);
   U2626 : HS65_LH_MX41X7 port map( D0 => registers_5_18_port, S0 => n6487, D1 
                           => registers_11_18_port, S1 => n6484, D2 => 
                           registers_7_18_port, S2 => n6481, D3 => 
                           registers_3_18_port, S3 => n6478, Z => n1191);
   U2627 : HS65_LH_MX41X7 port map( D0 => registers_5_19_port, S0 => n6487, D1 
                           => registers_11_19_port, S1 => n6484, D2 => 
                           registers_7_19_port, S2 => n6481, D3 => 
                           registers_3_19_port, S3 => n6478, Z => n1177);
   U2628 : HS65_LH_MX41X7 port map( D0 => registers_5_20_port, S0 => n6488, D1 
                           => registers_11_20_port, S1 => n6485, D2 => 
                           registers_7_20_port, S2 => n6482, D3 => 
                           registers_3_20_port, S3 => n6479, Z => n1149);
   U2629 : HS65_LH_MX41X7 port map( D0 => registers_5_21_port, S0 => n6488, D1 
                           => registers_11_21_port, S1 => n6485, D2 => 
                           registers_7_21_port, S2 => n6482, D3 => 
                           registers_3_21_port, S3 => n6479, Z => n1135);
   U2630 : HS65_LH_MX41X7 port map( D0 => registers_5_22_port, S0 => n6488, D1 
                           => registers_11_22_port, S1 => n6485, D2 => 
                           registers_7_22_port, S2 => n6482, D3 => 
                           registers_3_22_port, S3 => n6479, Z => n1121);
   U2631 : HS65_LH_MX41X7 port map( D0 => registers_5_23_port, S0 => n6488, D1 
                           => registers_11_23_port, S1 => n6485, D2 => 
                           registers_7_23_port, S2 => n6482, D3 => 
                           registers_3_23_port, S3 => n6479, Z => n1107);
   U2632 : HS65_LH_MX41X7 port map( D0 => registers_5_24_port, S0 => n6488, D1 
                           => registers_11_24_port, S1 => n6485, D2 => 
                           registers_7_24_port, S2 => n6482, D3 => 
                           registers_3_24_port, S3 => n6479, Z => n1093);
   U2633 : HS65_LH_MX41X7 port map( D0 => registers_5_25_port, S0 => n6488, D1 
                           => registers_11_25_port, S1 => n6485, D2 => 
                           registers_7_25_port, S2 => n6482, D3 => 
                           registers_3_25_port, S3 => n6479, Z => n1079);
   U2634 : HS65_LH_MX41X7 port map( D0 => registers_5_26_port, S0 => n6488, D1 
                           => registers_11_26_port, S1 => n6485, D2 => 
                           registers_7_26_port, S2 => n6482, D3 => 
                           registers_3_26_port, S3 => n6479, Z => n1065);
   U2635 : HS65_LH_MX41X7 port map( D0 => registers_5_27_port, S0 => n6488, D1 
                           => registers_11_27_port, S1 => n6485, D2 => 
                           registers_7_27_port, S2 => n6482, D3 => 
                           registers_3_27_port, S3 => n6479, Z => n1051);
   U2636 : HS65_LH_MX41X7 port map( D0 => registers_5_28_port, S0 => n6488, D1 
                           => registers_11_28_port, S1 => n6485, D2 => 
                           registers_7_28_port, S2 => n6482, D3 => 
                           registers_3_28_port, S3 => n6479, Z => n1037);
   U2637 : HS65_LH_MX41X7 port map( D0 => registers_5_29_port, S0 => n6488, D1 
                           => registers_11_29_port, S1 => n6485, D2 => 
                           registers_7_29_port, S2 => n6482, D3 => 
                           registers_3_29_port, S3 => n6479, Z => n1023);
   U2638 : HS65_LH_MX41X7 port map( D0 => registers_5_30_port, S0 => n6488, D1 
                           => registers_11_30_port, S1 => n6485, D2 => 
                           registers_7_30_port, S2 => n6482, D3 => 
                           registers_3_30_port, S3 => n6479, Z => n995);
   U2639 : HS65_LH_MX41X7 port map( D0 => registers_5_31_port, S0 => n6489, D1 
                           => registers_11_31_port, S1 => n6486, D2 => 
                           registers_7_31_port, S2 => n6483, D3 => 
                           registers_3_31_port, S3 => n6480, Z => n981);
   U2640 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n768, D1 => 
                           registers_30_0_port, S1 => n6448, D2 => n6445, S2 =>
                           n672, D3 => registers_20_0_port, S3 => n6442, Z => 
                           n1333);
   U2641 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n767, D1 => 
                           registers_30_1_port, S1 => n6448, D2 => n6445, S2 =>
                           n671, D3 => registers_20_1_port, S3 => n6442, Z => 
                           n1169);
   U2642 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n766, D1 => 
                           registers_30_2_port, S1 => n6449, D2 => n6446, S2 =>
                           n670, D3 => registers_20_2_port, S3 => n6443, Z => 
                           n1015);
   U2643 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n765, D1 => 
                           registers_30_3_port, S1 => n6450, D2 => n6446, S2 =>
                           n669, D3 => registers_20_3_port, S3 => n6444, Z => 
                           n973);
   U2644 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n764, D1 => 
                           registers_30_4_port, S1 => n6450, D2 => n6447, S2 =>
                           n668, D3 => registers_20_4_port, S3 => n6444, Z => 
                           n959);
   U2645 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n763, D1 => 
                           registers_30_5_port, S1 => n6450, D2 => n6447, S2 =>
                           n667, D3 => registers_20_5_port, S3 => n6444, Z => 
                           n945);
   U2646 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n762, D1 => 
                           registers_30_6_port, S1 => n6450, D2 => n6447, S2 =>
                           n666, D3 => registers_20_6_port, S3 => n6444, Z => 
                           n931);
   U2647 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n761, D1 => 
                           registers_30_7_port, S1 => n6450, D2 => n6447, S2 =>
                           n665, D3 => registers_20_7_port, S3 => n6444, Z => 
                           n917);
   U2648 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n760, D1 => 
                           registers_30_8_port, S1 => n6450, D2 => n6447, S2 =>
                           n664, D3 => registers_20_8_port, S3 => n6444, Z => 
                           n903);
   U2649 : HS65_LH_MX41X7 port map( D0 => n6453, S0 => n759, D1 => 
                           registers_30_9_port, S1 => n6450, D2 => n6447, S2 =>
                           n663, D3 => registers_20_9_port, S3 => n6444, Z => 
                           n873);
   U2650 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n757, D1 => 
                           registers_30_11_port, S1 => n6448, D2 => n6445, S2 
                           => n661, D3 => registers_20_11_port, S3 => n6442, Z 
                           => n1295);
   U2651 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n756, D1 => 
                           registers_30_12_port, S1 => n6448, D2 => n6445, S2 
                           => n660, D3 => registers_20_12_port, S3 => n6442, Z 
                           => n1281);
   U2652 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n755, D1 => 
                           registers_30_13_port, S1 => n6448, D2 => n6445, S2 
                           => n659, D3 => registers_20_13_port, S3 => n6442, Z 
                           => n1267);
   U2653 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n754, D1 => 
                           registers_30_14_port, S1 => n6448, D2 => n6445, S2 
                           => n658, D3 => registers_20_14_port, S3 => n6442, Z 
                           => n1253);
   U2654 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n753, D1 => 
                           registers_30_15_port, S1 => n6448, D2 => n6445, S2 
                           => n657, D3 => registers_20_15_port, S3 => n6442, Z 
                           => n1239);
   U2655 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n752, D1 => 
                           registers_30_16_port, S1 => n6448, D2 => n6445, S2 
                           => n656, D3 => registers_20_16_port, S3 => n6442, Z 
                           => n1225);
   U2656 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n751, D1 => 
                           registers_30_17_port, S1 => n6448, D2 => n6445, S2 
                           => n655, D3 => registers_20_17_port, S3 => n6442, Z 
                           => n1211);
   U2657 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n750, D1 => 
                           registers_30_18_port, S1 => n6448, D2 => n6445, S2 
                           => n654, D3 => registers_20_18_port, S3 => n6442, Z 
                           => n1197);
   U2658 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n749, D1 => 
                           registers_30_19_port, S1 => n6448, D2 => n6445, S2 
                           => n653, D3 => registers_20_19_port, S3 => n6442, Z 
                           => n1183);
   U2659 : HS65_LH_MX41X7 port map( D0 => n6451, S0 => n748, D1 => 
                           registers_30_20_port, S1 => n6449, D2 => n6445, S2 
                           => n652, D3 => registers_20_20_port, S3 => n6443, Z 
                           => n1155);
   U2660 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n747, D1 => 
                           registers_30_21_port, S1 => n6449, D2 => n6446, S2 
                           => n651, D3 => registers_20_21_port, S3 => n6443, Z 
                           => n1141);
   U2661 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n746, D1 => 
                           registers_30_22_port, S1 => n6449, D2 => n6446, S2 
                           => n650, D3 => registers_20_22_port, S3 => n6443, Z 
                           => n1127);
   U2662 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n745, D1 => 
                           registers_30_23_port, S1 => n6449, D2 => n6446, S2 
                           => n649, D3 => registers_20_23_port, S3 => n6443, Z 
                           => n1113);
   U2663 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n744, D1 => 
                           registers_30_24_port, S1 => n6449, D2 => n6446, S2 
                           => n648, D3 => registers_20_24_port, S3 => n6443, Z 
                           => n1099);
   U2664 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n743, D1 => 
                           registers_30_25_port, S1 => n6449, D2 => n6446, S2 
                           => n647, D3 => registers_20_25_port, S3 => n6443, Z 
                           => n1085);
   U2665 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n742, D1 => 
                           registers_30_26_port, S1 => n6449, D2 => n6446, S2 
                           => n646, D3 => registers_20_26_port, S3 => n6443, Z 
                           => n1071);
   U2666 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n741, D1 => 
                           registers_30_27_port, S1 => n6449, D2 => n6446, S2 
                           => n645, D3 => registers_20_27_port, S3 => n6443, Z 
                           => n1057);
   U2667 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n740, D1 => 
                           registers_30_28_port, S1 => n6449, D2 => n6446, S2 
                           => n644, D3 => registers_20_28_port, S3 => n6443, Z 
                           => n1043);
   U2668 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n739, D1 => 
                           registers_30_29_port, S1 => n6449, D2 => n6446, S2 
                           => n643, D3 => registers_20_29_port, S3 => n6443, Z 
                           => n1029);
   U2669 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n738, D1 => 
                           registers_30_30_port, S1 => n6449, D2 => n6446, S2 
                           => n642, D3 => registers_20_30_port, S3 => n6443, Z 
                           => n1001);
   U2670 : HS65_LH_MX41X7 port map( D0 => n6452, S0 => n737, D1 => 
                           registers_30_31_port, S1 => n6450, D2 => n6446, S2 
                           => n641, D3 => registers_20_31_port, S3 => n6444, Z 
                           => n987);
   U2671 : HS65_LH_MX41X7 port map( D0 => registers_2_0_port, S0 => n6499, D1 
                           => n6496, S1 => n640, D2 => n6493, S2 => n576, D3 =>
                           registers_23_0_port, S3 => n6490, Z => n1318);
   U2672 : HS65_LH_IVX9 port map( A => n160, Z => n576);
   U2673 : HS65_LH_MX41X7 port map( D0 => registers_2_1_port, S0 => n6499, D1 
                           => n6496, S1 => n639, D2 => n6493, S2 => n575, D3 =>
                           registers_23_1_port, S3 => n6490, Z => n1164);
   U2674 : HS65_LH_IVX9 port map( A => n159, Z => n575);
   U2675 : HS65_LH_MX41X7 port map( D0 => registers_2_2_port, S0 => n6500, D1 
                           => n6497, S1 => n638, D2 => n6494, S2 => n574, D3 =>
                           registers_23_2_port, S3 => n6491, Z => n1010);
   U2676 : HS65_LH_IVX9 port map( A => n158, Z => n574);
   U2677 : HS65_LH_MX41X7 port map( D0 => registers_2_3_port, S0 => n6501, D1 
                           => n6498, S1 => n637, D2 => n6494, S2 => n573, D3 =>
                           registers_23_3_port, S3 => n6492, Z => n968);
   U2678 : HS65_LH_IVX9 port map( A => n157, Z => n573);
   U2679 : HS65_LH_MX41X7 port map( D0 => registers_2_4_port, S0 => n6501, D1 
                           => n6498, S1 => n636, D2 => n6495, S2 => n572, D3 =>
                           registers_23_4_port, S3 => n6492, Z => n954);
   U2680 : HS65_LH_IVX9 port map( A => n156, Z => n572);
   U2681 : HS65_LH_MX41X7 port map( D0 => registers_2_5_port, S0 => n6501, D1 
                           => n6498, S1 => n635, D2 => n6495, S2 => n571, D3 =>
                           registers_23_5_port, S3 => n6492, Z => n940);
   U2682 : HS65_LH_IVX9 port map( A => n155, Z => n571);
   U2683 : HS65_LH_MX41X7 port map( D0 => registers_2_6_port, S0 => n6501, D1 
                           => n6498, S1 => n634, D2 => n6495, S2 => n570, D3 =>
                           registers_23_6_port, S3 => n6492, Z => n926);
   U2684 : HS65_LH_IVX9 port map( A => n154, Z => n570);
   U2685 : HS65_LH_MX41X7 port map( D0 => registers_2_7_port, S0 => n6501, D1 
                           => n6498, S1 => n633, D2 => n6495, S2 => n569, D3 =>
                           registers_23_7_port, S3 => n6492, Z => n912);
   U2686 : HS65_LH_IVX9 port map( A => n153, Z => n569);
   U2687 : HS65_LH_MX41X7 port map( D0 => registers_2_8_port, S0 => n6501, D1 
                           => n6498, S1 => n632, D2 => n6495, S2 => n568, D3 =>
                           registers_23_8_port, S3 => n6492, Z => n898);
   U2688 : HS65_LH_IVX9 port map( A => n152, Z => n568);
   U2689 : HS65_LH_MX41X7 port map( D0 => registers_2_9_port, S0 => n6501, D1 
                           => n6498, S1 => n631, D2 => n6495, S2 => n567, D3 =>
                           registers_23_9_port, S3 => n6492, Z => n853);
   U2690 : HS65_LH_IVX9 port map( A => n151, Z => n567);
   U2691 : HS65_LH_MX41X7 port map( D0 => registers_2_10_port, S0 => n6499, D1 
                           => n6496, S1 => n630, D2 => n6493, S2 => n566, D3 =>
                           registers_23_10_port, S3 => n6490, Z => n1304);
   U2692 : HS65_LH_IVX9 port map( A => n150, Z => n566);
   U2693 : HS65_LH_MX41X7 port map( D0 => registers_2_11_port, S0 => n6499, D1 
                           => n6496, S1 => n629, D2 => n6493, S2 => n565, D3 =>
                           registers_23_11_port, S3 => n6490, Z => n1290);
   U2694 : HS65_LH_IVX9 port map( A => n149, Z => n565);
   U2695 : HS65_LH_MX41X7 port map( D0 => registers_2_12_port, S0 => n6499, D1 
                           => n6496, S1 => n628, D2 => n6493, S2 => n564, D3 =>
                           registers_23_12_port, S3 => n6490, Z => n1276);
   U2696 : HS65_LH_IVX9 port map( A => n148, Z => n564);
   U2697 : HS65_LH_MX41X7 port map( D0 => registers_2_13_port, S0 => n6499, D1 
                           => n6496, S1 => n627, D2 => n6493, S2 => n563, D3 =>
                           registers_23_13_port, S3 => n6490, Z => n1262);
   U2698 : HS65_LH_IVX9 port map( A => n147, Z => n563);
   U2699 : HS65_LH_MX41X7 port map( D0 => registers_2_14_port, S0 => n6499, D1 
                           => n6496, S1 => n626, D2 => n6493, S2 => n562, D3 =>
                           registers_23_14_port, S3 => n6490, Z => n1248);
   U2700 : HS65_LH_IVX9 port map( A => n146, Z => n562);
   U2701 : HS65_LH_MX41X7 port map( D0 => registers_2_15_port, S0 => n6499, D1 
                           => n6496, S1 => n625, D2 => n6493, S2 => n561, D3 =>
                           registers_23_15_port, S3 => n6490, Z => n1234);
   U2702 : HS65_LH_IVX9 port map( A => n145, Z => n561);
   U2703 : HS65_LH_MX41X7 port map( D0 => registers_2_16_port, S0 => n6499, D1 
                           => n6496, S1 => n624, D2 => n6493, S2 => n560, D3 =>
                           registers_23_16_port, S3 => n6490, Z => n1220);
   U2704 : HS65_LH_IVX9 port map( A => n144, Z => n560);
   U2705 : HS65_LH_MX41X7 port map( D0 => registers_2_17_port, S0 => n6499, D1 
                           => n6496, S1 => n623, D2 => n6493, S2 => n559, D3 =>
                           registers_23_17_port, S3 => n6490, Z => n1206);
   U2706 : HS65_LH_IVX9 port map( A => n143, Z => n559);
   U2707 : HS65_LH_MX41X7 port map( D0 => registers_2_18_port, S0 => n6499, D1 
                           => n6496, S1 => n622, D2 => n6493, S2 => n558, D3 =>
                           registers_23_18_port, S3 => n6490, Z => n1192);
   U2708 : HS65_LH_IVX9 port map( A => n142, Z => n558);
   U2709 : HS65_LH_MX41X7 port map( D0 => registers_2_19_port, S0 => n6499, D1 
                           => n6496, S1 => n621, D2 => n6493, S2 => n557, D3 =>
                           registers_23_19_port, S3 => n6490, Z => n1178);
   U2710 : HS65_LH_IVX9 port map( A => n141, Z => n557);
   U2711 : HS65_LH_MX41X7 port map( D0 => registers_2_20_port, S0 => n6500, D1 
                           => n6497, S1 => n620, D2 => n6493, S2 => n556, D3 =>
                           registers_23_20_port, S3 => n6491, Z => n1150);
   U2712 : HS65_LH_IVX9 port map( A => n140, Z => n556);
   U2713 : HS65_LH_MX41X7 port map( D0 => registers_2_21_port, S0 => n6500, D1 
                           => n6497, S1 => n619, D2 => n6494, S2 => n555, D3 =>
                           registers_23_21_port, S3 => n6491, Z => n1136);
   U2714 : HS65_LH_IVX9 port map( A => n139, Z => n555);
   U2715 : HS65_LH_MX41X7 port map( D0 => registers_2_22_port, S0 => n6500, D1 
                           => n6497, S1 => n618, D2 => n6494, S2 => n554, D3 =>
                           registers_23_22_port, S3 => n6491, Z => n1122);
   U2716 : HS65_LH_IVX9 port map( A => n138, Z => n554);
   U2717 : HS65_LH_MX41X7 port map( D0 => registers_2_23_port, S0 => n6500, D1 
                           => n6497, S1 => n617, D2 => n6494, S2 => n553, D3 =>
                           registers_23_23_port, S3 => n6491, Z => n1108);
   U2718 : HS65_LH_IVX9 port map( A => n137, Z => n553);
   U2719 : HS65_LH_MX41X7 port map( D0 => registers_2_24_port, S0 => n6500, D1 
                           => n6497, S1 => n616, D2 => n6494, S2 => n552, D3 =>
                           registers_23_24_port, S3 => n6491, Z => n1094);
   U2720 : HS65_LH_IVX9 port map( A => n136, Z => n552);
   U2721 : HS65_LH_MX41X7 port map( D0 => registers_2_25_port, S0 => n6500, D1 
                           => n6497, S1 => n615, D2 => n6494, S2 => n551, D3 =>
                           registers_23_25_port, S3 => n6491, Z => n1080);
   U2722 : HS65_LH_IVX9 port map( A => n135, Z => n551);
   U2723 : HS65_LH_MX41X7 port map( D0 => registers_2_26_port, S0 => n6500, D1 
                           => n6497, S1 => n614, D2 => n6494, S2 => n550, D3 =>
                           registers_23_26_port, S3 => n6491, Z => n1066);
   U2724 : HS65_LH_IVX9 port map( A => n134, Z => n550);
   U2725 : HS65_LH_MX41X7 port map( D0 => registers_2_27_port, S0 => n6500, D1 
                           => n6497, S1 => n613, D2 => n6494, S2 => n549, D3 =>
                           registers_23_27_port, S3 => n6491, Z => n1052);
   U2726 : HS65_LH_IVX9 port map( A => n133, Z => n549);
   U2727 : HS65_LH_MX41X7 port map( D0 => registers_2_28_port, S0 => n6500, D1 
                           => n6497, S1 => n612, D2 => n6494, S2 => n548, D3 =>
                           registers_23_28_port, S3 => n6491, Z => n1038);
   U2728 : HS65_LH_IVX9 port map( A => n132, Z => n548);
   U2729 : HS65_LH_MX41X7 port map( D0 => registers_2_29_port, S0 => n6500, D1 
                           => n6497, S1 => n611, D2 => n6494, S2 => n547, D3 =>
                           registers_23_29_port, S3 => n6491, Z => n1024);
   U2730 : HS65_LH_IVX9 port map( A => n131, Z => n547);
   U2731 : HS65_LH_MX41X7 port map( D0 => registers_2_30_port, S0 => n6500, D1 
                           => n6497, S1 => n610, D2 => n6494, S2 => n546, D3 =>
                           registers_23_30_port, S3 => n6491, Z => n996);
   U2732 : HS65_LH_IVX9 port map( A => n130, Z => n546);
   U2733 : HS65_LH_MX41X7 port map( D0 => registers_2_31_port, S0 => n6501, D1 
                           => n6498, S1 => n609, D2 => n6494, S2 => n545, D3 =>
                           registers_23_31_port, S3 => n6492, Z => n982);
   U2734 : HS65_LH_IVX9 port map( A => n129, Z => n545);
   U2735 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_0_port, D1 
                           => n6391, S1 => registers_4_0_port, D2 => n6388, S2 
                           => registers_5_0_port, D3 => n6385, S3 => 
                           registers_1_0_port, Z => n2800);
   U2736 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_1_port, D1 
                           => n6391, S1 => registers_4_1_port, D2 => n6388, S2 
                           => registers_5_1_port, D3 => n6385, S3 => 
                           registers_1_1_port, Z => n2646);
   U2737 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_2_port, D1 
                           => n6392, S1 => registers_4_2_port, D2 => n6389, S2 
                           => registers_5_2_port, D3 => n6386, S3 => 
                           registers_1_2_port, Z => n2492);
   U2738 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_3_port, D1 
                           => n6393, S1 => registers_4_3_port, D2 => n6389, S2 
                           => registers_5_3_port, D3 => n6387, S3 => 
                           registers_1_3_port, Z => n2450);
   U2739 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_4_port, D1 
                           => n6393, S1 => registers_4_4_port, D2 => n6390, S2 
                           => registers_5_4_port, D3 => n6387, S3 => 
                           registers_1_4_port, Z => n2436);
   U2740 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_5_port, D1 
                           => n6393, S1 => registers_4_5_port, D2 => n6390, S2 
                           => registers_5_5_port, D3 => n6387, S3 => 
                           registers_1_5_port, Z => n1430);
   U2741 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_6_port, D1 
                           => n6393, S1 => registers_4_6_port, D2 => n6390, S2 
                           => registers_5_6_port, D3 => n6387, S3 => 
                           registers_1_6_port, Z => n1416);
   U2742 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_7_port, D1 
                           => n6393, S1 => registers_4_7_port, D2 => n6390, S2 
                           => registers_5_7_port, D3 => n6387, S3 => 
                           registers_1_7_port, Z => n1402);
   U2743 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_8_port, D1 
                           => n6393, S1 => registers_4_8_port, D2 => n6390, S2 
                           => registers_5_8_port, D3 => n6387, S3 => 
                           registers_1_8_port, Z => n1388);
   U2744 : HS65_LH_MX41X7 port map( D0 => n6396, S0 => registers_7_9_port, D1 
                           => n6393, S1 => registers_4_9_port, D2 => n6390, S2 
                           => registers_5_9_port, D3 => n6387, S3 => 
                           registers_1_9_port, Z => n1343);
   U2745 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_10_port, D1 
                           => n6391, S1 => registers_4_10_port, D2 => n6388, S2
                           => registers_5_10_port, D3 => n6385, S3 => 
                           registers_1_10_port, Z => n2786);
   U2746 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_11_port, D1 
                           => n6391, S1 => registers_4_11_port, D2 => n6388, S2
                           => registers_5_11_port, D3 => n6385, S3 => 
                           registers_1_11_port, Z => n2772);
   U2747 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_12_port, D1 
                           => n6391, S1 => registers_4_12_port, D2 => n6388, S2
                           => registers_5_12_port, D3 => n6385, S3 => 
                           registers_1_12_port, Z => n2758);
   U2748 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_13_port, D1 
                           => n6391, S1 => registers_4_13_port, D2 => n6388, S2
                           => registers_5_13_port, D3 => n6385, S3 => 
                           registers_1_13_port, Z => n2744);
   U2749 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_14_port, D1 
                           => n6391, S1 => registers_4_14_port, D2 => n6388, S2
                           => registers_5_14_port, D3 => n6385, S3 => 
                           registers_1_14_port, Z => n2730);
   U2750 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_15_port, D1 
                           => n6391, S1 => registers_4_15_port, D2 => n6388, S2
                           => registers_5_15_port, D3 => n6385, S3 => 
                           registers_1_15_port, Z => n2716);
   U2751 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_16_port, D1 
                           => n6391, S1 => registers_4_16_port, D2 => n6388, S2
                           => registers_5_16_port, D3 => n6385, S3 => 
                           registers_1_16_port, Z => n2702);
   U2752 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_17_port, D1 
                           => n6391, S1 => registers_4_17_port, D2 => n6388, S2
                           => registers_5_17_port, D3 => n6385, S3 => 
                           registers_1_17_port, Z => n2688);
   U2753 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_18_port, D1 
                           => n6391, S1 => registers_4_18_port, D2 => n6388, S2
                           => registers_5_18_port, D3 => n6385, S3 => 
                           registers_1_18_port, Z => n2674);
   U2754 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_19_port, D1 
                           => n6391, S1 => registers_4_19_port, D2 => n6388, S2
                           => registers_5_19_port, D3 => n6385, S3 => 
                           registers_1_19_port, Z => n2660);
   U2755 : HS65_LH_MX41X7 port map( D0 => n6394, S0 => registers_7_20_port, D1 
                           => n6392, S1 => registers_4_20_port, D2 => n6388, S2
                           => registers_5_20_port, D3 => n6386, S3 => 
                           registers_1_20_port, Z => n2632);
   U2756 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_21_port, D1 
                           => n6392, S1 => registers_4_21_port, D2 => n6389, S2
                           => registers_5_21_port, D3 => n6386, S3 => 
                           registers_1_21_port, Z => n2618);
   U2757 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_22_port, D1 
                           => n6392, S1 => registers_4_22_port, D2 => n6389, S2
                           => registers_5_22_port, D3 => n6386, S3 => 
                           registers_1_22_port, Z => n2604);
   U2758 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_23_port, D1 
                           => n6392, S1 => registers_4_23_port, D2 => n6389, S2
                           => registers_5_23_port, D3 => n6386, S3 => 
                           registers_1_23_port, Z => n2590);
   U2759 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_24_port, D1 
                           => n6392, S1 => registers_4_24_port, D2 => n6389, S2
                           => registers_5_24_port, D3 => n6386, S3 => 
                           registers_1_24_port, Z => n2576);
   U2760 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_25_port, D1 
                           => n6392, S1 => registers_4_25_port, D2 => n6389, S2
                           => registers_5_25_port, D3 => n6386, S3 => 
                           registers_1_25_port, Z => n2562);
   U2761 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_26_port, D1 
                           => n6392, S1 => registers_4_26_port, D2 => n6389, S2
                           => registers_5_26_port, D3 => n6386, S3 => 
                           registers_1_26_port, Z => n2548);
   U2762 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_27_port, D1 
                           => n6392, S1 => registers_4_27_port, D2 => n6389, S2
                           => registers_5_27_port, D3 => n6386, S3 => 
                           registers_1_27_port, Z => n2534);
   U2763 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_28_port, D1 
                           => n6392, S1 => registers_4_28_port, D2 => n6389, S2
                           => registers_5_28_port, D3 => n6386, S3 => 
                           registers_1_28_port, Z => n2520);
   U2764 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_29_port, D1 
                           => n6392, S1 => registers_4_29_port, D2 => n6389, S2
                           => registers_5_29_port, D3 => n6386, S3 => 
                           registers_1_29_port, Z => n2506);
   U2765 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_30_port, D1 
                           => n6392, S1 => registers_4_30_port, D2 => n6389, S2
                           => registers_5_30_port, D3 => n6386, S3 => 
                           registers_1_30_port, Z => n2478);
   U2766 : HS65_LH_MX41X7 port map( D0 => n6395, S0 => registers_7_31_port, D1 
                           => n6393, S1 => registers_4_31_port, D2 => n6389, S2
                           => registers_5_31_port, D3 => n6387, S3 => 
                           registers_1_31_port, Z => n2464);
   U2767 : HS65_LH_MX41X7 port map( D0 => registers_22_0_port, S0 => n6439, D1 
                           => registers_21_0_port, S1 => n6436, D2 => 
                           registers_19_0_port, S2 => n6433, D3 => n6430, S3 =>
                           n608, Z => n1332);
   U2768 : HS65_LH_MX41X7 port map( D0 => registers_22_1_port, S0 => n6439, D1 
                           => registers_21_1_port, S1 => n6436, D2 => 
                           registers_19_1_port, S2 => n6433, D3 => n6430, S3 =>
                           n607, Z => n1168);
   U2769 : HS65_LH_MX41X7 port map( D0 => registers_22_2_port, S0 => n6440, D1 
                           => registers_21_2_port, S1 => n6437, D2 => 
                           registers_19_2_port, S2 => n6434, D3 => n6431, S3 =>
                           n606, Z => n1014);
   U2770 : HS65_LH_MX41X7 port map( D0 => registers_22_3_port, S0 => n6441, D1 
                           => registers_21_3_port, S1 => n6438, D2 => 
                           registers_19_3_port, S2 => n6435, D3 => n6432, S3 =>
                           n605, Z => n972);
   U2771 : HS65_LH_MX41X7 port map( D0 => registers_22_4_port, S0 => n6441, D1 
                           => registers_21_4_port, S1 => n6438, D2 => 
                           registers_19_4_port, S2 => n6435, D3 => n6432, S3 =>
                           n604, Z => n958);
   U2772 : HS65_LH_MX41X7 port map( D0 => registers_22_5_port, S0 => n6441, D1 
                           => registers_21_5_port, S1 => n6438, D2 => 
                           registers_19_5_port, S2 => n6435, D3 => n6432, S3 =>
                           n603, Z => n944);
   U2773 : HS65_LH_MX41X7 port map( D0 => registers_22_6_port, S0 => n6441, D1 
                           => registers_21_6_port, S1 => n6438, D2 => 
                           registers_19_6_port, S2 => n6435, D3 => n6432, S3 =>
                           n602, Z => n930);
   U2774 : HS65_LH_MX41X7 port map( D0 => registers_22_7_port, S0 => n6441, D1 
                           => registers_21_7_port, S1 => n6438, D2 => 
                           registers_19_7_port, S2 => n6435, D3 => n6432, S3 =>
                           n601, Z => n916);
   U2775 : HS65_LH_MX41X7 port map( D0 => registers_22_8_port, S0 => n6441, D1 
                           => registers_21_8_port, S1 => n6438, D2 => 
                           registers_19_8_port, S2 => n6435, D3 => n6432, S3 =>
                           n600, Z => n902);
   U2776 : HS65_LH_MX41X7 port map( D0 => registers_22_9_port, S0 => n6441, D1 
                           => registers_21_9_port, S1 => n6438, D2 => 
                           registers_19_9_port, S2 => n6435, D3 => n6432, S3 =>
                           n599, Z => n872);
   U2777 : HS65_LH_MX41X7 port map( D0 => registers_22_11_port, S0 => n6439, D1
                           => registers_21_11_port, S1 => n6436, D2 => 
                           registers_19_11_port, S2 => n6433, D3 => n6430, S3 
                           => n597, Z => n1294);
   U2778 : HS65_LH_MX41X7 port map( D0 => registers_22_12_port, S0 => n6439, D1
                           => registers_21_12_port, S1 => n6436, D2 => 
                           registers_19_12_port, S2 => n6433, D3 => n6430, S3 
                           => n596, Z => n1280);
   U2779 : HS65_LH_MX41X7 port map( D0 => registers_22_13_port, S0 => n6439, D1
                           => registers_21_13_port, S1 => n6436, D2 => 
                           registers_19_13_port, S2 => n6433, D3 => n6430, S3 
                           => n595, Z => n1266);
   U2780 : HS65_LH_MX41X7 port map( D0 => registers_22_14_port, S0 => n6439, D1
                           => registers_21_14_port, S1 => n6436, D2 => 
                           registers_19_14_port, S2 => n6433, D3 => n6430, S3 
                           => n594, Z => n1252);
   U2781 : HS65_LH_MX41X7 port map( D0 => registers_22_15_port, S0 => n6439, D1
                           => registers_21_15_port, S1 => n6436, D2 => 
                           registers_19_15_port, S2 => n6433, D3 => n6430, S3 
                           => n593, Z => n1238);
   U2782 : HS65_LH_MX41X7 port map( D0 => registers_22_16_port, S0 => n6439, D1
                           => registers_21_16_port, S1 => n6436, D2 => 
                           registers_19_16_port, S2 => n6433, D3 => n6430, S3 
                           => n592, Z => n1224);
   U2783 : HS65_LH_MX41X7 port map( D0 => registers_22_17_port, S0 => n6439, D1
                           => registers_21_17_port, S1 => n6436, D2 => 
                           registers_19_17_port, S2 => n6433, D3 => n6430, S3 
                           => n591, Z => n1210);
   U2784 : HS65_LH_MX41X7 port map( D0 => registers_22_18_port, S0 => n6439, D1
                           => registers_21_18_port, S1 => n6436, D2 => 
                           registers_19_18_port, S2 => n6433, D3 => n6430, S3 
                           => n590, Z => n1196);
   U2785 : HS65_LH_MX41X7 port map( D0 => registers_22_19_port, S0 => n6439, D1
                           => registers_21_19_port, S1 => n6436, D2 => 
                           registers_19_19_port, S2 => n6433, D3 => n6430, S3 
                           => n589, Z => n1182);
   U2786 : HS65_LH_MX41X7 port map( D0 => registers_22_20_port, S0 => n6440, D1
                           => registers_21_20_port, S1 => n6437, D2 => 
                           registers_19_20_port, S2 => n6434, D3 => n6431, S3 
                           => n588, Z => n1154);
   U2787 : HS65_LH_MX41X7 port map( D0 => registers_22_21_port, S0 => n6440, D1
                           => registers_21_21_port, S1 => n6437, D2 => 
                           registers_19_21_port, S2 => n6434, D3 => n6431, S3 
                           => n587, Z => n1140);
   U2788 : HS65_LH_MX41X7 port map( D0 => registers_22_22_port, S0 => n6440, D1
                           => registers_21_22_port, S1 => n6437, D2 => 
                           registers_19_22_port, S2 => n6434, D3 => n6431, S3 
                           => n586, Z => n1126);
   U2789 : HS65_LH_MX41X7 port map( D0 => registers_22_23_port, S0 => n6440, D1
                           => registers_21_23_port, S1 => n6437, D2 => 
                           registers_19_23_port, S2 => n6434, D3 => n6431, S3 
                           => n585, Z => n1112);
   U2790 : HS65_LH_MX41X7 port map( D0 => registers_22_24_port, S0 => n6440, D1
                           => registers_21_24_port, S1 => n6437, D2 => 
                           registers_19_24_port, S2 => n6434, D3 => n6431, S3 
                           => n584, Z => n1098);
   U2791 : HS65_LH_MX41X7 port map( D0 => registers_22_25_port, S0 => n6440, D1
                           => registers_21_25_port, S1 => n6437, D2 => 
                           registers_19_25_port, S2 => n6434, D3 => n6431, S3 
                           => n583, Z => n1084);
   U2792 : HS65_LH_MX41X7 port map( D0 => registers_22_26_port, S0 => n6440, D1
                           => registers_21_26_port, S1 => n6437, D2 => 
                           registers_19_26_port, S2 => n6434, D3 => n6431, S3 
                           => n582, Z => n1070);
   U2793 : HS65_LH_MX41X7 port map( D0 => registers_22_27_port, S0 => n6440, D1
                           => registers_21_27_port, S1 => n6437, D2 => 
                           registers_19_27_port, S2 => n6434, D3 => n6431, S3 
                           => n581, Z => n1056);
   U2794 : HS65_LH_MX41X7 port map( D0 => registers_22_28_port, S0 => n6440, D1
                           => registers_21_28_port, S1 => n6437, D2 => 
                           registers_19_28_port, S2 => n6434, D3 => n6431, S3 
                           => n580, Z => n1042);
   U2795 : HS65_LH_MX41X7 port map( D0 => registers_22_29_port, S0 => n6440, D1
                           => registers_21_29_port, S1 => n6437, D2 => 
                           registers_19_29_port, S2 => n6434, D3 => n6431, S3 
                           => n579, Z => n1028);
   U2796 : HS65_LH_MX41X7 port map( D0 => registers_22_30_port, S0 => n6440, D1
                           => registers_21_30_port, S1 => n6437, D2 => 
                           registers_19_30_port, S2 => n6434, D3 => n6431, S3 
                           => n578, Z => n1000);
   U2797 : HS65_LH_MX41X7 port map( D0 => registers_22_31_port, S0 => n6441, D1
                           => registers_21_31_port, S1 => n6438, D2 => 
                           registers_19_31_port, S2 => n6435, D3 => n6432, S3 
                           => n577, Z => n986);
   U2798 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n704, D1 => n6355, S1 =>
                           registers_30_0_port, D2 => n6352, S2 => n608, D3 => 
                           n6349, S3 => registers_20_0_port, Z => n2815);
   U2799 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n703, D1 => n6355, S1 =>
                           registers_30_1_port, D2 => n6352, S2 => n607, D3 => 
                           n6349, S3 => registers_20_1_port, Z => n2652);
   U2800 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n702, D1 => n6356, S1 =>
                           registers_30_2_port, D2 => n6353, S2 => n606, D3 => 
                           n6350, S3 => registers_20_2_port, Z => n2498);
   U2801 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n701, D1 => n6357, S1 =>
                           registers_30_3_port, D2 => n6353, S2 => n605, D3 => 
                           n6351, S3 => registers_20_3_port, Z => n2456);
   U2802 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n700, D1 => n6357, S1 =>
                           registers_30_4_port, D2 => n6354, S2 => n604, D3 => 
                           n6351, S3 => registers_20_4_port, Z => n2442);
   U2803 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n699, D1 => n6357, S1 =>
                           registers_30_5_port, D2 => n6354, S2 => n603, D3 => 
                           n6351, S3 => registers_20_5_port, Z => n2428);
   U2804 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n698, D1 => n6357, S1 =>
                           registers_30_6_port, D2 => n6354, S2 => n602, D3 => 
                           n6351, S3 => registers_20_6_port, Z => n1422);
   U2805 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n697, D1 => n6357, S1 =>
                           registers_30_7_port, D2 => n6354, S2 => n601, D3 => 
                           n6351, S3 => registers_20_7_port, Z => n1408);
   U2806 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n696, D1 => n6357, S1 =>
                           registers_30_8_port, D2 => n6354, S2 => n600, D3 => 
                           n6351, S3 => registers_20_8_port, Z => n1394);
   U2807 : HS65_LH_MX41X7 port map( D0 => n6360, S0 => n695, D1 => n6357, S1 =>
                           registers_30_9_port, D2 => n6354, S2 => n599, D3 => 
                           n6351, S3 => registers_20_9_port, Z => n1364);
   U2808 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n694, D1 => n6355, S1 =>
                           registers_30_10_port, D2 => n6352, S2 => n598, D3 =>
                           n6349, S3 => registers_20_10_port, Z => n2792);
   U2809 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n693, D1 => n6355, S1 =>
                           registers_30_11_port, D2 => n6352, S2 => n597, D3 =>
                           n6349, S3 => registers_20_11_port, Z => n2778);
   U2810 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n692, D1 => n6355, S1 =>
                           registers_30_12_port, D2 => n6352, S2 => n596, D3 =>
                           n6349, S3 => registers_20_12_port, Z => n2764);
   U2811 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n691, D1 => n6355, S1 =>
                           registers_30_13_port, D2 => n6352, S2 => n595, D3 =>
                           n6349, S3 => registers_20_13_port, Z => n2750);
   U2812 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n690, D1 => n6355, S1 =>
                           registers_30_14_port, D2 => n6352, S2 => n594, D3 =>
                           n6349, S3 => registers_20_14_port, Z => n2736);
   U2813 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n689, D1 => n6355, S1 =>
                           registers_30_15_port, D2 => n6352, S2 => n593, D3 =>
                           n6349, S3 => registers_20_15_port, Z => n2722);
   U2814 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n688, D1 => n6355, S1 =>
                           registers_30_16_port, D2 => n6352, S2 => n592, D3 =>
                           n6349, S3 => registers_20_16_port, Z => n2708);
   U2815 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n687, D1 => n6355, S1 =>
                           registers_30_17_port, D2 => n6352, S2 => n591, D3 =>
                           n6349, S3 => registers_20_17_port, Z => n2694);
   U2816 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n686, D1 => n6355, S1 =>
                           registers_30_18_port, D2 => n6352, S2 => n590, D3 =>
                           n6349, S3 => registers_20_18_port, Z => n2680);
   U2817 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n685, D1 => n6355, S1 =>
                           registers_30_19_port, D2 => n6352, S2 => n589, D3 =>
                           n6349, S3 => registers_20_19_port, Z => n2666);
   U2818 : HS65_LH_MX41X7 port map( D0 => n6358, S0 => n684, D1 => n6356, S1 =>
                           registers_30_20_port, D2 => n6352, S2 => n588, D3 =>
                           n6350, S3 => registers_20_20_port, Z => n2638);
   U2819 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n683, D1 => n6356, S1 =>
                           registers_30_21_port, D2 => n6353, S2 => n587, D3 =>
                           n6350, S3 => registers_20_21_port, Z => n2624);
   U2820 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n682, D1 => n6356, S1 =>
                           registers_30_22_port, D2 => n6353, S2 => n586, D3 =>
                           n6350, S3 => registers_20_22_port, Z => n2610);
   U2821 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n681, D1 => n6356, S1 =>
                           registers_30_23_port, D2 => n6353, S2 => n585, D3 =>
                           n6350, S3 => registers_20_23_port, Z => n2596);
   U2822 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n680, D1 => n6356, S1 =>
                           registers_30_24_port, D2 => n6353, S2 => n584, D3 =>
                           n6350, S3 => registers_20_24_port, Z => n2582);
   U2823 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n679, D1 => n6356, S1 =>
                           registers_30_25_port, D2 => n6353, S2 => n583, D3 =>
                           n6350, S3 => registers_20_25_port, Z => n2568);
   U2824 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n678, D1 => n6356, S1 =>
                           registers_30_26_port, D2 => n6353, S2 => n582, D3 =>
                           n6350, S3 => registers_20_26_port, Z => n2554);
   U2825 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n677, D1 => n6356, S1 =>
                           registers_30_27_port, D2 => n6353, S2 => n581, D3 =>
                           n6350, S3 => registers_20_27_port, Z => n2540);
   U2826 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n676, D1 => n6356, S1 =>
                           registers_30_28_port, D2 => n6353, S2 => n580, D3 =>
                           n6350, S3 => registers_20_28_port, Z => n2526);
   U2827 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n675, D1 => n6356, S1 =>
                           registers_30_29_port, D2 => n6353, S2 => n579, D3 =>
                           n6350, S3 => registers_20_29_port, Z => n2512);
   U2828 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n674, D1 => n6356, S1 =>
                           registers_30_30_port, D2 => n6353, S2 => n578, D3 =>
                           n6350, S3 => registers_20_30_port, Z => n2484);
   U2829 : HS65_LH_MX41X7 port map( D0 => n6359, S0 => n673, D1 => n6357, S1 =>
                           registers_30_31_port, D2 => n6353, S2 => n577, D3 =>
                           n6351, S3 => registers_20_31_port, Z => n2470);
   U2830 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_0_port, D1 
                           => n6343, S1 => registers_21_0_port, D2 => n6340, S2
                           => registers_23_0_port, D3 => n6337, S3 => 
                           registers_12_0_port, Z => n2814);
   U2831 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_1_port, D1 
                           => n6343, S1 => registers_21_1_port, D2 => n6340, S2
                           => registers_23_1_port, D3 => n6337, S3 => 
                           registers_12_1_port, Z => n2651);
   U2832 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_2_port, D1 
                           => n6344, S1 => registers_21_2_port, D2 => n6341, S2
                           => registers_23_2_port, D3 => n6338, S3 => 
                           registers_12_2_port, Z => n2497);
   U2833 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_3_port, D1 
                           => n6345, S1 => registers_21_3_port, D2 => n6341, S2
                           => registers_23_3_port, D3 => n6339, S3 => 
                           registers_12_3_port, Z => n2455);
   U2834 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_4_port, D1 
                           => n6345, S1 => registers_21_4_port, D2 => n6342, S2
                           => registers_23_4_port, D3 => n6339, S3 => 
                           registers_12_4_port, Z => n2441);
   U2835 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_5_port, D1 
                           => n6345, S1 => registers_21_5_port, D2 => n6342, S2
                           => registers_23_5_port, D3 => n6339, S3 => 
                           registers_12_5_port, Z => n2427);
   U2836 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_6_port, D1 
                           => n6345, S1 => registers_21_6_port, D2 => n6342, S2
                           => registers_23_6_port, D3 => n6339, S3 => 
                           registers_12_6_port, Z => n1421);
   U2837 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_7_port, D1 
                           => n6345, S1 => registers_21_7_port, D2 => n6342, S2
                           => registers_23_7_port, D3 => n6339, S3 => 
                           registers_12_7_port, Z => n1407);
   U2838 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_8_port, D1 
                           => n6345, S1 => registers_21_8_port, D2 => n6342, S2
                           => registers_23_8_port, D3 => n6339, S3 => 
                           registers_12_8_port, Z => n1393);
   U2839 : HS65_LH_MX41X7 port map( D0 => n6348, S0 => registers_22_9_port, D1 
                           => n6345, S1 => registers_21_9_port, D2 => n6342, S2
                           => registers_23_9_port, D3 => n6339, S3 => 
                           registers_12_9_port, Z => n1363);
   U2840 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_10_port, D1
                           => n6343, S1 => registers_21_10_port, D2 => n6340, 
                           S2 => registers_23_10_port, D3 => n6337, S3 => 
                           registers_12_10_port, Z => n2791);
   U2841 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_11_port, D1
                           => n6343, S1 => registers_21_11_port, D2 => n6340, 
                           S2 => registers_23_11_port, D3 => n6337, S3 => 
                           registers_12_11_port, Z => n2777);
   U2842 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_12_port, D1
                           => n6343, S1 => registers_21_12_port, D2 => n6340, 
                           S2 => registers_23_12_port, D3 => n6337, S3 => 
                           registers_12_12_port, Z => n2763);
   U2843 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_13_port, D1
                           => n6343, S1 => registers_21_13_port, D2 => n6340, 
                           S2 => registers_23_13_port, D3 => n6337, S3 => 
                           registers_12_13_port, Z => n2749);
   U2844 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_14_port, D1
                           => n6343, S1 => registers_21_14_port, D2 => n6340, 
                           S2 => registers_23_14_port, D3 => n6337, S3 => 
                           registers_12_14_port, Z => n2735);
   U2845 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_15_port, D1
                           => n6343, S1 => registers_21_15_port, D2 => n6340, 
                           S2 => registers_23_15_port, D3 => n6337, S3 => 
                           registers_12_15_port, Z => n2721);
   U2846 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_16_port, D1
                           => n6343, S1 => registers_21_16_port, D2 => n6340, 
                           S2 => registers_23_16_port, D3 => n6337, S3 => 
                           registers_12_16_port, Z => n2707);
   U2847 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_17_port, D1
                           => n6343, S1 => registers_21_17_port, D2 => n6340, 
                           S2 => registers_23_17_port, D3 => n6337, S3 => 
                           registers_12_17_port, Z => n2693);
   U2848 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_18_port, D1
                           => n6343, S1 => registers_21_18_port, D2 => n6340, 
                           S2 => registers_23_18_port, D3 => n6337, S3 => 
                           registers_12_18_port, Z => n2679);
   U2849 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_19_port, D1
                           => n6343, S1 => registers_21_19_port, D2 => n6340, 
                           S2 => registers_23_19_port, D3 => n6337, S3 => 
                           registers_12_19_port, Z => n2665);
   U2850 : HS65_LH_MX41X7 port map( D0 => n6346, S0 => registers_22_20_port, D1
                           => n6344, S1 => registers_21_20_port, D2 => n6340, 
                           S2 => registers_23_20_port, D3 => n6338, S3 => 
                           registers_12_20_port, Z => n2637);
   U2851 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_21_port, D1
                           => n6344, S1 => registers_21_21_port, D2 => n6341, 
                           S2 => registers_23_21_port, D3 => n6338, S3 => 
                           registers_12_21_port, Z => n2623);
   U2852 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_22_port, D1
                           => n6344, S1 => registers_21_22_port, D2 => n6341, 
                           S2 => registers_23_22_port, D3 => n6338, S3 => 
                           registers_12_22_port, Z => n2609);
   U2853 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_23_port, D1
                           => n6344, S1 => registers_21_23_port, D2 => n6341, 
                           S2 => registers_23_23_port, D3 => n6338, S3 => 
                           registers_12_23_port, Z => n2595);
   U2854 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_24_port, D1
                           => n6344, S1 => registers_21_24_port, D2 => n6341, 
                           S2 => registers_23_24_port, D3 => n6338, S3 => 
                           registers_12_24_port, Z => n2581);
   U2855 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_25_port, D1
                           => n6344, S1 => registers_21_25_port, D2 => n6341, 
                           S2 => registers_23_25_port, D3 => n6338, S3 => 
                           registers_12_25_port, Z => n2567);
   U2856 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_26_port, D1
                           => n6344, S1 => registers_21_26_port, D2 => n6341, 
                           S2 => registers_23_26_port, D3 => n6338, S3 => 
                           registers_12_26_port, Z => n2553);
   U2857 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_27_port, D1
                           => n6344, S1 => registers_21_27_port, D2 => n6341, 
                           S2 => registers_23_27_port, D3 => n6338, S3 => 
                           registers_12_27_port, Z => n2539);
   U2858 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_28_port, D1
                           => n6344, S1 => registers_21_28_port, D2 => n6341, 
                           S2 => registers_23_28_port, D3 => n6338, S3 => 
                           registers_12_28_port, Z => n2525);
   U2859 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_29_port, D1
                           => n6344, S1 => registers_21_29_port, D2 => n6341, 
                           S2 => registers_23_29_port, D3 => n6338, S3 => 
                           registers_12_29_port, Z => n2511);
   U2860 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_30_port, D1
                           => n6344, S1 => registers_21_30_port, D2 => n6341, 
                           S2 => registers_23_30_port, D3 => n6338, S3 => 
                           registers_12_30_port, Z => n2483);
   U2861 : HS65_LH_MX41X7 port map( D0 => n6347, S0 => registers_22_31_port, D1
                           => n6345, S1 => registers_21_31_port, D2 => n6341, 
                           S2 => registers_23_31_port, D3 => n6339, S3 => 
                           registers_12_31_port, Z => n2469);
   U2862 : HS65_LH_IVX9 port map( A => regfile_i(40), Z => n778);
   U2863 : HS65_LH_IVX9 port map( A => regfile_i(45), Z => n773);
   U2864 : HS65_LH_IVX9 port map( A => regfile_i(37), Z => n812);
   U2865 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n640, D1 => n6403, S1 =>
                           registers_2_0_port, D2 => n6400, S2 => 
                           registers_3_0_port, D3 => n6397, S3 => n768, Z => 
                           n2801);
   U2866 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n639, D1 => n6403, S1 =>
                           registers_2_1_port, D2 => n6400, S2 => 
                           registers_3_1_port, D3 => n6397, S3 => n767, Z => 
                           n2647);
   U2867 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n638, D1 => n6404, S1 =>
                           registers_2_2_port, D2 => n6401, S2 => 
                           registers_3_2_port, D3 => n6398, S3 => n766, Z => 
                           n2493);
   U2868 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n630, D1 => n6403, S1 =>
                           registers_2_10_port, D2 => n6400, S2 => 
                           registers_3_10_port, D3 => n6397, S3 => n758, Z => 
                           n2787);
   U2869 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n629, D1 => n6403, S1 =>
                           registers_2_11_port, D2 => n6400, S2 => 
                           registers_3_11_port, D3 => n6397, S3 => n757, Z => 
                           n2773);
   U2870 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n628, D1 => n6403, S1 =>
                           registers_2_12_port, D2 => n6400, S2 => 
                           registers_3_12_port, D3 => n6397, S3 => n756, Z => 
                           n2759);
   U2871 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n627, D1 => n6403, S1 =>
                           registers_2_13_port, D2 => n6400, S2 => 
                           registers_3_13_port, D3 => n6397, S3 => n755, Z => 
                           n2745);
   U2872 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n626, D1 => n6403, S1 =>
                           registers_2_14_port, D2 => n6400, S2 => 
                           registers_3_14_port, D3 => n6397, S3 => n754, Z => 
                           n2731);
   U2873 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n625, D1 => n6403, S1 =>
                           registers_2_15_port, D2 => n6400, S2 => 
                           registers_3_15_port, D3 => n6397, S3 => n753, Z => 
                           n2717);
   U2874 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n624, D1 => n6403, S1 =>
                           registers_2_16_port, D2 => n6400, S2 => 
                           registers_3_16_port, D3 => n6397, S3 => n752, Z => 
                           n2703);
   U2875 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n623, D1 => n6403, S1 =>
                           registers_2_17_port, D2 => n6400, S2 => 
                           registers_3_17_port, D3 => n6397, S3 => n751, Z => 
                           n2689);
   U2876 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n622, D1 => n6403, S1 =>
                           registers_2_18_port, D2 => n6400, S2 => 
                           registers_3_18_port, D3 => n6397, S3 => n750, Z => 
                           n2675);
   U2877 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n621, D1 => n6403, S1 =>
                           registers_2_19_port, D2 => n6400, S2 => 
                           registers_3_19_port, D3 => n6397, S3 => n749, Z => 
                           n2661);
   U2878 : HS65_LH_MX41X7 port map( D0 => n6406, S0 => n620, D1 => n6404, S1 =>
                           registers_2_20_port, D2 => n6400, S2 => 
                           registers_3_20_port, D3 => n6398, S3 => n748, Z => 
                           n2633);
   U2879 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n619, D1 => n6404, S1 =>
                           registers_2_21_port, D2 => n6401, S2 => 
                           registers_3_21_port, D3 => n6398, S3 => n747, Z => 
                           n2619);
   U2880 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n618, D1 => n6404, S1 =>
                           registers_2_22_port, D2 => n6401, S2 => 
                           registers_3_22_port, D3 => n6398, S3 => n746, Z => 
                           n2605);
   U2881 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n617, D1 => n6404, S1 =>
                           registers_2_23_port, D2 => n6401, S2 => 
                           registers_3_23_port, D3 => n6398, S3 => n745, Z => 
                           n2591);
   U2882 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n616, D1 => n6404, S1 =>
                           registers_2_24_port, D2 => n6401, S2 => 
                           registers_3_24_port, D3 => n6398, S3 => n744, Z => 
                           n2577);
   U2883 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n615, D1 => n6404, S1 =>
                           registers_2_25_port, D2 => n6401, S2 => 
                           registers_3_25_port, D3 => n6398, S3 => n743, Z => 
                           n2563);
   U2884 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n614, D1 => n6404, S1 =>
                           registers_2_26_port, D2 => n6401, S2 => 
                           registers_3_26_port, D3 => n6398, S3 => n742, Z => 
                           n2549);
   U2885 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n613, D1 => n6404, S1 =>
                           registers_2_27_port, D2 => n6401, S2 => 
                           registers_3_27_port, D3 => n6398, S3 => n741, Z => 
                           n2535);
   U2886 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n612, D1 => n6404, S1 =>
                           registers_2_28_port, D2 => n6401, S2 => 
                           registers_3_28_port, D3 => n6398, S3 => n740, Z => 
                           n2521);
   U2887 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n611, D1 => n6404, S1 =>
                           registers_2_29_port, D2 => n6401, S2 => 
                           registers_3_29_port, D3 => n6398, S3 => n739, Z => 
                           n2507);
   U2888 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n610, D1 => n6404, S1 =>
                           registers_2_30_port, D2 => n6401, S2 => 
                           registers_3_30_port, D3 => n6398, S3 => n738, Z => 
                           n2479);
   U2889 : HS65_LH_IVX9 port map( A => regfile_i(3), Z => n846);
   U2890 : HS65_LH_IVX9 port map( A => regfile_i(4), Z => n845);
   U2891 : HS65_LH_IVX9 port map( A => regfile_i(5), Z => n844);
   U2892 : HS65_LH_IVX9 port map( A => regfile_i(6), Z => n843);
   U2893 : HS65_LH_IVX9 port map( A => regfile_i(7), Z => n842);
   U2894 : HS65_LH_IVX9 port map( A => regfile_i(8), Z => n841);
   U2895 : HS65_LH_IVX9 port map( A => regfile_i(9), Z => n840);
   U2896 : HS65_LH_IVX9 port map( A => regfile_i(10), Z => n839);
   U2897 : HS65_LH_IVX9 port map( A => regfile_i(11), Z => n838);
   U2898 : HS65_LH_IVX9 port map( A => regfile_i(12), Z => n837);
   U2899 : HS65_LH_IVX9 port map( A => regfile_i(13), Z => n836);
   U2900 : HS65_LH_IVX9 port map( A => regfile_i(14), Z => n835);
   U2901 : HS65_LH_IVX9 port map( A => regfile_i(15), Z => n834);
   U2902 : HS65_LH_IVX9 port map( A => regfile_i(16), Z => n833);
   U2903 : HS65_LH_IVX9 port map( A => regfile_i(17), Z => n832);
   U2904 : HS65_LH_IVX9 port map( A => regfile_i(18), Z => n831);
   U2905 : HS65_LH_IVX9 port map( A => regfile_i(19), Z => n830);
   U2906 : HS65_LH_IVX9 port map( A => regfile_i(20), Z => n829);
   U2907 : HS65_LH_IVX9 port map( A => regfile_i(21), Z => n828);
   U2908 : HS65_LH_IVX9 port map( A => regfile_i(22), Z => n827);
   U2909 : HS65_LH_IVX9 port map( A => regfile_i(23), Z => n826);
   U2910 : HS65_LH_IVX9 port map( A => regfile_i(24), Z => n825);
   U2911 : HS65_LH_IVX9 port map( A => regfile_i(25), Z => n824);
   U2912 : HS65_LH_IVX9 port map( A => regfile_i(26), Z => n823);
   U2913 : HS65_LH_IVX9 port map( A => regfile_i(27), Z => n822);
   U2914 : HS65_LH_IVX9 port map( A => regfile_i(28), Z => n821);
   U2915 : HS65_LH_IVX9 port map( A => regfile_i(29), Z => n820);
   U2916 : HS65_LH_IVX9 port map( A => regfile_i(30), Z => n819);
   U2917 : HS65_LH_IVX9 port map( A => regfile_i(31), Z => n818);
   U2918 : HS65_LH_IVX9 port map( A => regfile_i(32), Z => n817);
   U2919 : HS65_LH_IVX9 port map( A => regfile_i(33), Z => n816);
   U2920 : HS65_LH_IVX9 port map( A => regfile_i(34), Z => n815);
   U2921 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n637, D1 => n6405, S1 =>
                           registers_2_3_port, D2 => n6401, S2 => 
                           registers_3_3_port, D3 => n6399, S3 => n765, Z => 
                           n2451);
   U2922 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n636, D1 => n6405, S1 =>
                           registers_2_4_port, D2 => n6402, S2 => 
                           registers_3_4_port, D3 => n6399, S3 => n764, Z => 
                           n2437);
   U2923 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n635, D1 => n6405, S1 =>
                           registers_2_5_port, D2 => n6402, S2 => 
                           registers_3_5_port, D3 => n6399, S3 => n763, Z => 
                           n1431);
   U2924 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n634, D1 => n6405, S1 =>
                           registers_2_6_port, D2 => n6402, S2 => 
                           registers_3_6_port, D3 => n6399, S3 => n762, Z => 
                           n1417);
   U2925 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n633, D1 => n6405, S1 =>
                           registers_2_7_port, D2 => n6402, S2 => 
                           registers_3_7_port, D3 => n6399, S3 => n761, Z => 
                           n1403);
   U2926 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n632, D1 => n6405, S1 =>
                           registers_2_8_port, D2 => n6402, S2 => 
                           registers_3_8_port, D3 => n6399, S3 => n760, Z => 
                           n1389);
   U2927 : HS65_LH_MX41X7 port map( D0 => n6408, S0 => n631, D1 => n6405, S1 =>
                           registers_2_9_port, D2 => n6402, S2 => 
                           registers_3_9_port, D3 => n6399, S3 => n759, Z => 
                           n1344);
   U2928 : HS65_LH_MX41X7 port map( D0 => n6407, S0 => n609, D1 => n6405, S1 =>
                           registers_2_31_port, D2 => n6401, S2 => 
                           registers_3_31_port, D3 => n6399, S3 => n737, Z => 
                           n2465);
   U2929 : HS65_LH_BFX9 port map( A => rst_n, Z => n6536);
   U2930 : HS65_LH_IVX9 port map( A => n96, Z => n544);
   U2931 : HS65_LH_IVX9 port map( A => n95, Z => n543);
   U2932 : HS65_LH_IVX9 port map( A => n94, Z => n542);
   U2933 : HS65_LH_IVX9 port map( A => n93, Z => n541);
   U2934 : HS65_LH_IVX9 port map( A => n92, Z => n540);
   U2935 : HS65_LH_IVX9 port map( A => n91, Z => n539);
   U2936 : HS65_LH_IVX9 port map( A => n90, Z => n538);
   U2937 : HS65_LH_IVX9 port map( A => n89, Z => n537);
   U2938 : HS65_LH_IVX9 port map( A => n88, Z => n536);
   U2939 : HS65_LH_IVX9 port map( A => n87, Z => n535);
   U2940 : HS65_LH_IVX9 port map( A => n86, Z => n534);
   U2941 : HS65_LH_IVX9 port map( A => n85, Z => n533);
   U2942 : HS65_LH_IVX9 port map( A => n84, Z => n532);
   U2943 : HS65_LH_IVX9 port map( A => n83, Z => n531);
   U2944 : HS65_LH_IVX9 port map( A => n82, Z => n530);
   U2945 : HS65_LH_IVX9 port map( A => n81, Z => n529);
   U2946 : HS65_LH_IVX9 port map( A => n80, Z => n528);
   U2947 : HS65_LH_IVX9 port map( A => n79, Z => n527);
   U2948 : HS65_LH_IVX9 port map( A => n78, Z => n526);
   U2949 : HS65_LH_IVX9 port map( A => n77, Z => n525);
   U2950 : HS65_LH_IVX9 port map( A => n76, Z => n524);
   U2951 : HS65_LH_IVX9 port map( A => n75, Z => n523);
   U2952 : HS65_LH_IVX9 port map( A => n74, Z => n522);
   U2953 : HS65_LH_IVX9 port map( A => n73, Z => n521);
   U2954 : HS65_LH_IVX9 port map( A => n72, Z => n520);
   U2955 : HS65_LH_IVX9 port map( A => n71, Z => n519);
   U2956 : HS65_LH_IVX9 port map( A => n70, Z => n518);
   U2957 : HS65_LH_IVX9 port map( A => n69, Z => n517);
   U2958 : HS65_LH_IVX9 port map( A => n68, Z => n516);
   U2959 : HS65_LH_IVX9 port map( A => n67, Z => n515);
   U2960 : HS65_LH_IVX9 port map( A => n66, Z => n514);
   U2961 : HS65_LH_IVX9 port map( A => n65, Z => n513);
   U2962 : HS65_LH_IVX9 port map( A => n32, Z => n704);
   U2963 : HS65_LH_IVX9 port map( A => n31, Z => n703);
   U2964 : HS65_LH_IVX9 port map( A => n30, Z => n702);
   U2965 : HS65_LH_IVX9 port map( A => n29, Z => n701);
   U2966 : HS65_LH_IVX9 port map( A => n28, Z => n700);
   U2967 : HS65_LH_IVX9 port map( A => n27, Z => n699);
   U2968 : HS65_LH_IVX9 port map( A => n26, Z => n698);
   U2969 : HS65_LH_IVX9 port map( A => n25, Z => n697);
   U2970 : HS65_LH_IVX9 port map( A => n24, Z => n696);
   U2971 : HS65_LH_IVX9 port map( A => n23, Z => n695);
   U2972 : HS65_LH_IVX9 port map( A => n22, Z => n694);
   U2973 : HS65_LH_IVX9 port map( A => n21, Z => n693);
   U2974 : HS65_LH_IVX9 port map( A => n20, Z => n692);
   U2975 : HS65_LH_IVX9 port map( A => n19, Z => n691);
   U2976 : HS65_LH_IVX9 port map( A => n18, Z => n690);
   U2977 : HS65_LH_IVX9 port map( A => n17, Z => n689);
   U2978 : HS65_LH_IVX9 port map( A => n16, Z => n688);
   U2979 : HS65_LH_IVX9 port map( A => n15, Z => n687);
   U2980 : HS65_LH_IVX9 port map( A => n14, Z => n686);
   U2981 : HS65_LH_IVX9 port map( A => n13, Z => n685);
   U2982 : HS65_LH_IVX9 port map( A => n12, Z => n684);
   U2983 : HS65_LH_IVX9 port map( A => n11, Z => n683);
   U2984 : HS65_LH_IVX9 port map( A => n10, Z => n682);
   U2985 : HS65_LH_IVX9 port map( A => n9, Z => n681);
   U2986 : HS65_LH_IVX9 port map( A => n8, Z => n680);
   U2987 : HS65_LH_IVX9 port map( A => n7, Z => n679);
   U2988 : HS65_LH_IVX9 port map( A => n6, Z => n678);
   U2989 : HS65_LH_IVX9 port map( A => n5, Z => n677);
   U2990 : HS65_LH_IVX9 port map( A => n4, Z => n676);
   U2991 : HS65_LH_IVX9 port map( A => n3, Z => n675);
   U2992 : HS65_LH_IVX9 port map( A => n2, Z => n674);
   U2993 : HS65_LH_IVX9 port map( A => n1, Z => n673);
   U2994 : HS65_LH_IVX9 port map( A => regfile_i(42), Z => n776);
   U2995 : HS65_LH_IVX9 port map( A => regfile_i(47), Z => n771);
   U2996 : HS65_LH_IVX9 port map( A => n128, Z => n672);
   U2997 : HS65_LH_IVX9 port map( A => n127, Z => n671);
   U2998 : HS65_LH_IVX9 port map( A => n126, Z => n670);
   U2999 : HS65_LH_IVX9 port map( A => n125, Z => n669);
   U3000 : HS65_LH_IVX9 port map( A => n124, Z => n668);
   U3001 : HS65_LH_IVX9 port map( A => n123, Z => n667);
   U3002 : HS65_LH_IVX9 port map( A => n122, Z => n666);
   U3003 : HS65_LH_IVX9 port map( A => n121, Z => n665);
   U3004 : HS65_LH_IVX9 port map( A => n120, Z => n664);
   U3005 : HS65_LH_IVX9 port map( A => n119, Z => n663);
   U3006 : HS65_LH_IVX9 port map( A => n118, Z => n662);
   U3007 : HS65_LH_IVX9 port map( A => n117, Z => n661);
   U3008 : HS65_LH_IVX9 port map( A => n116, Z => n660);
   U3009 : HS65_LH_IVX9 port map( A => n115, Z => n659);
   U3010 : HS65_LH_IVX9 port map( A => n114, Z => n658);
   U3011 : HS65_LH_IVX9 port map( A => n113, Z => n657);
   U3012 : HS65_LH_IVX9 port map( A => n112, Z => n656);
   U3013 : HS65_LH_IVX9 port map( A => n111, Z => n655);
   U3014 : HS65_LH_IVX9 port map( A => n110, Z => n654);
   U3015 : HS65_LH_IVX9 port map( A => n109, Z => n653);
   U3016 : HS65_LH_IVX9 port map( A => n108, Z => n652);
   U3017 : HS65_LH_IVX9 port map( A => n107, Z => n651);
   U3018 : HS65_LH_IVX9 port map( A => n106, Z => n650);
   U3019 : HS65_LH_IVX9 port map( A => n105, Z => n649);
   U3020 : HS65_LH_IVX9 port map( A => n104, Z => n648);
   U3021 : HS65_LH_IVX9 port map( A => n103, Z => n647);
   U3022 : HS65_LH_IVX9 port map( A => n102, Z => n646);
   U3023 : HS65_LH_IVX9 port map( A => n101, Z => n645);
   U3024 : HS65_LH_IVX9 port map( A => n100, Z => n644);
   U3025 : HS65_LH_IVX9 port map( A => n99, Z => n643);
   U3026 : HS65_LH_IVX9 port map( A => n98, Z => n642);
   U3027 : HS65_LH_IVX9 port map( A => n97, Z => n641);
   U3028 : HS65_LH_IVX9 port map( A => regfile_i(41), Z => n777);
   U3029 : HS65_LH_IVX9 port map( A => regfile_i(46), Z => n772);
   U3030 : HS65_LH_IVX9 port map( A => n256, Z => n768);
   U3031 : HS65_LH_IVX9 port map( A => n255, Z => n767);
   U3032 : HS65_LH_IVX9 port map( A => n254, Z => n766);
   U3033 : HS65_LH_IVX9 port map( A => n253, Z => n765);
   U3034 : HS65_LH_IVX9 port map( A => n252, Z => n764);
   U3035 : HS65_LH_IVX9 port map( A => n251, Z => n763);
   U3036 : HS65_LH_IVX9 port map( A => n250, Z => n762);
   U3037 : HS65_LH_IVX9 port map( A => n249, Z => n761);
   U3038 : HS65_LH_IVX9 port map( A => n248, Z => n760);
   U3039 : HS65_LH_IVX9 port map( A => n247, Z => n759);
   U3040 : HS65_LH_IVX9 port map( A => n246, Z => n758);
   U3041 : HS65_LH_IVX9 port map( A => n245, Z => n757);
   U3042 : HS65_LH_IVX9 port map( A => n244, Z => n756);
   U3043 : HS65_LH_IVX9 port map( A => n243, Z => n755);
   U3044 : HS65_LH_IVX9 port map( A => n242, Z => n754);
   U3045 : HS65_LH_IVX9 port map( A => n241, Z => n753);
   U3046 : HS65_LH_IVX9 port map( A => n240, Z => n752);
   U3047 : HS65_LH_IVX9 port map( A => n239, Z => n751);
   U3048 : HS65_LH_IVX9 port map( A => n238, Z => n750);
   U3049 : HS65_LH_IVX9 port map( A => n237, Z => n749);
   U3050 : HS65_LH_IVX9 port map( A => n236, Z => n748);
   U3051 : HS65_LH_IVX9 port map( A => n235, Z => n747);
   U3052 : HS65_LH_IVX9 port map( A => n234, Z => n746);
   U3053 : HS65_LH_IVX9 port map( A => n233, Z => n745);
   U3054 : HS65_LH_IVX9 port map( A => n232, Z => n744);
   U3055 : HS65_LH_IVX9 port map( A => n231, Z => n743);
   U3056 : HS65_LH_IVX9 port map( A => n230, Z => n742);
   U3057 : HS65_LH_IVX9 port map( A => n229, Z => n741);
   U3058 : HS65_LH_IVX9 port map( A => n228, Z => n740);
   U3059 : HS65_LH_IVX9 port map( A => n227, Z => n739);
   U3060 : HS65_LH_IVX9 port map( A => n226, Z => n738);
   U3061 : HS65_LH_IVX9 port map( A => n225, Z => n737);
   U3062 : HS65_LH_IVX9 port map( A => n64, Z => n608);
   U3063 : HS65_LH_IVX9 port map( A => n63, Z => n607);
   U3064 : HS65_LH_IVX9 port map( A => n62, Z => n606);
   U3065 : HS65_LH_IVX9 port map( A => n61, Z => n605);
   U3066 : HS65_LH_IVX9 port map( A => n60, Z => n604);
   U3067 : HS65_LH_IVX9 port map( A => n59, Z => n603);
   U3068 : HS65_LH_IVX9 port map( A => n58, Z => n602);
   U3069 : HS65_LH_IVX9 port map( A => n57, Z => n601);
   U3070 : HS65_LH_IVX9 port map( A => n56, Z => n600);
   U3071 : HS65_LH_IVX9 port map( A => n55, Z => n599);
   U3072 : HS65_LH_IVX9 port map( A => n54, Z => n598);
   U3073 : HS65_LH_IVX9 port map( A => n53, Z => n597);
   U3074 : HS65_LH_IVX9 port map( A => n52, Z => n596);
   U3075 : HS65_LH_IVX9 port map( A => n51, Z => n595);
   U3076 : HS65_LH_IVX9 port map( A => n50, Z => n594);
   U3077 : HS65_LH_IVX9 port map( A => n49, Z => n593);
   U3078 : HS65_LH_IVX9 port map( A => n48, Z => n592);
   U3079 : HS65_LH_IVX9 port map( A => n47, Z => n591);
   U3080 : HS65_LH_IVX9 port map( A => n46, Z => n590);
   U3081 : HS65_LH_IVX9 port map( A => n45, Z => n589);
   U3082 : HS65_LH_IVX9 port map( A => n44, Z => n588);
   U3083 : HS65_LH_IVX9 port map( A => n43, Z => n587);
   U3084 : HS65_LH_IVX9 port map( A => n42, Z => n586);
   U3085 : HS65_LH_IVX9 port map( A => n41, Z => n585);
   U3086 : HS65_LH_IVX9 port map( A => n40, Z => n584);
   U3087 : HS65_LH_IVX9 port map( A => n39, Z => n583);
   U3088 : HS65_LH_IVX9 port map( A => n38, Z => n582);
   U3089 : HS65_LH_IVX9 port map( A => n37, Z => n581);
   U3090 : HS65_LH_IVX9 port map( A => n36, Z => n580);
   U3091 : HS65_LH_IVX9 port map( A => n35, Z => n579);
   U3092 : HS65_LH_IVX9 port map( A => n34, Z => n578);
   U3093 : HS65_LH_IVX9 port map( A => n33, Z => n577);
   U3094 : HS65_LH_IVX9 port map( A => n192, Z => n640);
   U3095 : HS65_LH_IVX9 port map( A => n191, Z => n639);
   U3096 : HS65_LH_IVX9 port map( A => n190, Z => n638);
   U3097 : HS65_LH_IVX9 port map( A => n189, Z => n637);
   U3098 : HS65_LH_IVX9 port map( A => n188, Z => n636);
   U3099 : HS65_LH_IVX9 port map( A => n187, Z => n635);
   U3100 : HS65_LH_IVX9 port map( A => n186, Z => n634);
   U3101 : HS65_LH_IVX9 port map( A => n185, Z => n633);
   U3102 : HS65_LH_IVX9 port map( A => n184, Z => n632);
   U3103 : HS65_LH_IVX9 port map( A => n183, Z => n631);
   U3104 : HS65_LH_IVX9 port map( A => n182, Z => n630);
   U3105 : HS65_LH_IVX9 port map( A => n181, Z => n629);
   U3106 : HS65_LH_IVX9 port map( A => n180, Z => n628);
   U3107 : HS65_LH_IVX9 port map( A => n179, Z => n627);
   U3108 : HS65_LH_IVX9 port map( A => n178, Z => n626);
   U3109 : HS65_LH_IVX9 port map( A => n177, Z => n625);
   U3110 : HS65_LH_IVX9 port map( A => n176, Z => n624);
   U3111 : HS65_LH_IVX9 port map( A => n175, Z => n623);
   U3112 : HS65_LH_IVX9 port map( A => n174, Z => n622);
   U3113 : HS65_LH_IVX9 port map( A => n173, Z => n621);
   U3114 : HS65_LH_IVX9 port map( A => n172, Z => n620);
   U3115 : HS65_LH_IVX9 port map( A => n171, Z => n619);
   U3116 : HS65_LH_IVX9 port map( A => n170, Z => n618);
   U3117 : HS65_LH_IVX9 port map( A => n169, Z => n617);
   U3118 : HS65_LH_IVX9 port map( A => n168, Z => n616);
   U3119 : HS65_LH_IVX9 port map( A => n167, Z => n615);
   U3120 : HS65_LH_IVX9 port map( A => n166, Z => n614);
   U3121 : HS65_LH_IVX9 port map( A => n165, Z => n613);
   U3122 : HS65_LH_IVX9 port map( A => n164, Z => n612);
   U3123 : HS65_LH_IVX9 port map( A => n163, Z => n611);
   U3124 : HS65_LH_IVX9 port map( A => n162, Z => n610);
   U3125 : HS65_LH_IVX9 port map( A => n161, Z => n609);
   U3126 : HS65_LH_IVX9 port map( A => regfile_i(39), Z => n795);
   U3127 : HS65_LH_IVX9 port map( A => regfile_i(38), Z => n811);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity id_top is

   port( clk, rst_n : in std_logic;  id_top_i : in std_logic_vector (71 downto 
         0);  id_top_o : out std_logic_vector (127 downto 0));

end id_top;

architecture SYN_Behavioral of id_top is

   component regfile
      port( clk, rst_n : in std_logic;  regfile_i : in std_logic_vector (49 
            downto 0);  regfile_o : out std_logic_vector (63 downto 0));
   end component;
   
   signal id_top_o_REG_A_31_port, id_top_o_REG_A_30_port, 
      id_top_o_REG_A_29_port, id_top_o_REG_A_28_port, id_top_o_REG_A_27_port, 
      id_top_o_REG_A_26_port, id_top_o_REG_A_25_port, id_top_o_REG_A_24_port, 
      id_top_o_REG_A_23_port, id_top_o_REG_A_22_port, id_top_o_REG_A_21_port, 
      id_top_o_REG_A_20_port, id_top_o_REG_A_19_port, id_top_o_REG_A_18_port, 
      id_top_o_REG_A_17_port, id_top_o_REG_A_16_port, id_top_o_REG_A_15_port, 
      id_top_o_REG_A_14_port, id_top_o_REG_A_13_port, id_top_o_REG_A_12_port, 
      id_top_o_REG_A_11_port, id_top_o_REG_A_10_port, id_top_o_REG_A_9_port, 
      id_top_o_REG_A_8_port, id_top_o_REG_A_7_port, id_top_o_REG_A_6_port, 
      id_top_o_REG_A_5_port, id_top_o_REG_A_4_port, id_top_o_REG_A_3_port, 
      id_top_o_REG_A_2_port, id_top_o_REG_A_1_port, id_top_o_REG_A_0_port, 
      id_top_o_REG_B_31_port, id_top_o_REG_B_30_port, id_top_o_REG_B_29_port, 
      id_top_o_REG_B_28_port, id_top_o_REG_B_27_port, id_top_o_REG_B_26_port, 
      id_top_o_REG_B_25_port, id_top_o_REG_B_24_port, id_top_o_REG_B_23_port, 
      id_top_o_REG_B_22_port, id_top_o_REG_B_21_port, id_top_o_REG_B_20_port, 
      id_top_o_REG_B_19_port, id_top_o_REG_B_18_port, id_top_o_REG_B_17_port, 
      id_top_o_REG_B_16_port, id_top_o_REG_B_15_port, id_top_o_REG_B_14_port, 
      id_top_o_REG_B_13_port, id_top_o_REG_B_12_port, id_top_o_REG_B_11_port, 
      id_top_o_REG_B_10_port, id_top_o_REG_B_9_port, id_top_o_REG_B_8_port, 
      id_top_o_REG_B_7_port, id_top_o_REG_B_6_port, id_top_o_REG_B_5_port, 
      id_top_o_REG_B_4_port, id_top_o_REG_B_3_port, id_top_o_REG_B_2_port, 
      id_top_o_REG_B_1_port, id_top_o_REG_B_0_port : std_logic;

begin
   id_top_o <= ( id_top_o_REG_A_31_port, id_top_o_REG_A_30_port, 
      id_top_o_REG_A_29_port, id_top_o_REG_A_28_port, id_top_o_REG_A_27_port, 
      id_top_o_REG_A_26_port, id_top_o_REG_A_25_port, id_top_o_REG_A_24_port, 
      id_top_o_REG_A_23_port, id_top_o_REG_A_22_port, id_top_o_REG_A_21_port, 
      id_top_o_REG_A_20_port, id_top_o_REG_A_19_port, id_top_o_REG_A_18_port, 
      id_top_o_REG_A_17_port, id_top_o_REG_A_16_port, id_top_o_REG_A_15_port, 
      id_top_o_REG_A_14_port, id_top_o_REG_A_13_port, id_top_o_REG_A_12_port, 
      id_top_o_REG_A_11_port, id_top_o_REG_A_10_port, id_top_o_REG_A_9_port, 
      id_top_o_REG_A_8_port, id_top_o_REG_A_7_port, id_top_o_REG_A_6_port, 
      id_top_o_REG_A_5_port, id_top_o_REG_A_4_port, id_top_o_REG_A_3_port, 
      id_top_o_REG_A_2_port, id_top_o_REG_A_1_port, id_top_o_REG_A_0_port, 
      id_top_o_REG_B_31_port, id_top_o_REG_B_30_port, id_top_o_REG_B_29_port, 
      id_top_o_REG_B_28_port, id_top_o_REG_B_27_port, id_top_o_REG_B_26_port, 
      id_top_o_REG_B_25_port, id_top_o_REG_B_24_port, id_top_o_REG_B_23_port, 
      id_top_o_REG_B_22_port, id_top_o_REG_B_21_port, id_top_o_REG_B_20_port, 
      id_top_o_REG_B_19_port, id_top_o_REG_B_18_port, id_top_o_REG_B_17_port, 
      id_top_o_REG_B_16_port, id_top_o_REG_B_15_port, id_top_o_REG_B_14_port, 
      id_top_o_REG_B_13_port, id_top_o_REG_B_12_port, id_top_o_REG_B_11_port, 
      id_top_o_REG_B_10_port, id_top_o_REG_B_9_port, id_top_o_REG_B_8_port, 
      id_top_o_REG_B_7_port, id_top_o_REG_B_6_port, id_top_o_REG_B_5_port, 
      id_top_o_REG_B_4_port, id_top_o_REG_B_3_port, id_top_o_REG_B_2_port, 
      id_top_o_REG_B_1_port, id_top_o_REG_B_0_port, id_top_i(71), id_top_i(70),
      id_top_i(69), id_top_i(68), id_top_i(67), id_top_i(66), id_top_i(65), 
      id_top_i(64), id_top_i(63), id_top_i(62), id_top_i(61), id_top_i(60), 
      id_top_i(59), id_top_i(58), id_top_i(57), id_top_i(56), id_top_i(55), 
      id_top_i(54), id_top_i(53), id_top_i(52), id_top_i(51), id_top_i(50), 
      id_top_i(49), id_top_i(48), id_top_i(47), id_top_i(46), id_top_i(45), 
      id_top_i(44), id_top_i(43), id_top_i(42), id_top_i(41), id_top_i(40), 
      id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), 
      id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), 
      id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), id_top_i(55), 
      id_top_i(55), id_top_i(55), id_top_i(54), id_top_i(53), id_top_i(52), 
      id_top_i(51), id_top_i(50), id_top_i(49), id_top_i(48), id_top_i(47), 
      id_top_i(46), id_top_i(45), id_top_i(44), id_top_i(43), id_top_i(42), 
      id_top_i(41), id_top_i(40) );
   
   regfile_inst : regfile port map( clk => clk, rst_n => rst_n, regfile_i(49) 
                           => id_top_i(65), regfile_i(48) => id_top_i(64), 
                           regfile_i(47) => id_top_i(63), regfile_i(46) => 
                           id_top_i(62), regfile_i(45) => id_top_i(61), 
                           regfile_i(44) => id_top_i(60), regfile_i(43) => 
                           id_top_i(59), regfile_i(42) => id_top_i(58), 
                           regfile_i(41) => id_top_i(57), regfile_i(40) => 
                           id_top_i(56), regfile_i(39) => id_top_i(4), 
                           regfile_i(38) => id_top_i(3), regfile_i(37) => 
                           id_top_i(2), regfile_i(36) => id_top_i(1), 
                           regfile_i(35) => id_top_i(0), regfile_i(34) => 
                           id_top_i(39), regfile_i(33) => id_top_i(38), 
                           regfile_i(32) => id_top_i(37), regfile_i(31) => 
                           id_top_i(36), regfile_i(30) => id_top_i(35), 
                           regfile_i(29) => id_top_i(34), regfile_i(28) => 
                           id_top_i(33), regfile_i(27) => id_top_i(32), 
                           regfile_i(26) => id_top_i(31), regfile_i(25) => 
                           id_top_i(30), regfile_i(24) => id_top_i(29), 
                           regfile_i(23) => id_top_i(28), regfile_i(22) => 
                           id_top_i(27), regfile_i(21) => id_top_i(26), 
                           regfile_i(20) => id_top_i(25), regfile_i(19) => 
                           id_top_i(24), regfile_i(18) => id_top_i(23), 
                           regfile_i(17) => id_top_i(22), regfile_i(16) => 
                           id_top_i(21), regfile_i(15) => id_top_i(20), 
                           regfile_i(14) => id_top_i(19), regfile_i(13) => 
                           id_top_i(18), regfile_i(12) => id_top_i(17), 
                           regfile_i(11) => id_top_i(16), regfile_i(10) => 
                           id_top_i(15), regfile_i(9) => id_top_i(14), 
                           regfile_i(8) => id_top_i(13), regfile_i(7) => 
                           id_top_i(12), regfile_i(6) => id_top_i(11), 
                           regfile_i(5) => id_top_i(10), regfile_i(4) => 
                           id_top_i(9), regfile_i(3) => id_top_i(8), 
                           regfile_i(2) => id_top_i(7), regfile_i(1) => 
                           id_top_i(6), regfile_i(0) => id_top_i(5), 
                           regfile_o(63) => id_top_o_REG_A_31_port, 
                           regfile_o(62) => id_top_o_REG_A_30_port, 
                           regfile_o(61) => id_top_o_REG_A_29_port, 
                           regfile_o(60) => id_top_o_REG_A_28_port, 
                           regfile_o(59) => id_top_o_REG_A_27_port, 
                           regfile_o(58) => id_top_o_REG_A_26_port, 
                           regfile_o(57) => id_top_o_REG_A_25_port, 
                           regfile_o(56) => id_top_o_REG_A_24_port, 
                           regfile_o(55) => id_top_o_REG_A_23_port, 
                           regfile_o(54) => id_top_o_REG_A_22_port, 
                           regfile_o(53) => id_top_o_REG_A_21_port, 
                           regfile_o(52) => id_top_o_REG_A_20_port, 
                           regfile_o(51) => id_top_o_REG_A_19_port, 
                           regfile_o(50) => id_top_o_REG_A_18_port, 
                           regfile_o(49) => id_top_o_REG_A_17_port, 
                           regfile_o(48) => id_top_o_REG_A_16_port, 
                           regfile_o(47) => id_top_o_REG_A_15_port, 
                           regfile_o(46) => id_top_o_REG_A_14_port, 
                           regfile_o(45) => id_top_o_REG_A_13_port, 
                           regfile_o(44) => id_top_o_REG_A_12_port, 
                           regfile_o(43) => id_top_o_REG_A_11_port, 
                           regfile_o(42) => id_top_o_REG_A_10_port, 
                           regfile_o(41) => id_top_o_REG_A_9_port, 
                           regfile_o(40) => id_top_o_REG_A_8_port, 
                           regfile_o(39) => id_top_o_REG_A_7_port, 
                           regfile_o(38) => id_top_o_REG_A_6_port, 
                           regfile_o(37) => id_top_o_REG_A_5_port, 
                           regfile_o(36) => id_top_o_REG_A_4_port, 
                           regfile_o(35) => id_top_o_REG_A_3_port, 
                           regfile_o(34) => id_top_o_REG_A_2_port, 
                           regfile_o(33) => id_top_o_REG_A_1_port, 
                           regfile_o(32) => id_top_o_REG_A_0_port, 
                           regfile_o(31) => id_top_o_REG_B_31_port, 
                           regfile_o(30) => id_top_o_REG_B_30_port, 
                           regfile_o(29) => id_top_o_REG_B_29_port, 
                           regfile_o(28) => id_top_o_REG_B_28_port, 
                           regfile_o(27) => id_top_o_REG_B_27_port, 
                           regfile_o(26) => id_top_o_REG_B_26_port, 
                           regfile_o(25) => id_top_o_REG_B_25_port, 
                           regfile_o(24) => id_top_o_REG_B_24_port, 
                           regfile_o(23) => id_top_o_REG_B_23_port, 
                           regfile_o(22) => id_top_o_REG_B_22_port, 
                           regfile_o(21) => id_top_o_REG_B_21_port, 
                           regfile_o(20) => id_top_o_REG_B_20_port, 
                           regfile_o(19) => id_top_o_REG_B_19_port, 
                           regfile_o(18) => id_top_o_REG_B_18_port, 
                           regfile_o(17) => id_top_o_REG_B_17_port, 
                           regfile_o(16) => id_top_o_REG_B_16_port, 
                           regfile_o(15) => id_top_o_REG_B_15_port, 
                           regfile_o(14) => id_top_o_REG_B_14_port, 
                           regfile_o(13) => id_top_o_REG_B_13_port, 
                           regfile_o(12) => id_top_o_REG_B_12_port, 
                           regfile_o(11) => id_top_o_REG_B_11_port, 
                           regfile_o(10) => id_top_o_REG_B_10_port, 
                           regfile_o(9) => id_top_o_REG_B_9_port, regfile_o(8) 
                           => id_top_o_REG_B_8_port, regfile_o(7) => 
                           id_top_o_REG_B_7_port, regfile_o(6) => 
                           id_top_o_REG_B_6_port, regfile_o(5) => 
                           id_top_o_REG_B_5_port, regfile_o(4) => 
                           id_top_o_REG_B_4_port, regfile_o(3) => 
                           id_top_o_REG_B_3_port, regfile_o(2) => 
                           id_top_o_REG_B_2_port, regfile_o(1) => 
                           id_top_o_REG_B_1_port, regfile_o(0) => 
                           id_top_o_REG_B_0_port);

end SYN_Behavioral;
