
library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_mult_uns_0 is

   port( a, b : in std_logic_vector (31 downto 0);  product : out 
         std_logic_vector (63 downto 0));

end alu_DW_mult_uns_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_mult_uns_0 is

   component HS65_LHS_XOR2X3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X4
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_HA1X4
      port( A0, B0 : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   signal n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n292, n293, n294, n295, n296, n297, n299, n300, 
      n302, n303, n304, n305, n306, n307, n308, n309, n311, n312, n313, n314, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n330, n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n354, 
      n355, n356, n357, n358, n359, n360, n361, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n385, n386, n387, n388, n389, n390, n391, n392, 
      n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, 
      n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, 
      n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
      n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105 : std_logic
      ;

begin
   
   U228 : HS65_LH_FA1X4 port map( A0 => n293, B0 => n292, CI => n228, CO => 
                           n227, S0 => product(62));
   U229 : HS65_LH_FA1X4 port map( A0 => n295, B0 => n294, CI => n229, CO => 
                           n228, S0 => product(61));
   U230 : HS65_LH_FA1X4 port map( A0 => n296, B0 => n299, CI => n230, CO => 
                           n229, S0 => product(60));
   U231 : HS65_LH_FA1X4 port map( A0 => n300, B0 => n302, CI => n231, CO => 
                           n230, S0 => product(59));
   U232 : HS65_LH_FA1X4 port map( A0 => n303, B0 => n305, CI => n232, CO => 
                           n231, S0 => product(58));
   U233 : HS65_LH_FA1X4 port map( A0 => n306, B0 => n311, CI => n233, CO => 
                           n232, S0 => product(57));
   U234 : HS65_LH_FA1X4 port map( A0 => n312, B0 => n316, CI => n234, CO => 
                           n233, S0 => product(56));
   U235 : HS65_LH_FA1X4 port map( A0 => n317, B0 => n322, CI => n235, CO => 
                           n234, S0 => product(55));
   U236 : HS65_LH_FA1X4 port map( A0 => n323, B0 => n330, CI => n236, CO => 
                           n235, S0 => product(54));
   U237 : HS65_LH_FA1X4 port map( A0 => n331, B0 => n337, CI => n237, CO => 
                           n236, S0 => product(53));
   U238 : HS65_LH_FA1X4 port map( A0 => n338, B0 => n344, CI => n238, CO => 
                           n237, S0 => product(52));
   U239 : HS65_LH_FA1X4 port map( A0 => n345, B0 => n354, CI => n239, CO => 
                           n238, S0 => product(51));
   U240 : HS65_LH_FA1X4 port map( A0 => n355, B0 => n363, CI => n240, CO => 
                           n239, S0 => product(50));
   U241 : HS65_LH_FA1X4 port map( A0 => n364, B0 => n373, CI => n241, CO => 
                           n240, S0 => product(49));
   U242 : HS65_LH_FA1X4 port map( A0 => n374, B0 => n385, CI => n242, CO => 
                           n241, S0 => product(48));
   U243 : HS65_LH_FA1X4 port map( A0 => n386, B0 => n396, CI => n243, CO => 
                           n242, S0 => product(47));
   U244 : HS65_LH_FA1X4 port map( A0 => n397, B0 => n407, CI => n244, CO => 
                           n243, S0 => product(46));
   U245 : HS65_LH_FA1X4 port map( A0 => n408, B0 => n421, CI => n245, CO => 
                           n244, S0 => product(45));
   U246 : HS65_LH_FA1X4 port map( A0 => n422, B0 => n434, CI => n246, CO => 
                           n245, S0 => product(44));
   U247 : HS65_LH_FA1X4 port map( A0 => n435, B0 => n448, CI => n247, CO => 
                           n246, S0 => product(43));
   U248 : HS65_LH_FA1X4 port map( A0 => n449, B0 => n464, CI => n248, CO => 
                           n247, S0 => product(42));
   U249 : HS65_LH_FA1X4 port map( A0 => n465, B0 => n479, CI => n249, CO => 
                           n248, S0 => product(41));
   U250 : HS65_LH_FA1X4 port map( A0 => n480, B0 => n494, CI => n250, CO => 
                           n249, S0 => product(40));
   U251 : HS65_LH_FA1X4 port map( A0 => n495, B0 => n512, CI => n251, CO => 
                           n250, S0 => product(39));
   U252 : HS65_LH_FA1X4 port map( A0 => n513, B0 => n529, CI => n252, CO => 
                           n251, S0 => product(38));
   U253 : HS65_LH_FA1X4 port map( A0 => n530, B0 => n546, CI => n253, CO => 
                           n252, S0 => product(37));
   U254 : HS65_LH_FA1X4 port map( A0 => n547, B0 => n564, CI => n254, CO => 
                           n253, S0 => product(36));
   U255 : HS65_LH_FA1X4 port map( A0 => n565, B0 => n582, CI => n255, CO => 
                           n254, S0 => product(35));
   U256 : HS65_LH_FA1X4 port map( A0 => n583, B0 => n600, CI => n256, CO => 
                           n255, S0 => product(34));
   U257 : HS65_LH_FA1X4 port map( A0 => n601, B0 => n1386, CI => n257, CO => 
                           n256, S0 => product(33));
   U258 : HS65_LH_FA1X4 port map( A0 => n1387, B0 => n619, CI => n258, CO => 
                           n257, S0 => product(32));
   U259 : HS65_LH_FA1X4 port map( A0 => n1388, B0 => n637, CI => n259, CO => 
                           n258, S0 => product(31));
   U260 : HS65_LH_FA1X4 port map( A0 => n1389, B0 => n655, CI => n260, CO => 
                           n259, S0 => product(30));
   U261 : HS65_LH_FA1X4 port map( A0 => n1390, B0 => n673, CI => n261, CO => 
                           n260, S0 => product(29));
   U262 : HS65_LH_FA1X4 port map( A0 => n1391, B0 => n691, CI => n262, CO => 
                           n261, S0 => product(28));
   U263 : HS65_LH_FA1X4 port map( A0 => n1392, B0 => n709, CI => n263, CO => 
                           n262, S0 => product(27));
   U264 : HS65_LH_FA1X4 port map( A0 => n1393, B0 => n727, CI => n264, CO => 
                           n263, S0 => product(26));
   U265 : HS65_LH_FA1X4 port map( A0 => n1394, B0 => n743, CI => n265, CO => 
                           n264, S0 => product(25));
   U266 : HS65_LH_FA1X4 port map( A0 => n1395, B0 => n759, CI => n266, CO => 
                           n265, S0 => product(24));
   U267 : HS65_LH_FA1X4 port map( A0 => n1396, B0 => n775, CI => n267, CO => 
                           n266, S0 => product(23));
   U268 : HS65_LH_FA1X4 port map( A0 => n1397, B0 => n789, CI => n268, CO => 
                           n267, S0 => product(22));
   U269 : HS65_LH_FA1X4 port map( A0 => n1398, B0 => n803, CI => n269, CO => 
                           n268, S0 => product(21));
   U270 : HS65_LH_FA1X4 port map( A0 => n1399, B0 => n817, CI => n270, CO => 
                           n269, S0 => product(20));
   U271 : HS65_LH_FA1X4 port map( A0 => n1400, B0 => n829, CI => n271, CO => 
                           n270, S0 => product(19));
   U272 : HS65_LH_FA1X4 port map( A0 => n1401, B0 => n841, CI => n272, CO => 
                           n271, S0 => product(18));
   U273 : HS65_LH_FA1X4 port map( A0 => n1402, B0 => n853, CI => n273, CO => 
                           n272, S0 => product(17));
   U274 : HS65_LH_FA1X4 port map( A0 => n1403, B0 => n863, CI => n274, CO => 
                           n273, S0 => product(16));
   U275 : HS65_LH_FA1X4 port map( A0 => n1404, B0 => n873, CI => n275, CO => 
                           n274, S0 => product(15));
   U276 : HS65_LH_FA1X4 port map( A0 => n1405, B0 => n883, CI => n276, CO => 
                           n275, S0 => product(14));
   U277 : HS65_LH_FA1X4 port map( A0 => n1406, B0 => n891, CI => n277, CO => 
                           n276, S0 => product(13));
   U278 : HS65_LH_FA1X4 port map( A0 => n1407, B0 => n899, CI => n278, CO => 
                           n277, S0 => product(12));
   U279 : HS65_LH_FA1X4 port map( A0 => n1408, B0 => n907, CI => n279, CO => 
                           n278, S0 => product(11));
   U280 : HS65_LH_FA1X4 port map( A0 => n1409, B0 => n913, CI => n280, CO => 
                           n279, S0 => product(10));
   U281 : HS65_LH_FA1X4 port map( A0 => n1410, B0 => n919, CI => n281, CO => 
                           n280, S0 => product(9));
   U282 : HS65_LH_FA1X4 port map( A0 => n1411, B0 => n925, CI => n282, CO => 
                           n281, S0 => product(8));
   U283 : HS65_LH_FA1X4 port map( A0 => n1412, B0 => n929, CI => n283, CO => 
                           n282, S0 => product(7));
   U284 : HS65_LH_FA1X4 port map( A0 => n1413, B0 => n933, CI => n284, CO => 
                           n283, S0 => product(6));
   U285 : HS65_LH_FA1X4 port map( A0 => n1414, B0 => n937, CI => n285, CO => 
                           n284, S0 => product(5));
   U286 : HS65_LH_FA1X4 port map( A0 => n1415, B0 => n939, CI => n286, CO => 
                           n285, S0 => product(4));
   U287 : HS65_LH_FA1X4 port map( A0 => n1416, B0 => n941, CI => n287, CO => 
                           n286, S0 => product(3));
   U288 : HS65_LH_HA1X4 port map( A0 => n1417, B0 => n288, CO => n287, S0 => 
                           product(2));
   U289 : HS65_LH_HA1X4 port map( A0 => n1418, B0 => n289, CO => n288, S0 => 
                           product(1));
   U290 : HS65_LH_HA1X4 port map( A0 => n2629, B0 => n1419, CO => n289, S0 => 
                           product(0));
   U293 : HS65_LH_FA1X4 port map( A0 => n297, B0 => n2657, CI => n1041, CO => 
                           n293, S0 => n294);
   U294 : HS65_LH_FA1X4 port map( A0 => n1042, B0 => n2658, CI => n1071, CO => 
                           n295, S0 => n296);
   U296 : HS65_LH_FA1X4 port map( A0 => n2658, B0 => n1043, CI => n1072, CO => 
                           n299, S0 => n300);
   U298 : HS65_LH_FA1X4 port map( A0 => n1073, B0 => n304, CI => n307, CO => 
                           n302, S0 => n303);
   U299 : HS65_LH_FA1X4 port map( A0 => n309, B0 => n2654, CI => n1044, CO => 
                           n297, S0 => n304);
   U300 : HS65_LH_FA1X4 port map( A0 => n1106, B0 => n1074, CI => n308, CO => 
                           n305, S0 => n306);
   U301 : HS65_LH_FA1X4 port map( A0 => n1045, B0 => n2663, CI => n313, CO => 
                           n307, S0 => n308);
   U303 : HS65_LH_FA1X4 port map( A0 => n314, B0 => n318, CI => n1107, CO => 
                           n311, S0 => n312);
   U304 : HS65_LH_FA1X4 port map( A0 => n2663, B0 => n320, CI => n1075, CO => 
                           n313, S0 => n314);
   U306 : HS65_LH_FA1X4 port map( A0 => n1108, B0 => n319, CI => n324, CO => 
                           n316, S0 => n317);
   U307 : HS65_LH_FA1X4 port map( A0 => n326, B0 => n321, CI => n1076, CO => 
                           n318, S0 => n319);
   U308 : HS65_LH_FA1X4 port map( A0 => n328, B0 => n2651, CI => n1046, CO => 
                           n320, S0 => n321);
   U309 : HS65_LH_FA1X4 port map( A0 => n1141, B0 => n1109, CI => n325, CO => 
                           n322, S0 => n323);
   U310 : HS65_LH_FA1X4 port map( A0 => n327, B0 => n334, CI => n332, CO => 
                           n324, S0 => n325);
   U311 : HS65_LH_FA1X4 port map( A0 => n1047, B0 => n2659, CI => n1077, CO => 
                           n326, S0 => n327);
   U313 : HS65_LH_FA1X4 port map( A0 => n333, B0 => n339, CI => n1142, CO => 
                           n330, S0 => n331);
   U314 : HS65_LH_FA1X4 port map( A0 => n335, B0 => n341, CI => n1110, CO => 
                           n332, S0 => n333);
   U315 : HS65_LH_FA1X4 port map( A0 => n2659, B0 => n1048, CI => n1078, CO => 
                           n334, S0 => n335);
   U317 : HS65_LH_FA1X4 port map( A0 => n1143, B0 => n340, CI => n346, CO => 
                           n337, S0 => n338);
   U318 : HS65_LH_FA1X4 port map( A0 => n348, B0 => n342, CI => n1111, CO => 
                           n339, S0 => n340);
   U319 : HS65_LH_FA1X4 port map( A0 => n1079, B0 => n343, CI => n350, CO => 
                           n341, S0 => n342);
   U320 : HS65_LH_FA1X4 port map( A0 => n352, B0 => n2648, CI => n1049, CO => 
                           n328, S0 => n343);
   U321 : HS65_LH_FA1X4 port map( A0 => n1176, B0 => n1144, CI => n347, CO => 
                           n344, S0 => n345);
   U322 : HS65_LH_FA1X4 port map( A0 => n349, B0 => n358, CI => n356, CO => 
                           n346, S0 => n347);
   U323 : HS65_LH_FA1X4 port map( A0 => n351, B0 => n1080, CI => n1112, CO => 
                           n348, S0 => n349);
   U324 : HS65_LH_FA1X4 port map( A0 => n1050, B0 => n2664, CI => n360, CO => 
                           n350, S0 => n351);
   U326 : HS65_LH_FA1X4 port map( A0 => n357, B0 => n365, CI => n1177, CO => 
                           n354, S0 => n355);
   U327 : HS65_LH_FA1X4 port map( A0 => n359, B0 => n367, CI => n1145, CO => 
                           n356, S0 => n357);
   U328 : HS65_LH_FA1X4 port map( A0 => n361, B0 => n369, CI => n1113, CO => 
                           n358, S0 => n359);
   U329 : HS65_LH_FA1X4 port map( A0 => n2664, B0 => n371, CI => n1081, CO => 
                           n360, S0 => n361);
   U331 : HS65_LH_FA1X4 port map( A0 => n1178, B0 => n366, CI => n375, CO => 
                           n363, S0 => n364);
   U332 : HS65_LH_FA1X4 port map( A0 => n377, B0 => n368, CI => n1146, CO => 
                           n365, S0 => n366);
   U333 : HS65_LH_FA1X4 port map( A0 => n1114, B0 => n370, CI => n379, CO => 
                           n367, S0 => n368);
   U334 : HS65_LH_FA1X4 port map( A0 => n381, B0 => n372, CI => n1082, CO => 
                           n369, S0 => n370);
   U335 : HS65_LH_FA1X4 port map( A0 => n383, B0 => n2645, CI => n1051, CO => 
                           n371, S0 => n372);
   U336 : HS65_LH_FA1X4 port map( A0 => n1211, B0 => n1179, CI => n376, CO => 
                           n373, S0 => n374);
   U337 : HS65_LH_FA1X4 port map( A0 => n378, B0 => n389, CI => n387, CO => 
                           n375, S0 => n376);
   U338 : HS65_LH_FA1X4 port map( A0 => n380, B0 => n1115, CI => n1147, CO => 
                           n377, S0 => n378);
   U339 : HS65_LH_FA1X4 port map( A0 => n382, B0 => n393, CI => n391, CO => 
                           n379, S0 => n380);
   U340 : HS65_LH_FA1X4 port map( A0 => n1052, B0 => n2660, CI => n1083, CO => 
                           n381, S0 => n382);
   U342 : HS65_LH_FA1X4 port map( A0 => n388, B0 => n398, CI => n1212, CO => 
                           n385, S0 => n386);
   U343 : HS65_LH_FA1X4 port map( A0 => n390, B0 => n400, CI => n1180, CO => 
                           n387, S0 => n388);
   U344 : HS65_LH_FA1X4 port map( A0 => n392, B0 => n402, CI => n1148, CO => 
                           n389, S0 => n390);
   U345 : HS65_LH_FA1X4 port map( A0 => n394, B0 => n404, CI => n1116, CO => 
                           n391, S0 => n392);
   U346 : HS65_LH_FA1X4 port map( A0 => n2660, B0 => n1053, CI => n1084, CO => 
                           n393, S0 => n394);
   U348 : HS65_LH_FA1X4 port map( A0 => n1213, B0 => n399, CI => n409, CO => 
                           n396, S0 => n397);
   U349 : HS65_LH_FA1X4 port map( A0 => n411, B0 => n401, CI => n1181, CO => 
                           n398, S0 => n399);
   U350 : HS65_LH_FA1X4 port map( A0 => n1149, B0 => n403, CI => n413, CO => 
                           n400, S0 => n401);
   U351 : HS65_LH_FA1X4 port map( A0 => n415, B0 => n405, CI => n1117, CO => 
                           n402, S0 => n403);
   U352 : HS65_LH_FA1X4 port map( A0 => n1085, B0 => n406, CI => n417, CO => 
                           n404, S0 => n405);
   U353 : HS65_LH_FA1X4 port map( A0 => n419, B0 => n2642, CI => n1054, CO => 
                           n383, S0 => n406);
   U354 : HS65_LH_FA1X4 port map( A0 => n1246, B0 => n1214, CI => n410, CO => 
                           n407, S0 => n408);
   U355 : HS65_LH_FA1X4 port map( A0 => n412, B0 => n425, CI => n423, CO => 
                           n409, S0 => n410);
   U356 : HS65_LH_FA1X4 port map( A0 => n414, B0 => n1150, CI => n1182, CO => 
                           n411, S0 => n412);
   U357 : HS65_LH_FA1X4 port map( A0 => n416, B0 => n429, CI => n427, CO => 
                           n413, S0 => n414);
   U358 : HS65_LH_FA1X4 port map( A0 => n418, B0 => n1086, CI => n1118, CO => 
                           n415, S0 => n416);
   U359 : HS65_LH_FA1X4 port map( A0 => n1055, B0 => n2665, CI => n431, CO => 
                           n417, S0 => n418);
   U361 : HS65_LH_FA1X4 port map( A0 => n424, B0 => n436, CI => n1247, CO => 
                           n421, S0 => n422);
   U362 : HS65_LH_FA1X4 port map( A0 => n426, B0 => n438, CI => n1215, CO => 
                           n423, S0 => n424);
   U363 : HS65_LH_FA1X4 port map( A0 => n428, B0 => n440, CI => n1183, CO => 
                           n425, S0 => n426);
   U364 : HS65_LH_FA1X4 port map( A0 => n430, B0 => n442, CI => n1151, CO => 
                           n427, S0 => n428);
   U365 : HS65_LH_FA1X4 port map( A0 => n432, B0 => n444, CI => n1119, CO => 
                           n429, S0 => n430);
   U366 : HS65_LH_FA1X4 port map( A0 => n2665, B0 => n446, CI => n1087, CO => 
                           n431, S0 => n432);
   U368 : HS65_LH_FA1X4 port map( A0 => n1248, B0 => n437, CI => n450, CO => 
                           n434, S0 => n435);
   U369 : HS65_LH_FA1X4 port map( A0 => n452, B0 => n439, CI => n1216, CO => 
                           n436, S0 => n437);
   U370 : HS65_LH_FA1X4 port map( A0 => n1184, B0 => n441, CI => n454, CO => 
                           n438, S0 => n439);
   U371 : HS65_LH_FA1X4 port map( A0 => n456, B0 => n443, CI => n1152, CO => 
                           n440, S0 => n441);
   U372 : HS65_LH_FA1X4 port map( A0 => n1120, B0 => n445, CI => n458, CO => 
                           n442, S0 => n443);
   U373 : HS65_LH_FA1X4 port map( A0 => n460, B0 => n447, CI => n1088, CO => 
                           n444, S0 => n445);
   U374 : HS65_LH_FA1X4 port map( A0 => n462, B0 => n2639, CI => n1056, CO => 
                           n446, S0 => n447);
   U375 : HS65_LH_FA1X4 port map( A0 => n1281, B0 => n1249, CI => n451, CO => 
                           n448, S0 => n449);
   U376 : HS65_LH_FA1X4 port map( A0 => n453, B0 => n468, CI => n466, CO => 
                           n450, S0 => n451);
   U377 : HS65_LH_FA1X4 port map( A0 => n455, B0 => n1185, CI => n1217, CO => 
                           n452, S0 => n453);
   U378 : HS65_LH_FA1X4 port map( A0 => n457, B0 => n472, CI => n470, CO => 
                           n454, S0 => n455);
   U379 : HS65_LH_FA1X4 port map( A0 => n459, B0 => n1121, CI => n1153, CO => 
                           n456, S0 => n457);
   U380 : HS65_LH_FA1X4 port map( A0 => n461, B0 => n476, CI => n474, CO => 
                           n458, S0 => n459);
   U381 : HS65_LH_FA1X4 port map( A0 => n1057, B0 => n2661, CI => n1089, CO => 
                           n460, S0 => n461);
   U383 : HS65_LH_FA1X4 port map( A0 => n467, B0 => n481, CI => n1282, CO => 
                           n464, S0 => n465);
   U384 : HS65_LH_FA1X4 port map( A0 => n469, B0 => n483, CI => n1250, CO => 
                           n466, S0 => n467);
   U385 : HS65_LH_FA1X4 port map( A0 => n471, B0 => n485, CI => n1218, CO => 
                           n468, S0 => n469);
   U386 : HS65_LH_FA1X4 port map( A0 => n473, B0 => n487, CI => n1186, CO => 
                           n470, S0 => n471);
   U387 : HS65_LH_FA1X4 port map( A0 => n475, B0 => n489, CI => n1154, CO => 
                           n472, S0 => n473);
   U388 : HS65_LH_FA1X4 port map( A0 => n477, B0 => n491, CI => n1122, CO => 
                           n474, S0 => n475);
   U389 : HS65_LH_FA1X4 port map( A0 => n2661, B0 => n1058, CI => n1090, CO => 
                           n476, S0 => n477);
   U391 : HS65_LH_FA1X4 port map( A0 => n1283, B0 => n482, CI => n496, CO => 
                           n479, S0 => n480);
   U392 : HS65_LH_FA1X4 port map( A0 => n498, B0 => n484, CI => n1251, CO => 
                           n481, S0 => n482);
   U393 : HS65_LH_FA1X4 port map( A0 => n1219, B0 => n486, CI => n500, CO => 
                           n483, S0 => n484);
   U394 : HS65_LH_FA1X4 port map( A0 => n502, B0 => n488, CI => n1187, CO => 
                           n485, S0 => n486);
   U395 : HS65_LH_FA1X4 port map( A0 => n1155, B0 => n490, CI => n504, CO => 
                           n487, S0 => n488);
   U396 : HS65_LH_FA1X4 port map( A0 => n506, B0 => n492, CI => n1123, CO => 
                           n489, S0 => n490);
   U397 : HS65_LH_FA1X4 port map( A0 => n1091, B0 => n493, CI => n508, CO => 
                           n491, S0 => n492);
   U398 : HS65_LH_FA1X4 port map( A0 => n510, B0 => n2636, CI => n1059, CO => 
                           n462, S0 => n493);
   U399 : HS65_LH_FA1X4 port map( A0 => n1316, B0 => n1284, CI => n497, CO => 
                           n494, S0 => n495);
   U400 : HS65_LH_FA1X4 port map( A0 => n499, B0 => n516, CI => n514, CO => 
                           n496, S0 => n497);
   U401 : HS65_LH_FA1X4 port map( A0 => n501, B0 => n1220, CI => n1252, CO => 
                           n498, S0 => n499);
   U402 : HS65_LH_FA1X4 port map( A0 => n503, B0 => n520, CI => n518, CO => 
                           n500, S0 => n501);
   U403 : HS65_LH_FA1X4 port map( A0 => n505, B0 => n1156, CI => n1188, CO => 
                           n502, S0 => n503);
   U404 : HS65_LH_FA1X4 port map( A0 => n507, B0 => n524, CI => n522, CO => 
                           n504, S0 => n505);
   U405 : HS65_LH_FA1X4 port map( A0 => n509, B0 => n1092, CI => n1124, CO => 
                           n506, S0 => n507);
   U406 : HS65_LH_FA1X4 port map( A0 => n1060, B0 => n2662, CI => n526, CO => 
                           n508, S0 => n509);
   U408 : HS65_LH_FA1X4 port map( A0 => n515, B0 => n531, CI => n1317, CO => 
                           n512, S0 => n513);
   U409 : HS65_LH_FA1X4 port map( A0 => n517, B0 => n533, CI => n1285, CO => 
                           n514, S0 => n515);
   U410 : HS65_LH_FA1X4 port map( A0 => n519, B0 => n535, CI => n1253, CO => 
                           n516, S0 => n517);
   U411 : HS65_LH_FA1X4 port map( A0 => n521, B0 => n537, CI => n1221, CO => 
                           n518, S0 => n519);
   U412 : HS65_LH_FA1X4 port map( A0 => n523, B0 => n539, CI => n1189, CO => 
                           n520, S0 => n521);
   U413 : HS65_LH_FA1X4 port map( A0 => n525, B0 => n541, CI => n1157, CO => 
                           n522, S0 => n523);
   U414 : HS65_LH_FA1X4 port map( A0 => n527, B0 => n543, CI => n1125, CO => 
                           n524, S0 => n525);
   U415 : HS65_LH_FA1X4 port map( A0 => n2662, B0 => n1061, CI => n1093, CO => 
                           n526, S0 => n527);
   U417 : HS65_LH_FA1X4 port map( A0 => n1318, B0 => n532, CI => n548, CO => 
                           n529, S0 => n530);
   U418 : HS65_LH_FA1X4 port map( A0 => n550, B0 => n534, CI => n1286, CO => 
                           n531, S0 => n532);
   U419 : HS65_LH_FA1X4 port map( A0 => n1254, B0 => n536, CI => n552, CO => 
                           n533, S0 => n534);
   U420 : HS65_LH_FA1X4 port map( A0 => n554, B0 => n538, CI => n1222, CO => 
                           n535, S0 => n536);
   U421 : HS65_LH_FA1X4 port map( A0 => n1190, B0 => n540, CI => n556, CO => 
                           n537, S0 => n538);
   U422 : HS65_LH_FA1X4 port map( A0 => n1158, B0 => n542, CI => n558, CO => 
                           n539, S0 => n540);
   U423 : HS65_LH_FA1X4 port map( A0 => n1126, B0 => n544, CI => n560, CO => 
                           n541, S0 => n542);
   U424 : HS65_LH_FA1X4 port map( A0 => n562, B0 => n545, CI => n1094, CO => 
                           n543, S0 => n544);
   U425 : HS65_LH_FA1X4 port map( A0 => n2633, B0 => n2630, CI => n1062, CO => 
                           n510, S0 => n545);
   U426 : HS65_LH_FA1X4 port map( A0 => n1351, B0 => n1319, CI => n549, CO => 
                           n546, S0 => n547);
   U427 : HS65_LH_FA1X4 port map( A0 => n551, B0 => n1287, CI => n566, CO => 
                           n548, S0 => n549);
   U428 : HS65_LH_FA1X4 port map( A0 => n553, B0 => n1255, CI => n568, CO => 
                           n550, S0 => n551);
   U429 : HS65_LH_FA1X4 port map( A0 => n555, B0 => n572, CI => n570, CO => 
                           n552, S0 => n553);
   U430 : HS65_LH_FA1X4 port map( A0 => n557, B0 => n1191, CI => n1223, CO => 
                           n554, S0 => n555);
   U431 : HS65_LH_FA1X4 port map( A0 => n559, B0 => n576, CI => n574, CO => 
                           n556, S0 => n557);
   U432 : HS65_LH_FA1X4 port map( A0 => n561, B0 => n1127, CI => n1159, CO => 
                           n558, S0 => n559);
   U433 : HS65_LH_FA1X4 port map( A0 => n563, B0 => n1095, CI => n578, CO => 
                           n560, S0 => n561);
   U434 : HS65_LH_FA1X4 port map( A0 => n1063, B0 => n2628, CI => n580, CO => 
                           n562, S0 => n563);
   U435 : HS65_LH_FA1X4 port map( A0 => n567, B0 => n1320, CI => n1352, CO => 
                           n564, S0 => n565);
   U436 : HS65_LH_FA1X4 port map( A0 => n569, B0 => n1288, CI => n584, CO => 
                           n566, S0 => n567);
   U437 : HS65_LH_FA1X4 port map( A0 => n571, B0 => n1256, CI => n586, CO => 
                           n568, S0 => n569);
   U438 : HS65_LH_FA1X4 port map( A0 => n573, B0 => n590, CI => n588, CO => 
                           n570, S0 => n571);
   U439 : HS65_LH_FA1X4 port map( A0 => n575, B0 => n1192, CI => n1224, CO => 
                           n572, S0 => n573);
   U440 : HS65_LH_FA1X4 port map( A0 => n577, B0 => n594, CI => n592, CO => 
                           n574, S0 => n575);
   U441 : HS65_LH_FA1X4 port map( A0 => n579, B0 => n1128, CI => n1160, CO => 
                           n576, S0 => n577);
   U442 : HS65_LH_FA1X4 port map( A0 => n581, B0 => n1096, CI => n596, CO => 
                           n578, S0 => n579);
   U443 : HS65_LH_FA1X4 port map( A0 => n1064, B0 => n2628, CI => n598, CO => 
                           n580, S0 => n581);
   U444 : HS65_LH_FA1X4 port map( A0 => n585, B0 => n602, CI => n1353, CO => 
                           n582, S0 => n583);
   U445 : HS65_LH_FA1X4 port map( A0 => n587, B0 => n604, CI => n1321, CO => 
                           n584, S0 => n585);
   U446 : HS65_LH_FA1X4 port map( A0 => n589, B0 => n606, CI => n1289, CO => 
                           n586, S0 => n587);
   U447 : HS65_LH_FA1X4 port map( A0 => n591, B0 => n608, CI => n1257, CO => 
                           n588, S0 => n589);
   U448 : HS65_LH_FA1X4 port map( A0 => n593, B0 => n610, CI => n1225, CO => 
                           n590, S0 => n591);
   U449 : HS65_LH_FA1X4 port map( A0 => n595, B0 => n612, CI => n1193, CO => 
                           n592, S0 => n593);
   U450 : HS65_LH_FA1X4 port map( A0 => n597, B0 => n614, CI => n1161, CO => 
                           n594, S0 => n595);
   U451 : HS65_LH_FA1X4 port map( A0 => n599, B0 => n616, CI => n1129, CO => 
                           n596, S0 => n597);
   U452 : HS65_LH_FA1X4 port map( A0 => n1065, B0 => n2628, CI => n1097, CO => 
                           n598, S0 => n599);
   U453 : HS65_LH_FA1X4 port map( A0 => n1354, B0 => n603, CI => n618, CO => 
                           n600, S0 => n601);
   U454 : HS65_LH_FA1X4 port map( A0 => n1322, B0 => n605, CI => n620, CO => 
                           n602, S0 => n603);
   U455 : HS65_LH_FA1X4 port map( A0 => n1290, B0 => n607, CI => n622, CO => 
                           n604, S0 => n605);
   U456 : HS65_LH_FA1X4 port map( A0 => n1258, B0 => n609, CI => n624, CO => 
                           n606, S0 => n607);
   U457 : HS65_LH_FA1X4 port map( A0 => n1226, B0 => n611, CI => n626, CO => 
                           n608, S0 => n609);
   U458 : HS65_LH_FA1X4 port map( A0 => n1194, B0 => n613, CI => n628, CO => 
                           n610, S0 => n611);
   U459 : HS65_LH_FA1X4 port map( A0 => n1162, B0 => n615, CI => n630, CO => 
                           n612, S0 => n613);
   U460 : HS65_LH_FA1X4 port map( A0 => n1130, B0 => n617, CI => n632, CO => 
                           n614, S0 => n615);
   U461 : HS65_LH_FA1X4 port map( A0 => n1098, B0 => n1066, CI => n634, CO => 
                           n616, S0 => n617);
   U462 : HS65_LH_FA1X4 port map( A0 => n1355, B0 => n621, CI => n636, CO => 
                           n618, S0 => n619);
   U463 : HS65_LH_FA1X4 port map( A0 => n1323, B0 => n623, CI => n638, CO => 
                           n620, S0 => n621);
   U464 : HS65_LH_FA1X4 port map( A0 => n1291, B0 => n625, CI => n640, CO => 
                           n622, S0 => n623);
   U465 : HS65_LH_FA1X4 port map( A0 => n1259, B0 => n627, CI => n642, CO => 
                           n624, S0 => n625);
   U466 : HS65_LH_FA1X4 port map( A0 => n1227, B0 => n629, CI => n644, CO => 
                           n626, S0 => n627);
   U467 : HS65_LH_FA1X4 port map( A0 => n1195, B0 => n631, CI => n646, CO => 
                           n628, S0 => n629);
   U468 : HS65_LH_FA1X4 port map( A0 => n1163, B0 => n633, CI => n648, CO => 
                           n630, S0 => n631);
   U469 : HS65_LH_FA1X4 port map( A0 => n1131, B0 => n635, CI => n650, CO => 
                           n632, S0 => n633);
   U470 : HS65_LH_FA1X4 port map( A0 => n1099, B0 => n1067, CI => n652, CO => 
                           n634, S0 => n635);
   U471 : HS65_LH_FA1X4 port map( A0 => n1356, B0 => n639, CI => n654, CO => 
                           n636, S0 => n637);
   U472 : HS65_LH_FA1X4 port map( A0 => n1324, B0 => n641, CI => n656, CO => 
                           n638, S0 => n639);
   U473 : HS65_LH_FA1X4 port map( A0 => n1292, B0 => n643, CI => n658, CO => 
                           n640, S0 => n641);
   U474 : HS65_LH_FA1X4 port map( A0 => n1260, B0 => n645, CI => n660, CO => 
                           n642, S0 => n643);
   U475 : HS65_LH_FA1X4 port map( A0 => n1228, B0 => n647, CI => n662, CO => 
                           n644, S0 => n645);
   U476 : HS65_LH_FA1X4 port map( A0 => n1196, B0 => n649, CI => n664, CO => 
                           n646, S0 => n647);
   U477 : HS65_LH_FA1X4 port map( A0 => n1164, B0 => n651, CI => n666, CO => 
                           n648, S0 => n649);
   U478 : HS65_LH_FA1X4 port map( A0 => n1132, B0 => n653, CI => n668, CO => 
                           n650, S0 => n651);
   U479 : HS65_LH_FA1X4 port map( A0 => n1100, B0 => n1068, CI => n670, CO => 
                           n652, S0 => n653);
   U480 : HS65_LH_FA1X4 port map( A0 => n1357, B0 => n657, CI => n672, CO => 
                           n654, S0 => n655);
   U481 : HS65_LH_FA1X4 port map( A0 => n1325, B0 => n659, CI => n674, CO => 
                           n656, S0 => n657);
   U482 : HS65_LH_FA1X4 port map( A0 => n1293, B0 => n661, CI => n676, CO => 
                           n658, S0 => n659);
   U483 : HS65_LH_FA1X4 port map( A0 => n1261, B0 => n663, CI => n678, CO => 
                           n660, S0 => n661);
   U484 : HS65_LH_FA1X4 port map( A0 => n1229, B0 => n665, CI => n680, CO => 
                           n662, S0 => n663);
   U485 : HS65_LH_FA1X4 port map( A0 => n1197, B0 => n667, CI => n682, CO => 
                           n664, S0 => n665);
   U486 : HS65_LH_FA1X4 port map( A0 => n1165, B0 => n669, CI => n684, CO => 
                           n666, S0 => n667);
   U487 : HS65_LH_FA1X4 port map( A0 => n1133, B0 => n671, CI => n686, CO => 
                           n668, S0 => n669);
   U488 : HS65_LH_FA1X4 port map( A0 => n1101, B0 => n1069, CI => n688, CO => 
                           n670, S0 => n671);
   U489 : HS65_LH_FA1X4 port map( A0 => n1358, B0 => n675, CI => n690, CO => 
                           n672, S0 => n673);
   U490 : HS65_LH_FA1X4 port map( A0 => n1326, B0 => n677, CI => n692, CO => 
                           n674, S0 => n675);
   U491 : HS65_LH_FA1X4 port map( A0 => n1294, B0 => n679, CI => n694, CO => 
                           n676, S0 => n677);
   U492 : HS65_LH_FA1X4 port map( A0 => n1262, B0 => n681, CI => n696, CO => 
                           n678, S0 => n679);
   U493 : HS65_LH_FA1X4 port map( A0 => n1230, B0 => n683, CI => n698, CO => 
                           n680, S0 => n681);
   U494 : HS65_LH_FA1X4 port map( A0 => n1198, B0 => n685, CI => n700, CO => 
                           n682, S0 => n683);
   U495 : HS65_LH_FA1X4 port map( A0 => n1166, B0 => n687, CI => n702, CO => 
                           n684, S0 => n685);
   U496 : HS65_LH_FA1X4 port map( A0 => n1134, B0 => n689, CI => n704, CO => 
                           n686, S0 => n687);
   U497 : HS65_LH_HA1X4 port map( A0 => n1102, B0 => n706, CO => n688, S0 => 
                           n689);
   U498 : HS65_LH_FA1X4 port map( A0 => n1359, B0 => n693, CI => n708, CO => 
                           n690, S0 => n691);
   U499 : HS65_LH_FA1X4 port map( A0 => n1327, B0 => n695, CI => n710, CO => 
                           n692, S0 => n693);
   U500 : HS65_LH_FA1X4 port map( A0 => n1295, B0 => n697, CI => n712, CO => 
                           n694, S0 => n695);
   U501 : HS65_LH_FA1X4 port map( A0 => n1263, B0 => n699, CI => n714, CO => 
                           n696, S0 => n697);
   U502 : HS65_LH_FA1X4 port map( A0 => n1231, B0 => n701, CI => n716, CO => 
                           n698, S0 => n699);
   U503 : HS65_LH_FA1X4 port map( A0 => n1199, B0 => n703, CI => n718, CO => 
                           n700, S0 => n701);
   U504 : HS65_LH_FA1X4 port map( A0 => n1167, B0 => n705, CI => n720, CO => 
                           n702, S0 => n703);
   U505 : HS65_LH_FA1X4 port map( A0 => n1135, B0 => n707, CI => n722, CO => 
                           n704, S0 => n705);
   U506 : HS65_LH_HA1X4 port map( A0 => n1103, B0 => n724, CO => n706, S0 => 
                           n707);
   U507 : HS65_LH_FA1X4 port map( A0 => n1360, B0 => n711, CI => n726, CO => 
                           n708, S0 => n709);
   U508 : HS65_LH_FA1X4 port map( A0 => n1328, B0 => n713, CI => n728, CO => 
                           n710, S0 => n711);
   U509 : HS65_LH_FA1X4 port map( A0 => n1296, B0 => n715, CI => n730, CO => 
                           n712, S0 => n713);
   U510 : HS65_LH_FA1X4 port map( A0 => n1264, B0 => n717, CI => n732, CO => 
                           n714, S0 => n715);
   U511 : HS65_LH_FA1X4 port map( A0 => n1232, B0 => n719, CI => n734, CO => 
                           n716, S0 => n717);
   U512 : HS65_LH_FA1X4 port map( A0 => n1200, B0 => n721, CI => n736, CO => 
                           n718, S0 => n719);
   U513 : HS65_LH_FA1X4 port map( A0 => n1168, B0 => n723, CI => n738, CO => 
                           n720, S0 => n721);
   U514 : HS65_LH_FA1X4 port map( A0 => n1136, B0 => n725, CI => n740, CO => 
                           n722, S0 => n723);
   U515 : HS65_LH_HA1X4 port map( A0 => n2656, B0 => n1104, CO => n724, S0 => 
                           n725);
   U516 : HS65_LH_FA1X4 port map( A0 => n1361, B0 => n729, CI => n742, CO => 
                           n726, S0 => n727);
   U517 : HS65_LH_FA1X4 port map( A0 => n1329, B0 => n731, CI => n744, CO => 
                           n728, S0 => n729);
   U518 : HS65_LH_FA1X4 port map( A0 => n1297, B0 => n733, CI => n746, CO => 
                           n730, S0 => n731);
   U519 : HS65_LH_FA1X4 port map( A0 => n1265, B0 => n735, CI => n748, CO => 
                           n732, S0 => n733);
   U520 : HS65_LH_FA1X4 port map( A0 => n1233, B0 => n737, CI => n750, CO => 
                           n734, S0 => n735);
   U521 : HS65_LH_FA1X4 port map( A0 => n1201, B0 => n739, CI => n752, CO => 
                           n736, S0 => n737);
   U522 : HS65_LH_FA1X4 port map( A0 => n1169, B0 => n741, CI => n754, CO => 
                           n738, S0 => n739);
   U523 : HS65_LH_HA1X4 port map( A0 => n1137, B0 => n756, CO => n740, S0 => 
                           n741);
   U524 : HS65_LH_FA1X4 port map( A0 => n1362, B0 => n745, CI => n758, CO => 
                           n742, S0 => n743);
   U525 : HS65_LH_FA1X4 port map( A0 => n1330, B0 => n747, CI => n760, CO => 
                           n744, S0 => n745);
   U526 : HS65_LH_FA1X4 port map( A0 => n1298, B0 => n749, CI => n762, CO => 
                           n746, S0 => n747);
   U527 : HS65_LH_FA1X4 port map( A0 => n1266, B0 => n751, CI => n764, CO => 
                           n748, S0 => n749);
   U528 : HS65_LH_FA1X4 port map( A0 => n1234, B0 => n753, CI => n766, CO => 
                           n750, S0 => n751);
   U529 : HS65_LH_FA1X4 port map( A0 => n1202, B0 => n755, CI => n768, CO => 
                           n752, S0 => n753);
   U530 : HS65_LH_FA1X4 port map( A0 => n1170, B0 => n757, CI => n770, CO => 
                           n754, S0 => n755);
   U531 : HS65_LH_HA1X4 port map( A0 => n1138, B0 => n772, CO => n756, S0 => 
                           n757);
   U532 : HS65_LH_FA1X4 port map( A0 => n1363, B0 => n761, CI => n774, CO => 
                           n758, S0 => n759);
   U533 : HS65_LH_FA1X4 port map( A0 => n1331, B0 => n763, CI => n776, CO => 
                           n760, S0 => n761);
   U534 : HS65_LH_FA1X4 port map( A0 => n1299, B0 => n765, CI => n778, CO => 
                           n762, S0 => n763);
   U535 : HS65_LH_FA1X4 port map( A0 => n1267, B0 => n767, CI => n780, CO => 
                           n764, S0 => n765);
   U536 : HS65_LH_FA1X4 port map( A0 => n1235, B0 => n769, CI => n782, CO => 
                           n766, S0 => n767);
   U537 : HS65_LH_FA1X4 port map( A0 => n1203, B0 => n771, CI => n784, CO => 
                           n768, S0 => n769);
   U538 : HS65_LH_FA1X4 port map( A0 => n1171, B0 => n773, CI => n786, CO => 
                           n770, S0 => n771);
   U539 : HS65_LH_HA1X4 port map( A0 => n2653, B0 => n1139, CO => n772, S0 => 
                           n773);
   U540 : HS65_LH_FA1X4 port map( A0 => n1364, B0 => n777, CI => n788, CO => 
                           n774, S0 => n775);
   U541 : HS65_LH_FA1X4 port map( A0 => n1332, B0 => n779, CI => n790, CO => 
                           n776, S0 => n777);
   U542 : HS65_LH_FA1X4 port map( A0 => n1300, B0 => n781, CI => n792, CO => 
                           n778, S0 => n779);
   U543 : HS65_LH_FA1X4 port map( A0 => n1268, B0 => n783, CI => n794, CO => 
                           n780, S0 => n781);
   U544 : HS65_LH_FA1X4 port map( A0 => n1236, B0 => n785, CI => n796, CO => 
                           n782, S0 => n783);
   U545 : HS65_LH_FA1X4 port map( A0 => n1204, B0 => n787, CI => n798, CO => 
                           n784, S0 => n785);
   U546 : HS65_LH_HA1X4 port map( A0 => n1172, B0 => n800, CO => n786, S0 => 
                           n787);
   U547 : HS65_LH_FA1X4 port map( A0 => n1365, B0 => n791, CI => n802, CO => 
                           n788, S0 => n789);
   U548 : HS65_LH_FA1X4 port map( A0 => n1333, B0 => n793, CI => n804, CO => 
                           n790, S0 => n791);
   U549 : HS65_LH_FA1X4 port map( A0 => n1301, B0 => n795, CI => n806, CO => 
                           n792, S0 => n793);
   U550 : HS65_LH_FA1X4 port map( A0 => n1269, B0 => n797, CI => n808, CO => 
                           n794, S0 => n795);
   U551 : HS65_LH_FA1X4 port map( A0 => n1237, B0 => n799, CI => n810, CO => 
                           n796, S0 => n797);
   U552 : HS65_LH_FA1X4 port map( A0 => n1205, B0 => n801, CI => n812, CO => 
                           n798, S0 => n799);
   U553 : HS65_LH_HA1X4 port map( A0 => n1173, B0 => n814, CO => n800, S0 => 
                           n801);
   U554 : HS65_LH_FA1X4 port map( A0 => n1366, B0 => n805, CI => n816, CO => 
                           n802, S0 => n803);
   U555 : HS65_LH_FA1X4 port map( A0 => n1334, B0 => n807, CI => n818, CO => 
                           n804, S0 => n805);
   U556 : HS65_LH_FA1X4 port map( A0 => n1302, B0 => n809, CI => n820, CO => 
                           n806, S0 => n807);
   U557 : HS65_LH_FA1X4 port map( A0 => n1270, B0 => n811, CI => n822, CO => 
                           n808, S0 => n809);
   U558 : HS65_LH_FA1X4 port map( A0 => n1238, B0 => n813, CI => n824, CO => 
                           n810, S0 => n811);
   U559 : HS65_LH_FA1X4 port map( A0 => n1206, B0 => n815, CI => n826, CO => 
                           n812, S0 => n813);
   U560 : HS65_LH_HA1X4 port map( A0 => n2650, B0 => n1174, CO => n814, S0 => 
                           n815);
   U561 : HS65_LH_FA1X4 port map( A0 => n1367, B0 => n819, CI => n828, CO => 
                           n816, S0 => n817);
   U562 : HS65_LH_FA1X4 port map( A0 => n1335, B0 => n821, CI => n830, CO => 
                           n818, S0 => n819);
   U563 : HS65_LH_FA1X4 port map( A0 => n1303, B0 => n823, CI => n832, CO => 
                           n820, S0 => n821);
   U564 : HS65_LH_FA1X4 port map( A0 => n1271, B0 => n825, CI => n834, CO => 
                           n822, S0 => n823);
   U565 : HS65_LH_FA1X4 port map( A0 => n1239, B0 => n827, CI => n836, CO => 
                           n824, S0 => n825);
   U566 : HS65_LH_HA1X4 port map( A0 => n1207, B0 => n838, CO => n826, S0 => 
                           n827);
   U567 : HS65_LH_FA1X4 port map( A0 => n1368, B0 => n831, CI => n840, CO => 
                           n828, S0 => n829);
   U568 : HS65_LH_FA1X4 port map( A0 => n1336, B0 => n833, CI => n842, CO => 
                           n830, S0 => n831);
   U569 : HS65_LH_FA1X4 port map( A0 => n1304, B0 => n835, CI => n844, CO => 
                           n832, S0 => n833);
   U570 : HS65_LH_FA1X4 port map( A0 => n1272, B0 => n837, CI => n846, CO => 
                           n834, S0 => n835);
   U571 : HS65_LH_FA1X4 port map( A0 => n1240, B0 => n839, CI => n848, CO => 
                           n836, S0 => n837);
   U572 : HS65_LH_HA1X4 port map( A0 => n1208, B0 => n850, CO => n838, S0 => 
                           n839);
   U573 : HS65_LH_FA1X4 port map( A0 => n1369, B0 => n843, CI => n852, CO => 
                           n840, S0 => n841);
   U574 : HS65_LH_FA1X4 port map( A0 => n1337, B0 => n845, CI => n854, CO => 
                           n842, S0 => n843);
   U575 : HS65_LH_FA1X4 port map( A0 => n1305, B0 => n847, CI => n856, CO => 
                           n844, S0 => n845);
   U576 : HS65_LH_FA1X4 port map( A0 => n1273, B0 => n849, CI => n858, CO => 
                           n846, S0 => n847);
   U577 : HS65_LH_FA1X4 port map( A0 => n1241, B0 => n851, CI => n860, CO => 
                           n848, S0 => n849);
   U578 : HS65_LH_HA1X4 port map( A0 => n2647, B0 => n1209, CO => n850, S0 => 
                           n851);
   U579 : HS65_LH_FA1X4 port map( A0 => n1370, B0 => n855, CI => n862, CO => 
                           n852, S0 => n853);
   U580 : HS65_LH_FA1X4 port map( A0 => n1338, B0 => n857, CI => n864, CO => 
                           n854, S0 => n855);
   U581 : HS65_LH_FA1X4 port map( A0 => n1306, B0 => n859, CI => n866, CO => 
                           n856, S0 => n857);
   U582 : HS65_LH_FA1X4 port map( A0 => n1274, B0 => n861, CI => n868, CO => 
                           n858, S0 => n859);
   U583 : HS65_LH_HA1X4 port map( A0 => n1242, B0 => n870, CO => n860, S0 => 
                           n861);
   U584 : HS65_LH_FA1X4 port map( A0 => n1371, B0 => n865, CI => n872, CO => 
                           n862, S0 => n863);
   U585 : HS65_LH_FA1X4 port map( A0 => n1339, B0 => n867, CI => n874, CO => 
                           n864, S0 => n865);
   U586 : HS65_LH_FA1X4 port map( A0 => n1307, B0 => n869, CI => n876, CO => 
                           n866, S0 => n867);
   U587 : HS65_LH_FA1X4 port map( A0 => n1275, B0 => n871, CI => n878, CO => 
                           n868, S0 => n869);
   U588 : HS65_LH_HA1X4 port map( A0 => n1243, B0 => n880, CO => n870, S0 => 
                           n871);
   U589 : HS65_LH_FA1X4 port map( A0 => n1372, B0 => n875, CI => n882, CO => 
                           n872, S0 => n873);
   U590 : HS65_LH_FA1X4 port map( A0 => n1340, B0 => n877, CI => n884, CO => 
                           n874, S0 => n875);
   U591 : HS65_LH_FA1X4 port map( A0 => n1308, B0 => n879, CI => n886, CO => 
                           n876, S0 => n877);
   U592 : HS65_LH_FA1X4 port map( A0 => n1276, B0 => n881, CI => n888, CO => 
                           n878, S0 => n879);
   U593 : HS65_LH_HA1X4 port map( A0 => n2644, B0 => n1244, CO => n880, S0 => 
                           n881);
   U594 : HS65_LH_FA1X4 port map( A0 => n1373, B0 => n885, CI => n890, CO => 
                           n882, S0 => n883);
   U595 : HS65_LH_FA1X4 port map( A0 => n1341, B0 => n887, CI => n892, CO => 
                           n884, S0 => n885);
   U596 : HS65_LH_FA1X4 port map( A0 => n1309, B0 => n889, CI => n894, CO => 
                           n886, S0 => n887);
   U597 : HS65_LH_HA1X4 port map( A0 => n1277, B0 => n896, CO => n888, S0 => 
                           n889);
   U598 : HS65_LH_FA1X4 port map( A0 => n1374, B0 => n893, CI => n898, CO => 
                           n890, S0 => n891);
   U599 : HS65_LH_FA1X4 port map( A0 => n1342, B0 => n895, CI => n900, CO => 
                           n892, S0 => n893);
   U600 : HS65_LH_FA1X4 port map( A0 => n1310, B0 => n897, CI => n902, CO => 
                           n894, S0 => n895);
   U601 : HS65_LH_HA1X4 port map( A0 => n1278, B0 => n904, CO => n896, S0 => 
                           n897);
   U602 : HS65_LH_FA1X4 port map( A0 => n1375, B0 => n901, CI => n906, CO => 
                           n898, S0 => n899);
   U603 : HS65_LH_FA1X4 port map( A0 => n1343, B0 => n903, CI => n908, CO => 
                           n900, S0 => n901);
   U604 : HS65_LH_FA1X4 port map( A0 => n1311, B0 => n905, CI => n910, CO => 
                           n902, S0 => n903);
   U605 : HS65_LH_HA1X4 port map( A0 => n2641, B0 => n1279, CO => n904, S0 => 
                           n905);
   U606 : HS65_LH_FA1X4 port map( A0 => n1376, B0 => n909, CI => n912, CO => 
                           n906, S0 => n907);
   U607 : HS65_LH_FA1X4 port map( A0 => n1344, B0 => n911, CI => n914, CO => 
                           n908, S0 => n909);
   U608 : HS65_LH_HA1X4 port map( A0 => n1312, B0 => n916, CO => n910, S0 => 
                           n911);
   U609 : HS65_LH_FA1X4 port map( A0 => n1377, B0 => n915, CI => n918, CO => 
                           n912, S0 => n913);
   U610 : HS65_LH_FA1X4 port map( A0 => n1345, B0 => n917, CI => n920, CO => 
                           n914, S0 => n915);
   U611 : HS65_LH_HA1X4 port map( A0 => n1313, B0 => n922, CO => n916, S0 => 
                           n917);
   U612 : HS65_LH_FA1X4 port map( A0 => n1378, B0 => n921, CI => n924, CO => 
                           n918, S0 => n919);
   U613 : HS65_LH_FA1X4 port map( A0 => n1346, B0 => n923, CI => n926, CO => 
                           n920, S0 => n921);
   U614 : HS65_LH_HA1X4 port map( A0 => n2638, B0 => n1314, CO => n922, S0 => 
                           n923);
   U615 : HS65_LH_FA1X4 port map( A0 => n1379, B0 => n927, CI => n928, CO => 
                           n924, S0 => n925);
   U616 : HS65_LH_HA1X4 port map( A0 => n1347, B0 => n930, CO => n926, S0 => 
                           n927);
   U617 : HS65_LH_FA1X4 port map( A0 => n1380, B0 => n931, CI => n932, CO => 
                           n928, S0 => n929);
   U618 : HS65_LH_HA1X4 port map( A0 => n1348, B0 => n934, CO => n930, S0 => 
                           n931);
   U619 : HS65_LH_FA1X4 port map( A0 => n1381, B0 => n935, CI => n936, CO => 
                           n932, S0 => n933);
   U620 : HS65_LH_HA1X4 port map( A0 => n2635, B0 => n1349, CO => n934, S0 => 
                           n935);
   U621 : HS65_LH_HA1X4 port map( A0 => n1382, B0 => n938, CO => n936, S0 => 
                           n937);
   U622 : HS65_LH_HA1X4 port map( A0 => n1383, B0 => n940, CO => n938, S0 => 
                           n939);
   U623 : HS65_LH_HA1X4 port map( A0 => n2632, B0 => n1384, CO => n940, S0 => 
                           n941);
   U1907 : HS65_LH_HA1X4 port map( A0 => n2626, B0 => n975, CO => n1006, S0 => 
                           n1007);
   U1908 : HS65_LH_FA1X4 port map( A0 => n2624, B0 => n2626, CI => n976, CO => 
                           n975, S0 => n1008);
   U1909 : HS65_LH_FA1X4 port map( A0 => n2622, B0 => n2624, CI => n977, CO => 
                           n976, S0 => n1009);
   U1910 : HS65_LH_FA1X4 port map( A0 => n2620, B0 => n2622, CI => n978, CO => 
                           n977, S0 => n1010);
   U1911 : HS65_LH_FA1X4 port map( A0 => n2618, B0 => n2620, CI => n979, CO => 
                           n978, S0 => n1011);
   U1912 : HS65_LH_FA1X4 port map( A0 => n2616, B0 => n2618, CI => n980, CO => 
                           n979, S0 => n1012);
   U1913 : HS65_LH_FA1X4 port map( A0 => n2614, B0 => n2616, CI => n981, CO => 
                           n980, S0 => n1013);
   U1914 : HS65_LH_FA1X4 port map( A0 => n2612, B0 => n2614, CI => n982, CO => 
                           n981, S0 => n1014);
   U1915 : HS65_LH_FA1X4 port map( A0 => n2610, B0 => n2612, CI => n983, CO => 
                           n982, S0 => n1015);
   U1916 : HS65_LH_FA1X4 port map( A0 => n2608, B0 => n2610, CI => n984, CO => 
                           n983, S0 => n1016);
   U1917 : HS65_LH_FA1X4 port map( A0 => n2606, B0 => n2608, CI => n985, CO => 
                           n984, S0 => n1017);
   U1918 : HS65_LH_FA1X4 port map( A0 => n2604, B0 => n2606, CI => n986, CO => 
                           n985, S0 => n1018);
   U1919 : HS65_LH_FA1X4 port map( A0 => n2602, B0 => n2604, CI => n987, CO => 
                           n986, S0 => n1019);
   U1920 : HS65_LH_FA1X4 port map( A0 => n2600, B0 => n2602, CI => n988, CO => 
                           n987, S0 => n1020);
   U1921 : HS65_LH_FA1X4 port map( A0 => n2598, B0 => n2600, CI => n989, CO => 
                           n988, S0 => n1021);
   U1922 : HS65_LH_FA1X4 port map( A0 => n2596, B0 => n2598, CI => n990, CO => 
                           n989, S0 => n1022);
   U1923 : HS65_LH_FA1X4 port map( A0 => n2594, B0 => n2596, CI => n991, CO => 
                           n990, S0 => n1023);
   U1924 : HS65_LH_FA1X4 port map( A0 => n2592, B0 => n2594, CI => n992, CO => 
                           n991, S0 => n1024);
   U1925 : HS65_LH_FA1X4 port map( A0 => n2590, B0 => n2592, CI => n993, CO => 
                           n992, S0 => n1025);
   U1926 : HS65_LH_FA1X4 port map( A0 => n2588, B0 => n2590, CI => n994, CO => 
                           n993, S0 => n1026);
   U1927 : HS65_LH_FA1X4 port map( A0 => n2586, B0 => n2588, CI => n995, CO => 
                           n994, S0 => n1027);
   U1928 : HS65_LH_FA1X4 port map( A0 => n2584, B0 => n2586, CI => n996, CO => 
                           n995, S0 => n1028);
   U1929 : HS65_LH_FA1X4 port map( A0 => n2582, B0 => n2584, CI => n997, CO => 
                           n996, S0 => n1029);
   U1930 : HS65_LH_FA1X4 port map( A0 => n2580, B0 => n2582, CI => n998, CO => 
                           n997, S0 => n1030);
   U1931 : HS65_LH_FA1X4 port map( A0 => n2578, B0 => n2580, CI => n999, CO => 
                           n998, S0 => n1031);
   U1932 : HS65_LH_FA1X4 port map( A0 => n2576, B0 => n2578, CI => n1000, CO =>
                           n999, S0 => n1032);
   U1933 : HS65_LH_FA1X4 port map( A0 => n2574, B0 => n2576, CI => n1001, CO =>
                           n1000, S0 => n1033);
   U1934 : HS65_LH_FA1X4 port map( A0 => n2572, B0 => n2574, CI => n1002, CO =>
                           n1001, S0 => n1034);
   U1935 : HS65_LH_FA1X4 port map( A0 => n2570, B0 => n2572, CI => n1003, CO =>
                           n1002, S0 => n1035);
   U1936 : HS65_LH_FA1X4 port map( A0 => n2568, B0 => n2570, CI => n1004, CO =>
                           n1003, S0 => n1036);
   U1937 : HS65_LH_FA1X4 port map( A0 => n2566, B0 => n2568, CI => n1005, CO =>
                           n1004, S0 => n1037);
   U1941 : HS65_LH_IVX9 port map( A => a(2), Z => n2630);
   U1942 : HS65_LH_IVX9 port map( A => n1007, Z => n2667);
   U1943 : HS65_LH_IVX9 port map( A => n2630, Z => n2628);
   U1944 : HS65_LH_IVX9 port map( A => n2630, Z => n2629);
   U1945 : HS65_LH_BFX9 port map( A => n2668, Z => n2422);
   U1946 : HS65_LH_BFX9 port map( A => n2445, Z => n2446);
   U1947 : HS65_LH_BFX9 port map( A => n2457, Z => n2454);
   U1948 : HS65_LH_BFX9 port map( A => n2457, Z => n2455);
   U1949 : HS65_LH_BFX9 port map( A => n2453, Z => n2450);
   U1950 : HS65_LH_BFX9 port map( A => n2466, Z => n2463);
   U1951 : HS65_LH_IVX9 port map( A => n2636, Z => n2635);
   U1952 : HS65_LH_IVX9 port map( A => n2633, Z => n2632);
   U1953 : HS65_LH_IVX9 port map( A => n2449, Z => n2448);
   U1954 : HS65_LH_BFX9 port map( A => n2668, Z => n2421);
   U1955 : HS65_LH_BFX9 port map( A => n2458, Z => n2459);
   U1956 : HS65_LH_BFX9 port map( A => n2484, Z => n2485);
   U1957 : HS65_LH_BFX9 port map( A => n2497, Z => n2498);
   U1958 : HS65_LH_BFX9 port map( A => n2510, Z => n2511);
   U1959 : HS65_LH_BFX9 port map( A => n2471, Z => n2472);
   U1960 : HS65_LH_BFX9 port map( A => n2453, Z => n2451);
   U1961 : HS65_LH_BFX9 port map( A => n2479, Z => n2477);
   U1962 : HS65_LH_BFX9 port map( A => n2470, Z => n2467);
   U1963 : HS65_LH_BFX9 port map( A => n2496, Z => n2493);
   U1964 : HS65_LH_BFX9 port map( A => n2509, Z => n2506);
   U1965 : HS65_LH_BFX9 port map( A => n2522, Z => n2519);
   U1966 : HS65_LH_BFX9 port map( A => n2470, Z => n2468);
   U1967 : HS65_LH_BFX9 port map( A => n2496, Z => n2494);
   U1968 : HS65_LH_BFX9 port map( A => n2509, Z => n2507);
   U1969 : HS65_LH_BFX9 port map( A => n2522, Z => n2520);
   U1970 : HS65_LH_BFX9 port map( A => n2483, Z => n2480);
   U1971 : HS65_LH_BFX9 port map( A => n2479, Z => n2476);
   U1972 : HS65_LH_BFX9 port map( A => n2492, Z => n2489);
   U1973 : HS65_LH_BFX9 port map( A => n2505, Z => n2502);
   U1974 : HS65_LH_BFX9 port map( A => n2518, Z => n2515);
   U1975 : HS65_LH_BFX9 port map( A => n2483, Z => n2481);
   U1976 : HS65_LH_IVX9 port map( A => n2642, Z => n2641);
   U1977 : HS65_LH_IVX9 port map( A => n2639, Z => n2638);
   U1978 : HS65_LH_IVX9 port map( A => n2648, Z => n2647);
   U1979 : HS65_LH_IVX9 port map( A => n2645, Z => n2644);
   U1980 : HS65_LH_IVX9 port map( A => n2462, Z => n2461);
   U1981 : HS65_LH_IVX9 port map( A => n2475, Z => n2474);
   U1982 : HS65_LH_IVX9 port map( A => n2488, Z => n2487);
   U1983 : HS65_LH_IVX9 port map( A => n2501, Z => n2500);
   U1984 : HS65_LH_IVX9 port map( A => n2514, Z => n2513);
   U1985 : HS65_LH_BFX9 port map( A => n2536, Z => n2537);
   U1986 : HS65_LH_BFX9 port map( A => n2549, Z => n2550);
   U1987 : HS65_LH_BFX9 port map( A => n2523, Z => n2524);
   U1988 : HS65_LH_BFX9 port map( A => n2535, Z => n2533);
   U1989 : HS65_LH_BFX9 port map( A => n2466, Z => n2464);
   U1990 : HS65_LH_BFX9 port map( A => n2492, Z => n2490);
   U1991 : HS65_LH_BFX9 port map( A => n2505, Z => n2503);
   U1992 : HS65_LH_BFX9 port map( A => n2518, Z => n2516);
   U1993 : HS65_LH_BFX9 port map( A => n2561, Z => n2558);
   U1994 : HS65_LH_BFX9 port map( A => n2548, Z => n2545);
   U1995 : HS65_LH_BFX9 port map( A => n2548, Z => n2546);
   U1996 : HS65_LH_BFX9 port map( A => n2561, Z => n2559);
   U1997 : HS65_LH_BFX9 port map( A => n2535, Z => n2532);
   U1998 : HS65_LH_BFX9 port map( A => n2531, Z => n2528);
   U1999 : HS65_LH_BFX9 port map( A => n2544, Z => n2541);
   U2000 : HS65_LH_BFX9 port map( A => n2557, Z => n2554);
   U2001 : HS65_LH_IVX9 port map( A => n2654, Z => n2653);
   U2002 : HS65_LH_IVX9 port map( A => n2657, Z => n2656);
   U2003 : HS65_LH_IVX9 port map( A => n2651, Z => n2650);
   U2004 : HS65_LH_IVX9 port map( A => n2527, Z => n2526);
   U2005 : HS65_LH_IVX9 port map( A => n2540, Z => n2539);
   U2006 : HS65_LH_IVX9 port map( A => n2553, Z => n2552);
   U2007 : HS65_LH_IVX9 port map( A => n510, Z => n2662);
   U2008 : HS65_LH_IVX9 port map( A => n462, Z => n2661);
   U2009 : HS65_LH_BFX9 port map( A => n2666, Z => n2418);
   U2010 : HS65_LH_BFX9 port map( A => n2668, Z => n2420);
   U2011 : HS65_LH_BFX9 port map( A => n2666, Z => n2419);
   U2012 : HS65_LH_BFX9 port map( A => n2433, Z => n2430);
   U2013 : HS65_LH_BFX9 port map( A => n2471, Z => n2473);
   U2014 : HS65_LH_BFX9 port map( A => n2531, Z => n2529);
   U2015 : HS65_LH_BFX9 port map( A => n2544, Z => n2542);
   U2016 : HS65_LH_BFX9 port map( A => n2557, Z => n2555);
   U2017 : HS65_LH_BFX9 port map( A => n2445, Z => n2447);
   U2018 : HS65_LH_BFX9 port map( A => n2458, Z => n2460);
   U2019 : HS65_LH_BFX9 port map( A => n2484, Z => n2486);
   U2020 : HS65_LH_BFX9 port map( A => n2433, Z => n2432);
   U2021 : HS65_LH_IVX9 port map( A => n419, Z => n2665);
   U2022 : HS65_LH_IVX9 port map( A => n352, Z => n2664);
   U2023 : HS65_LH_IVX9 port map( A => n383, Z => n2660);
   U2024 : HS65_LH_IVX9 port map( A => n328, Z => n2659);
   U2025 : HS65_LH_BFX9 port map( A => n2523, Z => n2525);
   U2026 : HS65_LH_BFX9 port map( A => n2497, Z => n2499);
   U2027 : HS65_LH_BFX9 port map( A => n2510, Z => n2512);
   U2028 : HS65_LH_BFX9 port map( A => n2457, Z => n2456);
   U2029 : HS65_LH_BFX9 port map( A => n2470, Z => n2469);
   U2030 : HS65_LH_BFX9 port map( A => n2453, Z => n2452);
   U2031 : HS65_LH_BFX9 port map( A => n2466, Z => n2465);
   U2032 : HS65_LH_BFX9 port map( A => n2479, Z => n2478);
   U2033 : HS65_LH_IVX9 port map( A => n309, Z => n2663);
   U2034 : HS65_LH_IVX9 port map( A => n297, Z => n2658);
   U2035 : HS65_LH_BFX9 port map( A => n2433, Z => n2431);
   U2036 : HS65_LH_BFX9 port map( A => n2536, Z => n2538);
   U2037 : HS65_LH_BFX9 port map( A => n2549, Z => n2551);
   U2038 : HS65_LH_BFX9 port map( A => n2496, Z => n2495);
   U2039 : HS65_LH_BFX9 port map( A => n2509, Z => n2508);
   U2040 : HS65_LH_BFX9 port map( A => n2483, Z => n2482);
   U2041 : HS65_LH_BFX9 port map( A => n2492, Z => n2491);
   U2042 : HS65_LH_BFX9 port map( A => n2505, Z => n2504);
   U2043 : HS65_LH_BFX9 port map( A => n2666, Z => n2417);
   U2044 : HS65_LH_BFX9 port map( A => n2522, Z => n2521);
   U2045 : HS65_LH_BFX9 port map( A => n2531, Z => n2530);
   U2046 : HS65_LH_BFX9 port map( A => n2518, Z => n2517);
   U2047 : HS65_LH_BFX9 port map( A => n2548, Z => n2547);
   U2048 : HS65_LH_BFX9 port map( A => n2561, Z => n2560);
   U2049 : HS65_LH_BFX9 port map( A => n2535, Z => n2534);
   U2050 : HS65_LH_BFX9 port map( A => n2544, Z => n2543);
   U2051 : HS65_LH_BFX9 port map( A => n2557, Z => n2556);
   U2052 : HS65_LH_IVX9 port map( A => n2713, Z => n2668);
   U2053 : HS65_LH_BFX9 port map( A => n2723, Z => n2457);
   U2054 : HS65_LH_BFX9 port map( A => n2721, Z => n2453);
   U2055 : HS65_LH_BFX9 port map( A => n2764, Z => n2466);
   U2056 : HS65_LH_IVX9 port map( A => a(5), Z => n2633);
   U2057 : HS65_LH_IVX9 port map( A => n2719, Z => n2449);
   U2058 : HS65_LH_IVX9 port map( A => n2762, Z => n2462);
   U2059 : HS65_LH_HA1X4 port map( A0 => n2566, B0 => n2563, CO => n1005, S0 =>
                           n1038);
   U2060 : HS65_LH_BFX9 port map( A => n2718, Z => n2445);
   U2061 : HS65_LH_BFX9 port map( A => b(2), Z => n2568);
   U2062 : HS65_LH_BFX9 port map( A => n2562, Z => n2563);
   U2063 : HS65_LH_BFX9 port map( A => n2436, Z => n2434);
   U2064 : HS65_LH_BFX9 port map( A => n2444, Z => n2441);
   U2065 : HS65_LH_BFX9 port map( A => n2444, Z => n2442);
   U2066 : HS65_LH_IVX9 port map( A => n2633, Z => n2631);
   U2067 : HS65_LH_BFX9 port map( A => n2444, Z => n2443);
   U2068 : HS65_LH_BFX9 port map( A => n2766, Z => n2470);
   U2069 : HS65_LH_BFX9 port map( A => n2809, Z => n2483);
   U2070 : HS65_LH_IVX9 port map( A => n2891, Z => n2501);
   U2071 : HS65_LH_IVX9 port map( A => n2934, Z => n2514);
   U2072 : HS65_LH_BFX9 port map( A => n2852, Z => n2496);
   U2073 : HS65_LH_BFX9 port map( A => n2895, Z => n2509);
   U2074 : HS65_LH_BFX9 port map( A => n2938, Z => n2522);
   U2075 : HS65_LH_BFX9 port map( A => n2850, Z => n2492);
   U2076 : HS65_LH_BFX9 port map( A => n2893, Z => n2505);
   U2077 : HS65_LH_BFX9 port map( A => n2936, Z => n2518);
   U2078 : HS65_LH_BFX9 port map( A => n2807, Z => n2479);
   U2079 : HS65_LH_IVX9 port map( A => a(14), Z => n2642);
   U2080 : HS65_LH_IVX9 port map( A => a(11), Z => n2639);
   U2081 : HS65_LH_IVX9 port map( A => a(20), Z => n2648);
   U2082 : HS65_LH_IVX9 port map( A => a(17), Z => n2645);
   U2083 : HS65_LH_IVX9 port map( A => n2848, Z => n2488);
   U2084 : HS65_LH_IVX9 port map( A => n2977, Z => n2527);
   U2085 : HS65_LH_IVX9 port map( A => n2805, Z => n2475);
   U2086 : HS65_LH_BFX9 port map( A => n2761, Z => n2458);
   U2087 : HS65_LH_BFX9 port map( A => n2804, Z => n2471);
   U2088 : HS65_LH_BFX9 port map( A => n2847, Z => n2484);
   U2089 : HS65_LH_BFX9 port map( A => n2890, Z => n2497);
   U2090 : HS65_LH_BFX9 port map( A => n2933, Z => n2510);
   U2091 : HS65_LH_BFX9 port map( A => b(3), Z => n2570);
   U2092 : HS65_LH_BFX9 port map( A => b(4), Z => n2572);
   U2093 : HS65_LH_BFX9 port map( A => n2562, Z => n2564);
   U2094 : HS65_LH_BFX9 port map( A => b(2), Z => n2569);
   U2095 : HS65_LH_BFX9 port map( A => b(3), Z => n2571);
   U2096 : HS65_LH_BFX9 port map( A => n2440, Z => n2437);
   U2097 : HS65_LH_BFX9 port map( A => b(4), Z => n2573);
   U2098 : HS65_LH_IVX9 port map( A => n2636, Z => n2634);
   U2099 : HS65_LH_IVX9 port map( A => a(8), Z => n2636);
   U2100 : HS65_LH_IVX9 port map( A => n2642, Z => n2640);
   U2101 : HS65_LH_IVX9 port map( A => n2639, Z => n2637);
   U2102 : HS65_LH_IVX9 port map( A => n2648, Z => n2646);
   U2103 : HS65_LH_IVX9 port map( A => n2645, Z => n2643);
   U2104 : HS65_LH_BFX9 port map( A => n2562, Z => n2565);
   U2105 : HS65_LH_BFX9 port map( A => n2440, Z => n2439);
   U2106 : HS65_LH_BFX9 port map( A => n3067, Z => n2561);
   U2107 : HS65_LH_BFX9 port map( A => n3022, Z => n2544);
   U2108 : HS65_LH_BFX9 port map( A => n2981, Z => n2535);
   U2109 : HS65_LH_BFX9 port map( A => n3024, Z => n2548);
   U2110 : HS65_LH_BFX9 port map( A => n2979, Z => n2531);
   U2111 : HS65_LH_BFX9 port map( A => n3065, Z => n2557);
   U2112 : HS65_LH_IVX9 port map( A => a(29), Z => n2657);
   U2113 : HS65_LH_IVX9 port map( A => n3020, Z => n2540);
   U2114 : HS65_LH_IVX9 port map( A => n3063, Z => n2553);
   U2115 : HS65_LH_BFX9 port map( A => n2976, Z => n2523);
   U2116 : HS65_LH_BFX9 port map( A => n3019, Z => n2536);
   U2117 : HS65_LH_BFX9 port map( A => n3062, Z => n2549);
   U2118 : HS65_LH_IVX9 port map( A => n2654, Z => n2652);
   U2119 : HS65_LH_IVX9 port map( A => a(26), Z => n2654);
   U2120 : HS65_LH_IVX9 port map( A => n2651, Z => n2649);
   U2121 : HS65_LH_IVX9 port map( A => a(23), Z => n2651);
   U2122 : HS65_LH_BFX9 port map( A => b(11), Z => n2586);
   U2123 : HS65_LH_BFX9 port map( A => b(11), Z => n2587);
   U2124 : HS65_LH_BFX9 port map( A => n2440, Z => n2438);
   U2125 : HS65_LH_BFX9 port map( A => n2436, Z => n2435);
   U2126 : HS65_LH_IVX9 port map( A => n2657, Z => n2655);
   U2127 : HS65_LH_BFX9 port map( A => n2429, Z => n2428);
   U2128 : HS65_LH_BFX9 port map( A => n2672, Z => n2433);
   U2129 : HS65_LH_IVX9 port map( A => n2673, Z => n2666);
   U2130 : HS65_LH_BFX9 port map( A => b(20), Z => n2604);
   U2131 : HS65_LH_BFX9 port map( A => n2425, Z => n2423);
   U2132 : HS65_LH_BFX9 port map( A => n2429, Z => n2426);
   U2133 : HS65_LH_BFX9 port map( A => b(27), Z => n2618);
   U2134 : HS65_LH_BFX9 port map( A => b(28), Z => n2620);
   U2135 : HS65_LH_BFX9 port map( A => n2425, Z => n2424);
   U2136 : HS65_LH_BFX9 port map( A => b(20), Z => n2605);
   U2137 : HS65_LH_BFX9 port map( A => b(31), Z => n2626);
   U2138 : HS65_LH_BFX9 port map( A => b(27), Z => n2619);
   U2139 : HS65_LH_BFX9 port map( A => b(28), Z => n2621);
   U2140 : HS65_LH_BFX9 port map( A => b(31), Z => n2627);
   U2141 : HS65_LH_BFX9 port map( A => n2429, Z => n2427);
   U2142 : HS65_LH_BFX9 port map( A => n2681, Z => n2444);
   U2143 : HS65_LH_BFX9 port map( A => n2677, Z => n2436);
   U2144 : HS65_LH_BFX9 port map( A => b(0), Z => n2562);
   U2145 : HS65_LH_BFX9 port map( A => n2679, Z => n2440);
   U2146 : HS65_LH_BFX9 port map( A => b(1), Z => n2566);
   U2147 : HS65_LH_BFX9 port map( A => b(5), Z => n2574);
   U2148 : HS65_LH_BFX9 port map( A => b(7), Z => n2578);
   U2149 : HS65_LH_BFX9 port map( A => b(6), Z => n2576);
   U2150 : HS65_LH_BFX9 port map( A => b(8), Z => n2580);
   U2151 : HS65_LH_BFX9 port map( A => b(5), Z => n2575);
   U2152 : HS65_LH_BFX9 port map( A => b(1), Z => n2567);
   U2153 : HS65_LH_BFX9 port map( A => b(6), Z => n2577);
   U2154 : HS65_LH_BFX9 port map( A => n2671, Z => n2429);
   U2155 : HS65_LH_BFX9 port map( A => b(12), Z => n2588);
   U2156 : HS65_LH_BFX9 port map( A => b(13), Z => n2590);
   U2157 : HS65_LH_BFX9 port map( A => b(9), Z => n2582);
   U2158 : HS65_LH_BFX9 port map( A => b(14), Z => n2592);
   U2159 : HS65_LH_BFX9 port map( A => b(10), Z => n2584);
   U2160 : HS65_LH_BFX9 port map( A => b(12), Z => n2589);
   U2161 : HS65_LH_BFX9 port map( A => b(7), Z => n2579);
   U2162 : HS65_LH_BFX9 port map( A => b(9), Z => n2583);
   U2163 : HS65_LH_BFX9 port map( A => b(8), Z => n2581);
   U2164 : HS65_LH_BFX9 port map( A => b(10), Z => n2585);
   U2165 : HS65_LH_BFX9 port map( A => n2670, Z => n2425);
   U2166 : HS65_LH_BFX9 port map( A => b(19), Z => n2602);
   U2167 : HS65_LH_BFX9 port map( A => b(18), Z => n2600);
   U2168 : HS65_LH_BFX9 port map( A => b(15), Z => n2594);
   U2169 : HS65_LH_BFX9 port map( A => b(17), Z => n2598);
   U2170 : HS65_LH_BFX9 port map( A => b(21), Z => n2606);
   U2171 : HS65_LH_BFX9 port map( A => b(16), Z => n2596);
   U2172 : HS65_LH_BFX9 port map( A => b(19), Z => n2603);
   U2173 : HS65_LH_BFX9 port map( A => b(13), Z => n2591);
   U2174 : HS65_LH_BFX9 port map( A => b(18), Z => n2601);
   U2175 : HS65_LH_BFX9 port map( A => b(15), Z => n2595);
   U2176 : HS65_LH_BFX9 port map( A => b(17), Z => n2599);
   U2177 : HS65_LH_BFX9 port map( A => b(14), Z => n2593);
   U2178 : HS65_LH_BFX9 port map( A => b(16), Z => n2597);
   U2179 : HS65_LH_BFX9 port map( A => b(23), Z => n2610);
   U2180 : HS65_LH_BFX9 port map( A => b(25), Z => n2614);
   U2181 : HS65_LH_BFX9 port map( A => b(24), Z => n2612);
   U2182 : HS65_LH_BFX9 port map( A => b(26), Z => n2616);
   U2183 : HS65_LH_BFX9 port map( A => b(22), Z => n2608);
   U2184 : HS65_LH_BFX9 port map( A => b(23), Z => n2611);
   U2185 : HS65_LH_BFX9 port map( A => b(25), Z => n2615);
   U2186 : HS65_LH_BFX9 port map( A => b(24), Z => n2613);
   U2187 : HS65_LH_BFX9 port map( A => b(21), Z => n2607);
   U2188 : HS65_LH_BFX9 port map( A => b(22), Z => n2609);
   U2189 : HS65_LH_BFX9 port map( A => b(29), Z => n2622);
   U2190 : HS65_LH_BFX9 port map( A => b(30), Z => n2624);
   U2191 : HS65_LH_BFX9 port map( A => b(26), Z => n2617);
   U2192 : HS65_LH_BFX9 port map( A => b(29), Z => n2623);
   U2193 : HS65_LH_BFX9 port map( A => b(30), Z => n2625);
   U2194 : HS65_LHS_XOR3X2 port map( A => n292, B => n227, C => n2669, Z => 
                           product(63));
   U2195 : HS65_LH_AO22X4 port map( A => n2627, B => n2423, C => n2419, D => 
                           n1006, Z => n2669);
   U2196 : HS65_LH_MX41X4 port map( D0 => n1025, S0 => n2419, D1 => n2593, S1 
                           => n2427, D2 => n2591, S2 => n2431, D3 => n2589, S3 
                           => n2423, Z => n419);
   U2197 : HS65_LH_MX41X4 port map( D0 => n1019, S0 => n2419, D1 => n2601, S1 
                           => n2423, D2 => n2603, S2 => n2430, D3 => n2605, S3 
                           => n2426, Z => n352);
   U2198 : HS65_LH_MX41X4 port map( D0 => n1013, S0 => n2419, D1 => n2613, S1 
                           => n2423, D2 => n2615, S2 => n2430, D3 => n2617, S3 
                           => n2426, Z => n309);
   U2199 : HS65_LH_OA12X4 port map( A => n2673, B => n2667, C => n2674, Z => 
                           n292);
   U2200 : HS65_LH_OAI22X1 port map( A => n2625, B => n2675, C => n2423, D => 
                           n2675, Z => n2674);
   U2201 : HS65_LH_AND2X4 port map( A => n2626, B => n2430, Z => n2675);
   U2202 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2676, Z => n1419);
   U2203 : HS65_LH_AO22X4 port map( A => n2565, B => n2434, C => n2422, D => 
                           n2564, Z => n2676);
   U2204 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2678, Z => n1418);
   U2205 : HS65_LH_AO222X4 port map( A => n2564, B => n2437, C => n2434, D => 
                           n2566, E => n2422, F => n1038, Z => n2678);
   U2206 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2680, Z => n1417);
   U2207 : HS65_LH_MX41X4 port map( D0 => n1037, S0 => n2422, D1 => n2442, S1 
                           => n2564, D2 => n2439, S2 => n2566, D3 => n2569, S3 
                           => n2434, Z => n2680);
   U2208 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2682, Z => n1416);
   U2209 : HS65_LH_MX41X4 port map( D0 => n1036, S0 => n2421, D1 => n2443, S1 
                           => n2567, D2 => n2569, S2 => n2437, D3 => n2571, S3 
                           => n2434, Z => n2682);
   U2210 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2683, Z => n1415);
   U2211 : HS65_LH_MX41X4 port map( D0 => n1035, S0 => n2422, D1 => n2443, S1 
                           => n2569, D2 => n2571, S2 => n2437, D3 => n2573, S3 
                           => n2434, Z => n2683);
   U2212 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2684, Z => n1414);
   U2213 : HS65_LH_MX41X4 port map( D0 => n1034, S0 => n2422, D1 => n2571, S1 
                           => n2441, D2 => n2573, S2 => n2437, D3 => n2575, S3 
                           => n2434, Z => n2684);
   U2214 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2685, Z => n1413);
   U2215 : HS65_LH_MX41X4 port map( D0 => n1033, S0 => n2421, D1 => n2573, S1 
                           => n2441, D2 => n2575, S2 => n2437, D3 => n2577, S3 
                           => n2434, Z => n2685);
   U2216 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2686, Z => n1412);
   U2217 : HS65_LH_MX41X4 port map( D0 => n1032, S0 => n2421, D1 => n2575, S1 
                           => n2441, D2 => n2577, S2 => n2437, D3 => n2579, S3 
                           => n2434, Z => n2686);
   U2218 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2687, Z => n1411);
   U2219 : HS65_LH_MX41X4 port map( D0 => n1031, S0 => n2421, D1 => n2577, S1 
                           => n2441, D2 => n2579, S2 => n2437, D3 => n2581, S3 
                           => n2434, Z => n2687);
   U2220 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2688, Z => n1410);
   U2221 : HS65_LH_MX41X4 port map( D0 => n1030, S0 => n2421, D1 => n2579, S1 
                           => n2441, D2 => n2581, S2 => n2437, D3 => n2583, S3 
                           => n2434, Z => n2688);
   U2222 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2689, Z => n1409);
   U2223 : HS65_LH_MX41X4 port map( D0 => n1029, S0 => n2421, D1 => n2581, S1 
                           => n2441, D2 => n2583, S2 => n2437, D3 => n2585, S3 
                           => n2434, Z => n2689);
   U2224 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2690, Z => n1408);
   U2225 : HS65_LH_MX41X4 port map( D0 => n1028, S0 => n2421, D1 => n2583, S1 
                           => n2441, D2 => n2585, S2 => n2437, D3 => n2587, S3 
                           => n2434, Z => n2690);
   U2226 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2691, Z => n1407);
   U2227 : HS65_LH_MX41X4 port map( D0 => n1027, S0 => n2421, D1 => n2585, S1 
                           => n2441, D2 => n2587, S2 => n2437, D3 => n2435, S3 
                           => n2589, Z => n2691);
   U2228 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2692, Z => n1406);
   U2229 : HS65_LH_MX41X4 port map( D0 => n1026, S0 => n2421, D1 => n2587, S1 
                           => n2441, D2 => n2438, S2 => n2588, D3 => n2435, S3 
                           => n2591, Z => n2692);
   U2230 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2693, Z => n1405);
   U2231 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1025, D1 => n2442, S1 
                           => n2589, D2 => n2438, S2 => n2590, D3 => n2435, S3 
                           => n2593, Z => n2693);
   U2232 : HS65_LHS_XOR2X3 port map( A => n2628, B => n2694, Z => n1404);
   U2233 : HS65_LH_MX41X4 port map( D0 => n1024, S0 => n2421, D1 => n2442, S1 
                           => n2591, D2 => n2438, S2 => n2592, D3 => n2595, S3 
                           => n2434, Z => n2694);
   U2234 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2695, Z => n1403);
   U2235 : HS65_LH_MX41X4 port map( D0 => n1023, S0 => n2421, D1 => n2442, S1 
                           => n2593, D2 => n2595, S2 => n2437, D3 => n2597, S3 
                           => n2434, Z => n2695);
   U2236 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2696, Z => n1402);
   U2237 : HS65_LH_MX41X4 port map( D0 => n1022, S0 => n2420, D1 => n2595, S1 
                           => n2441, D2 => n2597, S2 => n2437, D3 => n2599, S3 
                           => n2434, Z => n2696);
   U2238 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2697, Z => n1401);
   U2239 : HS65_LH_MX41X4 port map( D0 => n1021, S0 => n2420, D1 => n2597, S1 
                           => n2441, D2 => n2599, S2 => n2437, D3 => n2435, S3 
                           => n2601, Z => n2697);
   U2240 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2698, Z => n1400);
   U2241 : HS65_LH_MX41X4 port map( D0 => n1020, S0 => n2420, D1 => n2599, S1 
                           => n2441, D2 => n2438, S2 => n2600, D3 => n2435, S3 
                           => n2603, Z => n2698);
   U2242 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2699, Z => n1399);
   U2243 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1019, D1 => n2442, S1 
                           => n2601, D2 => n2438, S2 => n2602, D3 => n2435, S3 
                           => n2605, Z => n2699);
   U2244 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2700, Z => n1398);
   U2245 : HS65_LH_MX41X4 port map( D0 => n1018, S0 => n2420, D1 => n2442, S1 
                           => n2603, D2 => n2438, S2 => n2604, D3 => n2607, S3 
                           => n2435, Z => n2700);
   U2246 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2701, Z => n1397);
   U2247 : HS65_LH_MX41X4 port map( D0 => n1017, S0 => n2420, D1 => n2442, S1 
                           => n2605, D2 => n2607, S2 => n2438, D3 => n2609, S3 
                           => n2434, Z => n2701);
   U2248 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2702, Z => n1396);
   U2249 : HS65_LH_MX41X4 port map( D0 => n1016, S0 => n2420, D1 => n2607, S1 
                           => n2442, D2 => n2609, S2 => n2438, D3 => n2611, S3 
                           => n2435, Z => n2702);
   U2250 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2703, Z => n1395);
   U2251 : HS65_LH_MX41X4 port map( D0 => n1015, S0 => n2421, D1 => n2609, S1 
                           => n2442, D2 => n2611, S2 => n2438, D3 => n2435, S3 
                           => n2613, Z => n2703);
   U2252 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2704, Z => n1394);
   U2253 : HS65_LH_MX41X4 port map( D0 => n1014, S0 => n2420, D1 => n2611, S1 
                           => n2442, D2 => n2439, S2 => n2612, D3 => n2435, S3 
                           => n2615, Z => n2704);
   U2254 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2705, Z => n1393);
   U2255 : HS65_LH_MX41X4 port map( D0 => n2422, S0 => n1013, D1 => n2443, S1 
                           => n2613, D2 => n2438, S2 => n2614, D3 => n2435, S3 
                           => n2617, Z => n2705);
   U2256 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2706, Z => n1392);
   U2257 : HS65_LH_MX41X4 port map( D0 => n1012, S0 => n2420, D1 => n2443, S1 
                           => n2615, D2 => n2439, S2 => n2616, D3 => n2619, S3 
                           => n2435, Z => n2706);
   U2258 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2707, Z => n1391);
   U2259 : HS65_LH_MX41X4 port map( D0 => n1011, S0 => n2420, D1 => n2443, S1 
                           => n2617, D2 => n2619, S2 => n2438, D3 => n2621, S3 
                           => n2435, Z => n2707);
   U2260 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2708, Z => n1390);
   U2261 : HS65_LH_MX41X4 port map( D0 => n1010, S0 => n2420, D1 => n2619, S1 
                           => n2442, D2 => n2621, S2 => n2438, D3 => n2623, S3 
                           => n2435, Z => n2708);
   U2262 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2709, Z => n1389);
   U2263 : HS65_LH_MX41X4 port map( D0 => n1009, S0 => n2420, D1 => n2621, S1 
                           => n2442, D2 => n2623, S2 => n2438, D3 => n2625, S3 
                           => n2435, Z => n2709);
   U2264 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2710, Z => n1388);
   U2265 : HS65_LH_MX41X4 port map( D0 => n1008, S0 => n2420, D1 => n2623, S1 
                           => n2442, D2 => n2625, S2 => n2438, D3 => n2435, S3 
                           => n2627, Z => n2710);
   U2266 : HS65_LH_NOR2AX3 port map( A => a(0), B => n2711, Z => n2677);
   U2267 : HS65_LHS_XOR2X3 port map( A => n2629, B => n2712, Z => n1387);
   U2268 : HS65_LH_OAI12X2 port map( A => n2667, B => n2713, C => n2714, Z => 
                           n2712);
   U2269 : HS65_LH_OAI22X1 port map( A => n2625, B => n2715, C => n2441, D => 
                           n2715, Z => n2714);
   U2270 : HS65_LH_AND2X4 port map( A => n2438, B => n2626, Z => n2715);
   U2271 : HS65_LH_NOR2AX3 port map( A => a(1), B => a(0), Z => n2679);
   U2272 : HS65_LHS_XOR2X3 port map( A => n2630, B => n2716, Z => n1386);
   U2273 : HS65_LH_AOI22X1 port map( A => n2422, B => n1006, C => n2443, D => 
                           n2627, Z => n2716);
   U2274 : HS65_LH_NOR3AX2 port map( A => n2711, B => a(0), C => a(1), Z => 
                           n2681);
   U2275 : HS65_LH_NAND2X2 port map( A => a(0), B => n2711, Z => n2713);
   U2276 : HS65_LHS_XOR2X3 port map( A => n2629, B => a(1), Z => n2711);
   U2277 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2717, Z => n1384);
   U2278 : HS65_LH_AO22X4 port map( A => n2565, B => n2446, C => n2564, D => 
                           n2719, Z => n2717);
   U2279 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2720, Z => n1383);
   U2280 : HS65_LH_AO222X4 port map( A => n2567, B => n2446, C => n2563, D => 
                           n2450, E => n1038, F => n2448, Z => n2720);
   U2281 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2722, Z => n1382);
   U2282 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1037, D1 => n2455, S1 
                           => n2564, D2 => n2450, S2 => n2566, D3 => n2446, S3 
                           => n2569, Z => n2722);
   U2283 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2724, Z => n1381);
   U2284 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1036, D1 => n2454, S1 
                           => n2567, D2 => n2450, S2 => n2568, D3 => n2446, S3 
                           => n2571, Z => n2724);
   U2285 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2725, Z => n1380);
   U2286 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1035, D1 => n2454, S1 
                           => n2569, D2 => n2450, S2 => n2570, D3 => n2446, S3 
                           => n2573, Z => n2725);
   U2287 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2726, Z => n1379);
   U2288 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1034, D1 => n2454, S1 
                           => n2571, D2 => n2450, S2 => n2572, D3 => n2446, S3 
                           => n2575, Z => n2726);
   U2289 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2727, Z => n1378);
   U2290 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1033, D1 => n2454, S1 
                           => n2573, D2 => n2450, S2 => n2574, D3 => n2446, S3 
                           => n2577, Z => n2727);
   U2291 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2728, Z => n1377);
   U2292 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1032, D1 => n2454, S1 
                           => n2575, D2 => n2450, S2 => n2576, D3 => n2446, S3 
                           => n2579, Z => n2728);
   U2293 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2729, Z => n1376);
   U2294 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1031, D1 => n2454, S1 
                           => n2577, D2 => n2450, S2 => n2578, D3 => n2446, S3 
                           => n2581, Z => n2729);
   U2295 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2730, Z => n1375);
   U2296 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1030, D1 => n2454, S1 
                           => n2579, D2 => n2451, S2 => n2580, D3 => n2446, S3 
                           => n2583, Z => n2730);
   U2297 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2731, Z => n1374);
   U2298 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1029, D1 => n2454, S1 
                           => n2581, D2 => n2450, S2 => n2582, D3 => n2446, S3 
                           => n2585, Z => n2731);
   U2299 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2732, Z => n1373);
   U2300 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1028, D1 => n2454, S1 
                           => n2583, D2 => n2450, S2 => n2584, D3 => n2446, S3 
                           => n2587, Z => n2732);
   U2301 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2733, Z => n1372);
   U2302 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1027, D1 => n2454, S1 
                           => n2585, D2 => n2450, S2 => n2586, D3 => n2446, S3 
                           => n2589, Z => n2733);
   U2303 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2734, Z => n1371);
   U2304 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1026, D1 => n2454, S1 
                           => n2587, D2 => n2451, S2 => n2588, D3 => n2446, S3 
                           => n2591, Z => n2734);
   U2305 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2735, Z => n1370);
   U2306 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1025, D1 => n2454, S1 
                           => n2589, D2 => n2451, S2 => n2590, D3 => n2446, S3 
                           => n2592, Z => n2735);
   U2307 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2736, Z => n1369);
   U2308 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1024, D1 => n2455, S1 
                           => n2591, D2 => n2451, S2 => n2592, D3 => n2446, S3 
                           => n2595, Z => n2736);
   U2309 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2737, Z => n1368);
   U2310 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1023, D1 => n2455, S1 
                           => n2593, D2 => n2451, S2 => n2594, D3 => n2446, S3 
                           => n2597, Z => n2737);
   U2311 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2738, Z => n1367);
   U2312 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1022, D1 => n2455, S1 
                           => n2595, D2 => n2451, S2 => n2596, D3 => n2447, S3 
                           => n2599, Z => n2738);
   U2313 : HS65_LHS_XOR2X3 port map( A => n2631, B => n2739, Z => n1366);
   U2314 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1021, D1 => n2455, S1 
                           => n2597, D2 => n2451, S2 => n2598, D3 => n2447, S3 
                           => n2600, Z => n2739);
   U2315 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2740, Z => n1365);
   U2316 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1020, D1 => n2455, S1 
                           => n2599, D2 => n2451, S2 => n2600, D3 => n2447, S3 
                           => n2602, Z => n2740);
   U2317 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2741, Z => n1364);
   U2318 : HS65_LH_MX41X4 port map( D0 => n2448, S0 => n1019, D1 => n2455, S1 
                           => n2601, D2 => n2451, S2 => n2602, D3 => n2447, S3 
                           => n2604, Z => n2741);
   U2319 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2742, Z => n1363);
   U2320 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1018, D1 => n2455, S1 
                           => n2603, D2 => n2451, S2 => n2604, D3 => n2447, S3 
                           => n2607, Z => n2742);
   U2321 : HS65_LHS_XOR2X3 port map( A => a(5), B => n2743, Z => n1362);
   U2322 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1017, D1 => n2455, S1 
                           => n2605, D2 => n2451, S2 => n2606, D3 => n2447, S3 
                           => n2609, Z => n2743);
   U2323 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2744, Z => n1361);
   U2324 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1016, D1 => n2455, S1 
                           => n2607, D2 => n2451, S2 => n2608, D3 => n2447, S3 
                           => n2611, Z => n2744);
   U2325 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2745, Z => n1360);
   U2326 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1015, D1 => n2455, S1 
                           => n2609, D2 => n2451, S2 => n2610, D3 => n2447, S3 
                           => n2612, Z => n2745);
   U2327 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2746, Z => n1359);
   U2328 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1014, D1 => n2455, S1 
                           => n2611, D2 => n2451, S2 => n2612, D3 => n2447, S3 
                           => n2614, Z => n2746);
   U2329 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2747, Z => n1358);
   U2330 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1013, D1 => n2455, S1 
                           => n2613, D2 => n2452, S2 => n2614, D3 => n2447, S3 
                           => n2616, Z => n2747);
   U2331 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2748, Z => n1357);
   U2332 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1012, D1 => n2456, S1 
                           => n2615, D2 => n2452, S2 => n2616, D3 => n2447, S3 
                           => n2619, Z => n2748);
   U2333 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2749, Z => n1356);
   U2334 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1011, D1 => n2456, S1 
                           => n2617, D2 => n2452, S2 => n2618, D3 => n2447, S3 
                           => n2621, Z => n2749);
   U2335 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2750, Z => n1355);
   U2336 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1010, D1 => n2456, S1 
                           => n2619, D2 => n2452, S2 => n2620, D3 => n2447, S3 
                           => n2623, Z => n2750);
   U2337 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2751, Z => n1354);
   U2338 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1009, D1 => n2456, S1 
                           => n2621, D2 => n2452, S2 => n2622, D3 => n2447, S3 
                           => n2624, Z => n2751);
   U2339 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2752, Z => n1353);
   U2340 : HS65_LH_MX41X4 port map( D0 => n2719, S0 => n1008, D1 => n2456, S1 
                           => n2623, D2 => n2450, S2 => n2624, D3 => n2447, S3 
                           => n2627, Z => n2752);
   U2341 : HS65_LH_AND2X4 port map( A => n2753, B => n2754, Z => n2718);
   U2342 : HS65_LHS_XOR2X3 port map( A => n2632, B => n2755, Z => n1352);
   U2343 : HS65_LH_OAI12X2 port map( A => n2667, B => n2449, C => n2756, Z => 
                           n2755);
   U2344 : HS65_LH_OAI22X1 port map( A => n2625, B => n2757, C => n2454, D => 
                           n2757, Z => n2756);
   U2345 : HS65_LH_AND2X4 port map( A => n2450, B => n2626, Z => n2757);
   U2346 : HS65_LH_NOR2X2 port map( A => n2753, B => n2758, Z => n2721);
   U2347 : HS65_LHS_XOR2X3 port map( A => n2633, B => n2759, Z => n1351);
   U2348 : HS65_LH_AOI22X1 port map( A => n2719, B => n1006, C => n2456, D => 
                           n2627, Z => n2759);
   U2349 : HS65_LH_NOR3AX2 port map( A => n2758, B => n2754, C => n2753, Z => 
                           n2723);
   U2350 : HS65_LHS_XNOR2X3 port map( A => a(4), B => a(3), Z => n2758);
   U2351 : HS65_LH_NOR2AX3 port map( A => n2753, B => n2754, Z => n2719);
   U2352 : HS65_LHS_XNOR2X3 port map( A => n2632, B => a(4), Z => n2754);
   U2353 : HS65_LHS_XOR2X3 port map( A => n2628, B => a(3), Z => n2753);
   U2354 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2760, Z => n1349);
   U2355 : HS65_LH_AO22X4 port map( A => n2565, B => n2459, C => n2564, D => 
                           n2762, Z => n2760);
   U2356 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2763, Z => n1348);
   U2357 : HS65_LH_AO222X4 port map( A => n2567, B => n2459, C => n2563, D => 
                           n2463, E => n1038, F => n2461, Z => n2763);
   U2358 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2765, Z => n1347);
   U2359 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1037, D1 => n2468, S1 
                           => n2564, D2 => n2463, S2 => n2566, D3 => n2459, S3 
                           => n2569, Z => n2765);
   U2360 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2767, Z => n1346);
   U2361 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1036, D1 => n2467, S1 
                           => n2566, D2 => n2463, S2 => n2568, D3 => n2459, S3 
                           => n2571, Z => n2767);
   U2362 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2768, Z => n1345);
   U2363 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1035, D1 => n2467, S1 
                           => n2569, D2 => n2463, S2 => n2570, D3 => n2459, S3 
                           => n2573, Z => n2768);
   U2364 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2769, Z => n1344);
   U2365 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1034, D1 => n2467, S1 
                           => n2571, D2 => n2463, S2 => n2572, D3 => n2459, S3 
                           => n2575, Z => n2769);
   U2366 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2770, Z => n1343);
   U2367 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1033, D1 => n2467, S1 
                           => n2573, D2 => n2463, S2 => n2574, D3 => n2459, S3 
                           => n2577, Z => n2770);
   U2368 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2771, Z => n1342);
   U2369 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1032, D1 => n2467, S1 
                           => n2575, D2 => n2463, S2 => n2576, D3 => n2459, S3 
                           => n2579, Z => n2771);
   U2370 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2772, Z => n1341);
   U2371 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1031, D1 => n2467, S1 
                           => n2577, D2 => n2463, S2 => n2578, D3 => n2459, S3 
                           => n2581, Z => n2772);
   U2372 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2773, Z => n1340);
   U2373 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1030, D1 => n2467, S1 
                           => n2579, D2 => n2464, S2 => n2580, D3 => n2459, S3 
                           => n2583, Z => n2773);
   U2374 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2774, Z => n1339);
   U2375 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1029, D1 => n2467, S1 
                           => n2581, D2 => n2463, S2 => n2582, D3 => n2459, S3 
                           => n2585, Z => n2774);
   U2376 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2775, Z => n1338);
   U2377 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1028, D1 => n2467, S1 
                           => n2583, D2 => n2463, S2 => n2584, D3 => n2459, S3 
                           => n2587, Z => n2775);
   U2378 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2776, Z => n1337);
   U2379 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1027, D1 => n2467, S1 
                           => n2585, D2 => n2463, S2 => n2586, D3 => n2459, S3 
                           => n2589, Z => n2776);
   U2380 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2777, Z => n1336);
   U2381 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1026, D1 => n2467, S1 
                           => n2587, D2 => n2464, S2 => n2588, D3 => n2459, S3 
                           => n2591, Z => n2777);
   U2382 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2778, Z => n1335);
   U2383 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1025, D1 => n2467, S1 
                           => n2589, D2 => n2464, S2 => n2590, D3 => n2459, S3 
                           => n2593, Z => n2778);
   U2384 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2779, Z => n1334);
   U2385 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1024, D1 => n2468, S1 
                           => n2591, D2 => n2464, S2 => n2592, D3 => n2459, S3 
                           => n2595, Z => n2779);
   U2386 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2780, Z => n1333);
   U2387 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1023, D1 => n2468, S1 
                           => n2593, D2 => n2464, S2 => n2594, D3 => n2459, S3 
                           => n2597, Z => n2780);
   U2388 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2781, Z => n1332);
   U2389 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1022, D1 => n2468, S1 
                           => n2595, D2 => n2464, S2 => n2596, D3 => n2460, S3 
                           => n2599, Z => n2781);
   U2390 : HS65_LHS_XOR2X3 port map( A => n2634, B => n2782, Z => n1331);
   U2391 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1021, D1 => n2468, S1 
                           => n2597, D2 => n2464, S2 => n2598, D3 => n2460, S3 
                           => n2601, Z => n2782);
   U2392 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2783, Z => n1330);
   U2393 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1020, D1 => n2468, S1 
                           => n2599, D2 => n2464, S2 => n2600, D3 => n2460, S3 
                           => n2603, Z => n2783);
   U2394 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2784, Z => n1329);
   U2395 : HS65_LH_MX41X4 port map( D0 => n2461, S0 => n1019, D1 => n2468, S1 
                           => n2601, D2 => n2464, S2 => n2602, D3 => n2460, S3 
                           => n2605, Z => n2784);
   U2396 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2785, Z => n1328);
   U2397 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1018, D1 => n2468, S1 
                           => n2603, D2 => n2464, S2 => n2604, D3 => n2460, S3 
                           => n2607, Z => n2785);
   U2398 : HS65_LHS_XOR2X3 port map( A => a(8), B => n2786, Z => n1327);
   U2399 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1017, D1 => n2468, S1 
                           => n2605, D2 => n2464, S2 => n2606, D3 => n2460, S3 
                           => n2609, Z => n2786);
   U2400 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2787, Z => n1326);
   U2401 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1016, D1 => n2468, S1 
                           => n2607, D2 => n2464, S2 => n2608, D3 => n2460, S3 
                           => n2611, Z => n2787);
   U2402 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2788, Z => n1325);
   U2403 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1015, D1 => n2468, S1 
                           => n2609, D2 => n2464, S2 => n2610, D3 => n2460, S3 
                           => n2613, Z => n2788);
   U2404 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2789, Z => n1324);
   U2405 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1014, D1 => n2468, S1 
                           => n2611, D2 => n2464, S2 => n2612, D3 => n2460, S3 
                           => n2615, Z => n2789);
   U2406 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2790, Z => n1323);
   U2407 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1013, D1 => n2468, S1 
                           => n2613, D2 => n2465, S2 => n2614, D3 => n2460, S3 
                           => n2617, Z => n2790);
   U2408 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2791, Z => n1322);
   U2409 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1012, D1 => n2469, S1 
                           => n2615, D2 => n2465, S2 => n2616, D3 => n2460, S3 
                           => n2619, Z => n2791);
   U2410 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2792, Z => n1321);
   U2411 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1011, D1 => n2469, S1 
                           => n2617, D2 => n2465, S2 => n2618, D3 => n2460, S3 
                           => n2621, Z => n2792);
   U2412 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2793, Z => n1320);
   U2413 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1010, D1 => n2469, S1 
                           => n2619, D2 => n2465, S2 => n2620, D3 => n2460, S3 
                           => n2623, Z => n2793);
   U2414 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2794, Z => n1319);
   U2415 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1009, D1 => n2469, S1 
                           => n2621, D2 => n2465, S2 => n2622, D3 => n2460, S3 
                           => n2624, Z => n2794);
   U2416 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2795, Z => n1318);
   U2417 : HS65_LH_MX41X4 port map( D0 => n2762, S0 => n1008, D1 => n2469, S1 
                           => n2623, D2 => n2463, S2 => n2624, D3 => n2460, S3 
                           => n2627, Z => n2795);
   U2418 : HS65_LH_AND2X4 port map( A => n2796, B => n2797, Z => n2761);
   U2419 : HS65_LHS_XOR2X3 port map( A => n2635, B => n2798, Z => n1317);
   U2420 : HS65_LH_OAI12X2 port map( A => n2667, B => n2462, C => n2799, Z => 
                           n2798);
   U2421 : HS65_LH_OAI22X1 port map( A => n2625, B => n2800, C => n2467, D => 
                           n2800, Z => n2799);
   U2422 : HS65_LH_AND2X4 port map( A => n2463, B => n2626, Z => n2800);
   U2423 : HS65_LH_NOR2X2 port map( A => n2796, B => n2801, Z => n2764);
   U2424 : HS65_LHS_XOR2X3 port map( A => n2636, B => n2802, Z => n1316);
   U2425 : HS65_LH_AOI22X1 port map( A => n2762, B => n1006, C => n2469, D => 
                           n2627, Z => n2802);
   U2426 : HS65_LH_NOR3AX2 port map( A => n2801, B => n2797, C => n2796, Z => 
                           n2766);
   U2427 : HS65_LHS_XNOR2X3 port map( A => a(7), B => a(6), Z => n2801);
   U2428 : HS65_LH_NOR2AX3 port map( A => n2796, B => n2797, Z => n2762);
   U2429 : HS65_LHS_XNOR2X3 port map( A => n2635, B => a(7), Z => n2797);
   U2430 : HS65_LHS_XOR2X3 port map( A => n2631, B => a(6), Z => n2796);
   U2431 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2803, Z => n1314);
   U2432 : HS65_LH_AO22X4 port map( A => n2565, B => n2472, C => n2564, D => 
                           n2805, Z => n2803);
   U2433 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2806, Z => n1313);
   U2434 : HS65_LH_AO222X4 port map( A => n2567, B => n2472, C => n2563, D => 
                           n2476, E => n1038, F => n2474, Z => n2806);
   U2435 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2808, Z => n1312);
   U2436 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1037, D1 => n2472, S1 
                           => n2569, D2 => n2477, S2 => n2566, D3 => n2481, S3 
                           => n2564, Z => n2808);
   U2437 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2810, Z => n1311);
   U2438 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1036, D1 => n2472, S1 
                           => n2571, D2 => n2476, S2 => n2568, D3 => n2480, S3 
                           => n2566, Z => n2810);
   U2439 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2811, Z => n1310);
   U2440 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1035, D1 => n2472, S1 
                           => n2573, D2 => n2476, S2 => n2570, D3 => n2480, S3 
                           => n2569, Z => n2811);
   U2441 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2812, Z => n1309);
   U2442 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1034, D1 => n2472, S1 
                           => n2575, D2 => n2476, S2 => n2572, D3 => n2480, S3 
                           => n2571, Z => n2812);
   U2443 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2813, Z => n1308);
   U2444 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1033, D1 => n2472, S1 
                           => n2577, D2 => n2476, S2 => n2574, D3 => n2480, S3 
                           => n2573, Z => n2813);
   U2445 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2814, Z => n1307);
   U2446 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1032, D1 => n2472, S1 
                           => n2579, D2 => n2476, S2 => n2576, D3 => n2480, S3 
                           => n2575, Z => n2814);
   U2447 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2815, Z => n1306);
   U2448 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1031, D1 => n2472, S1 
                           => n2581, D2 => n2476, S2 => n2578, D3 => n2480, S3 
                           => n2577, Z => n2815);
   U2449 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2816, Z => n1305);
   U2450 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1030, D1 => n2472, S1 
                           => n2583, D2 => n2477, S2 => n2580, D3 => n2480, S3 
                           => n2579, Z => n2816);
   U2451 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2817, Z => n1304);
   U2452 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1029, D1 => n2472, S1 
                           => n2585, D2 => n2476, S2 => n2582, D3 => n2480, S3 
                           => n2581, Z => n2817);
   U2453 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2818, Z => n1303);
   U2454 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1028, D1 => n2472, S1 
                           => n2587, D2 => n2477, S2 => n2584, D3 => n2480, S3 
                           => n2583, Z => n2818);
   U2455 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2819, Z => n1302);
   U2456 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1027, D1 => n2472, S1 
                           => n2589, D2 => n2477, S2 => n2586, D3 => n2480, S3 
                           => n2585, Z => n2819);
   U2457 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2820, Z => n1301);
   U2458 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1026, D1 => n2472, S1 
                           => n2591, D2 => n2477, S2 => n2588, D3 => n2480, S3 
                           => n2587, Z => n2820);
   U2459 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2821, Z => n1300);
   U2460 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1025, D1 => n2472, S1 
                           => n2593, D2 => n2477, S2 => n2590, D3 => n2480, S3 
                           => n2589, Z => n2821);
   U2461 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2822, Z => n1299);
   U2462 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1024, D1 => n2476, S1 
                           => n2593, D2 => n2473, S2 => n2594, D3 => n2481, S3 
                           => n2591, Z => n2822);
   U2463 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2823, Z => n1298);
   U2464 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1023, D1 => n2476, S1 
                           => n2595, D2 => n2473, S2 => n2596, D3 => n2481, S3 
                           => n2593, Z => n2823);
   U2465 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2824, Z => n1297);
   U2466 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1022, D1 => n2473, S1 
                           => n2599, D2 => n2477, S2 => n2596, D3 => n2481, S3 
                           => n2595, Z => n2824);
   U2467 : HS65_LHS_XOR2X3 port map( A => n2637, B => n2825, Z => n1296);
   U2468 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1021, D1 => n2473, S1 
                           => n2601, D2 => n2477, S2 => n2598, D3 => n2481, S3 
                           => n2597, Z => n2825);
   U2469 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2826, Z => n1295);
   U2470 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1020, D1 => n2472, S1 
                           => n2603, D2 => n2477, S2 => n2600, D3 => n2481, S3 
                           => n2599, Z => n2826);
   U2471 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2827, Z => n1294);
   U2472 : HS65_LH_MX41X4 port map( D0 => n2474, S0 => n1019, D1 => n2473, S1 
                           => n2605, D2 => n2477, S2 => n2602, D3 => n2481, S3 
                           => n2601, Z => n2827);
   U2473 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2828, Z => n1293);
   U2474 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1018, D1 => n2473, S1 
                           => n2607, D2 => n2477, S2 => n2604, D3 => n2481, S3 
                           => n2603, Z => n2828);
   U2475 : HS65_LHS_XOR2X3 port map( A => a(11), B => n2829, Z => n1292);
   U2476 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1017, D1 => n2473, S1 
                           => n2609, D2 => n2477, S2 => n2606, D3 => n2481, S3 
                           => n2605, Z => n2829);
   U2477 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2830, Z => n1291);
   U2478 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1016, D1 => n2473, S1 
                           => n2611, D2 => n2477, S2 => n2608, D3 => n2481, S3 
                           => n2607, Z => n2830);
   U2479 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2831, Z => n1290);
   U2480 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1015, D1 => n2473, S1 
                           => n2613, D2 => n2477, S2 => n2610, D3 => n2481, S3 
                           => n2609, Z => n2831);
   U2481 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2832, Z => n1289);
   U2482 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1014, D1 => n2473, S1 
                           => n2615, D2 => n2478, S2 => n2612, D3 => n2481, S3 
                           => n2611, Z => n2832);
   U2483 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2833, Z => n1288);
   U2484 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1013, D1 => n2473, S1 
                           => n2617, D2 => n2478, S2 => n2614, D3 => n2481, S3 
                           => n2613, Z => n2833);
   U2485 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2834, Z => n1287);
   U2486 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1012, D1 => n2473, S1 
                           => n2619, D2 => n2478, S2 => n2616, D3 => n2482, S3 
                           => n2615, Z => n2834);
   U2487 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2835, Z => n1286);
   U2488 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1011, D1 => n2473, S1 
                           => n2621, D2 => n2478, S2 => n2618, D3 => n2482, S3 
                           => n2617, Z => n2835);
   U2489 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2836, Z => n1285);
   U2490 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1010, D1 => n2473, S1 
                           => n2623, D2 => n2478, S2 => n2620, D3 => n2482, S3 
                           => n2619, Z => n2836);
   U2491 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2837, Z => n1284);
   U2492 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1009, D1 => n2473, S1 
                           => n2624, D2 => n2476, S2 => n2622, D3 => n2482, S3 
                           => n2621, Z => n2837);
   U2493 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2838, Z => n1283);
   U2494 : HS65_LH_MX41X4 port map( D0 => n2805, S0 => n1008, D1 => n2476, S1 
                           => n2624, D2 => n2473, S2 => n2626, D3 => n2482, S3 
                           => n2623, Z => n2838);
   U2495 : HS65_LH_AND2X4 port map( A => n2839, B => n2840, Z => n2804);
   U2496 : HS65_LHS_XOR2X3 port map( A => n2638, B => n2841, Z => n1282);
   U2497 : HS65_LH_OAI12X2 port map( A => n2667, B => n2475, C => n2842, Z => 
                           n2841);
   U2498 : HS65_LH_OAI22X1 port map( A => n2625, B => n2843, C => n2480, D => 
                           n2843, Z => n2842);
   U2499 : HS65_LH_AND2X4 port map( A => n2476, B => n2626, Z => n2843);
   U2500 : HS65_LH_NOR2X2 port map( A => n2839, B => n2844, Z => n2807);
   U2501 : HS65_LHS_XOR2X3 port map( A => n2639, B => n2845, Z => n1281);
   U2502 : HS65_LH_AOI22X1 port map( A => n2805, B => n1006, C => n2482, D => 
                           n2627, Z => n2845);
   U2503 : HS65_LH_NOR3AX2 port map( A => n2844, B => n2840, C => n2839, Z => 
                           n2809);
   U2504 : HS65_LHS_XNOR2X3 port map( A => a(9), B => a(10), Z => n2844);
   U2505 : HS65_LH_NOR2AX3 port map( A => n2839, B => n2840, Z => n2805);
   U2506 : HS65_LHS_XNOR2X3 port map( A => n2638, B => a(10), Z => n2840);
   U2507 : HS65_LHS_XOR2X3 port map( A => n2634, B => a(9), Z => n2839);
   U2508 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2846, Z => n1279);
   U2509 : HS65_LH_AO22X4 port map( A => n2565, B => n2485, C => n2564, D => 
                           n2848, Z => n2846);
   U2510 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2849, Z => n1278);
   U2511 : HS65_LH_AO222X4 port map( A => n2567, B => n2485, C => n2563, D => 
                           n2489, E => n1038, F => n2487, Z => n2849);
   U2512 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2851, Z => n1277);
   U2513 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1037, D1 => n2494, S1 
                           => n2563, D2 => n2489, S2 => n2566, D3 => n2485, S3 
                           => n2569, Z => n2851);
   U2514 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2853, Z => n1276);
   U2515 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1036, D1 => n2493, S1 
                           => n2566, D2 => n2489, S2 => n2568, D3 => n2485, S3 
                           => n2571, Z => n2853);
   U2516 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2854, Z => n1275);
   U2517 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1035, D1 => n2493, S1 
                           => n2569, D2 => n2489, S2 => n2570, D3 => n2485, S3 
                           => n2573, Z => n2854);
   U2518 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2855, Z => n1274);
   U2519 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1034, D1 => n2493, S1 
                           => n2571, D2 => n2489, S2 => n2572, D3 => n2485, S3 
                           => n2575, Z => n2855);
   U2520 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2856, Z => n1273);
   U2521 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1033, D1 => n2493, S1 
                           => n2573, D2 => n2489, S2 => n2574, D3 => n2485, S3 
                           => n2577, Z => n2856);
   U2522 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2857, Z => n1272);
   U2523 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1032, D1 => n2493, S1 
                           => n2575, D2 => n2489, S2 => n2576, D3 => n2485, S3 
                           => n2579, Z => n2857);
   U2524 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2858, Z => n1271);
   U2525 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1031, D1 => n2493, S1 
                           => n2577, D2 => n2489, S2 => n2578, D3 => n2485, S3 
                           => n2581, Z => n2858);
   U2526 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2859, Z => n1270);
   U2527 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1030, D1 => n2493, S1 
                           => n2579, D2 => n2490, S2 => n2580, D3 => n2485, S3 
                           => n2583, Z => n2859);
   U2528 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2860, Z => n1269);
   U2529 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1029, D1 => n2493, S1 
                           => n2581, D2 => n2489, S2 => n2582, D3 => n2485, S3 
                           => n2585, Z => n2860);
   U2530 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2861, Z => n1268);
   U2531 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1028, D1 => n2493, S1 
                           => n2583, D2 => n2489, S2 => n2584, D3 => n2485, S3 
                           => n2587, Z => n2861);
   U2532 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2862, Z => n1267);
   U2533 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1027, D1 => n2493, S1 
                           => n2585, D2 => n2489, S2 => n2586, D3 => n2485, S3 
                           => n2589, Z => n2862);
   U2534 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2863, Z => n1266);
   U2535 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1026, D1 => n2493, S1 
                           => n2587, D2 => n2490, S2 => n2588, D3 => n2485, S3 
                           => n2591, Z => n2863);
   U2536 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2864, Z => n1265);
   U2537 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1025, D1 => n2493, S1 
                           => n2589, D2 => n2490, S2 => n2590, D3 => n2485, S3 
                           => n2593, Z => n2864);
   U2538 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2865, Z => n1264);
   U2539 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1024, D1 => n2494, S1 
                           => n2591, D2 => n2490, S2 => n2592, D3 => n2485, S3 
                           => n2595, Z => n2865);
   U2540 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2866, Z => n1263);
   U2541 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1023, D1 => n2494, S1 
                           => n2593, D2 => n2490, S2 => n2594, D3 => n2485, S3 
                           => n2597, Z => n2866);
   U2542 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2867, Z => n1262);
   U2543 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1022, D1 => n2494, S1 
                           => n2595, D2 => n2490, S2 => n2596, D3 => n2486, S3 
                           => n2599, Z => n2867);
   U2544 : HS65_LHS_XOR2X3 port map( A => n2640, B => n2868, Z => n1261);
   U2545 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1021, D1 => n2494, S1 
                           => n2597, D2 => n2490, S2 => n2598, D3 => n2486, S3 
                           => n2601, Z => n2868);
   U2546 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2869, Z => n1260);
   U2547 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1020, D1 => n2494, S1 
                           => n2599, D2 => n2490, S2 => n2600, D3 => n2486, S3 
                           => n2603, Z => n2869);
   U2548 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2870, Z => n1259);
   U2549 : HS65_LH_MX41X4 port map( D0 => n2487, S0 => n1019, D1 => n2494, S1 
                           => n2601, D2 => n2490, S2 => n2602, D3 => n2486, S3 
                           => n2605, Z => n2870);
   U2550 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2871, Z => n1258);
   U2551 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1018, D1 => n2494, S1 
                           => n2603, D2 => n2490, S2 => n2604, D3 => n2486, S3 
                           => n2607, Z => n2871);
   U2552 : HS65_LHS_XOR2X3 port map( A => a(14), B => n2872, Z => n1257);
   U2553 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1017, D1 => n2494, S1 
                           => n2605, D2 => n2490, S2 => n2606, D3 => n2486, S3 
                           => n2609, Z => n2872);
   U2554 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2873, Z => n1256);
   U2555 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1016, D1 => n2494, S1 
                           => n2607, D2 => n2490, S2 => n2608, D3 => n2486, S3 
                           => n2611, Z => n2873);
   U2556 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2874, Z => n1255);
   U2557 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1015, D1 => n2494, S1 
                           => n2609, D2 => n2490, S2 => n2610, D3 => n2486, S3 
                           => n2613, Z => n2874);
   U2558 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2875, Z => n1254);
   U2559 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1014, D1 => n2494, S1 
                           => n2611, D2 => n2490, S2 => n2612, D3 => n2486, S3 
                           => n2615, Z => n2875);
   U2560 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2876, Z => n1253);
   U2561 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1013, D1 => n2494, S1 
                           => n2613, D2 => n2491, S2 => n2614, D3 => n2486, S3 
                           => n2617, Z => n2876);
   U2562 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2877, Z => n1252);
   U2563 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1012, D1 => n2495, S1 
                           => n2615, D2 => n2491, S2 => n2616, D3 => n2486, S3 
                           => n2619, Z => n2877);
   U2564 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2878, Z => n1251);
   U2565 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1011, D1 => n2495, S1 
                           => n2617, D2 => n2491, S2 => n2618, D3 => n2486, S3 
                           => n2621, Z => n2878);
   U2566 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2879, Z => n1250);
   U2567 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1010, D1 => n2495, S1 
                           => n2619, D2 => n2491, S2 => n2620, D3 => n2486, S3 
                           => n2623, Z => n2879);
   U2568 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2880, Z => n1249);
   U2569 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1009, D1 => n2495, S1 
                           => n2621, D2 => n2491, S2 => n2622, D3 => n2486, S3 
                           => n2624, Z => n2880);
   U2570 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2881, Z => n1248);
   U2571 : HS65_LH_MX41X4 port map( D0 => n2848, S0 => n1008, D1 => n2495, S1 
                           => n2623, D2 => n2489, S2 => n2624, D3 => n2486, S3 
                           => n2627, Z => n2881);
   U2572 : HS65_LH_AND2X4 port map( A => n2882, B => n2883, Z => n2847);
   U2573 : HS65_LHS_XOR2X3 port map( A => n2641, B => n2884, Z => n1247);
   U2574 : HS65_LH_OAI12X2 port map( A => n2667, B => n2488, C => n2885, Z => 
                           n2884);
   U2575 : HS65_LH_OAI22X1 port map( A => n2625, B => n2886, C => n2493, D => 
                           n2886, Z => n2885);
   U2576 : HS65_LH_AND2X4 port map( A => n2489, B => n2626, Z => n2886);
   U2577 : HS65_LH_NOR2X2 port map( A => n2882, B => n2887, Z => n2850);
   U2578 : HS65_LHS_XOR2X3 port map( A => n2642, B => n2888, Z => n1246);
   U2579 : HS65_LH_AOI22X1 port map( A => n2848, B => n1006, C => n2495, D => 
                           n2627, Z => n2888);
   U2580 : HS65_LH_NOR3AX2 port map( A => n2887, B => n2883, C => n2882, Z => 
                           n2852);
   U2581 : HS65_LHS_XNOR2X3 port map( A => a(13), B => a(12), Z => n2887);
   U2582 : HS65_LH_NOR2AX3 port map( A => n2882, B => n2883, Z => n2848);
   U2583 : HS65_LHS_XNOR2X3 port map( A => n2641, B => a(13), Z => n2883);
   U2584 : HS65_LHS_XOR2X3 port map( A => n2637, B => a(12), Z => n2882);
   U2585 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2889, Z => n1244);
   U2586 : HS65_LH_AO22X4 port map( A => n2564, B => n2498, C => n2564, D => 
                           n2891, Z => n2889);
   U2587 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2892, Z => n1243);
   U2588 : HS65_LH_AO222X4 port map( A => n2567, B => n2498, C => n2563, D => 
                           n2502, E => n1038, F => n2500, Z => n2892);
   U2589 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2894, Z => n1242);
   U2590 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1037, D1 => n2507, S1 
                           => n2563, D2 => n2502, S2 => n2566, D3 => n2498, S3 
                           => n2569, Z => n2894);
   U2591 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2896, Z => n1241);
   U2592 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1036, D1 => n2506, S1 
                           => n2566, D2 => n2502, S2 => n2568, D3 => n2498, S3 
                           => n2571, Z => n2896);
   U2593 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2897, Z => n1240);
   U2594 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1035, D1 => n2506, S1 
                           => n2568, D2 => n2502, S2 => n2570, D3 => n2498, S3 
                           => n2573, Z => n2897);
   U2595 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2898, Z => n1239);
   U2596 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1034, D1 => n2506, S1 
                           => n2570, D2 => n2502, S2 => n2572, D3 => n2498, S3 
                           => n2575, Z => n2898);
   U2597 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2899, Z => n1238);
   U2598 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1033, D1 => n2506, S1 
                           => n2572, D2 => n2502, S2 => n2574, D3 => n2498, S3 
                           => n2577, Z => n2899);
   U2599 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2900, Z => n1237);
   U2600 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1032, D1 => n2506, S1 
                           => n2574, D2 => n2502, S2 => n2576, D3 => n2498, S3 
                           => n2579, Z => n2900);
   U2601 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2901, Z => n1236);
   U2602 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1031, D1 => n2506, S1 
                           => n2576, D2 => n2502, S2 => n2578, D3 => n2498, S3 
                           => n2581, Z => n2901);
   U2603 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2902, Z => n1235);
   U2604 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1030, D1 => n2506, S1 
                           => n2578, D2 => n2503, S2 => n2580, D3 => n2498, S3 
                           => n2583, Z => n2902);
   U2605 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2903, Z => n1234);
   U2606 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1029, D1 => n2506, S1 
                           => n2580, D2 => n2502, S2 => n2582, D3 => n2498, S3 
                           => n2585, Z => n2903);
   U2607 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2904, Z => n1233);
   U2608 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1028, D1 => n2506, S1 
                           => n2582, D2 => n2502, S2 => n2584, D3 => n2498, S3 
                           => n2587, Z => n2904);
   U2609 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2905, Z => n1232);
   U2610 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1027, D1 => n2506, S1 
                           => n2584, D2 => n2502, S2 => n2586, D3 => n2498, S3 
                           => n2589, Z => n2905);
   U2611 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2906, Z => n1231);
   U2612 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1026, D1 => n2506, S1 
                           => n2586, D2 => n2503, S2 => n2588, D3 => n2498, S3 
                           => n2591, Z => n2906);
   U2613 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2907, Z => n1230);
   U2614 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1025, D1 => n2506, S1 
                           => n2589, D2 => n2503, S2 => n2590, D3 => n2498, S3 
                           => n2593, Z => n2907);
   U2615 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2908, Z => n1229);
   U2616 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1024, D1 => n2507, S1 
                           => n2591, D2 => n2503, S2 => n2592, D3 => n2498, S3 
                           => n2595, Z => n2908);
   U2617 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2909, Z => n1228);
   U2618 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1023, D1 => n2507, S1 
                           => n2593, D2 => n2503, S2 => n2594, D3 => n2498, S3 
                           => n2597, Z => n2909);
   U2619 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2910, Z => n1227);
   U2620 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1022, D1 => n2507, S1 
                           => n2594, D2 => n2503, S2 => n2596, D3 => n2499, S3 
                           => n2599, Z => n2910);
   U2621 : HS65_LHS_XOR2X3 port map( A => n2643, B => n2911, Z => n1226);
   U2622 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1021, D1 => n2507, S1 
                           => n2597, D2 => n2503, S2 => n2598, D3 => n2499, S3 
                           => n2601, Z => n2911);
   U2623 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2912, Z => n1225);
   U2624 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1020, D1 => n2507, S1 
                           => n2598, D2 => n2503, S2 => n2600, D3 => n2499, S3 
                           => n2603, Z => n2912);
   U2625 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2913, Z => n1224);
   U2626 : HS65_LH_MX41X4 port map( D0 => n2500, S0 => n1019, D1 => n2507, S1 
                           => n2601, D2 => n2503, S2 => n2602, D3 => n2499, S3 
                           => n2605, Z => n2913);
   U2627 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2914, Z => n1223);
   U2628 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1018, D1 => n2507, S1 
                           => n2603, D2 => n2503, S2 => n2604, D3 => n2499, S3 
                           => n2607, Z => n2914);
   U2629 : HS65_LHS_XOR2X3 port map( A => a(17), B => n2915, Z => n1222);
   U2630 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1017, D1 => n2507, S1 
                           => n2605, D2 => n2503, S2 => n2606, D3 => n2499, S3 
                           => n2609, Z => n2915);
   U2631 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2916, Z => n1221);
   U2632 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1016, D1 => n2507, S1 
                           => n2606, D2 => n2503, S2 => n2608, D3 => n2499, S3 
                           => n2611, Z => n2916);
   U2633 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2917, Z => n1220);
   U2634 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1015, D1 => n2507, S1 
                           => n2608, D2 => n2503, S2 => n2610, D3 => n2499, S3 
                           => n2613, Z => n2917);
   U2635 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2918, Z => n1219);
   U2636 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1014, D1 => n2507, S1 
                           => n2610, D2 => n2503, S2 => n2612, D3 => n2499, S3 
                           => n2615, Z => n2918);
   U2637 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2919, Z => n1218);
   U2638 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1013, D1 => n2507, S1 
                           => n2613, D2 => n2504, S2 => n2614, D3 => n2499, S3 
                           => n2617, Z => n2919);
   U2639 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2920, Z => n1217);
   U2640 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1012, D1 => n2508, S1 
                           => n2615, D2 => n2504, S2 => n2616, D3 => n2499, S3 
                           => n2619, Z => n2920);
   U2641 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2921, Z => n1216);
   U2642 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1011, D1 => n2508, S1 
                           => n2617, D2 => n2504, S2 => n2618, D3 => n2499, S3 
                           => n2621, Z => n2921);
   U2643 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2922, Z => n1215);
   U2644 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1010, D1 => n2508, S1 
                           => n2618, D2 => n2504, S2 => n2620, D3 => n2499, S3 
                           => n2623, Z => n2922);
   U2645 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2923, Z => n1214);
   U2646 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1009, D1 => n2508, S1 
                           => n2620, D2 => n2504, S2 => n2622, D3 => n2499, S3 
                           => n2624, Z => n2923);
   U2647 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2924, Z => n1213);
   U2648 : HS65_LH_MX41X4 port map( D0 => n2891, S0 => n1008, D1 => n2508, S1 
                           => n2622, D2 => n2502, S2 => n2624, D3 => n2499, S3 
                           => n2626, Z => n2924);
   U2649 : HS65_LH_AND2X4 port map( A => n2925, B => n2926, Z => n2890);
   U2650 : HS65_LHS_XOR2X3 port map( A => n2644, B => n2927, Z => n1212);
   U2651 : HS65_LH_OAI12X2 port map( A => n2667, B => n2501, C => n2928, Z => 
                           n2927);
   U2652 : HS65_LH_OAI22X1 port map( A => n2625, B => n2929, C => n2506, D => 
                           n2929, Z => n2928);
   U2653 : HS65_LH_AND2X4 port map( A => n2502, B => n2626, Z => n2929);
   U2654 : HS65_LH_NOR2X2 port map( A => n2925, B => n2930, Z => n2893);
   U2655 : HS65_LHS_XOR2X3 port map( A => n2645, B => n2931, Z => n1211);
   U2656 : HS65_LH_AOI22X1 port map( A => n2891, B => n1006, C => n2508, D => 
                           n2627, Z => n2931);
   U2657 : HS65_LH_NOR3AX2 port map( A => n2930, B => n2926, C => n2925, Z => 
                           n2895);
   U2658 : HS65_LHS_XNOR2X3 port map( A => a(16), B => a(15), Z => n2930);
   U2659 : HS65_LH_NOR2AX3 port map( A => n2925, B => n2926, Z => n2891);
   U2660 : HS65_LHS_XNOR2X3 port map( A => n2644, B => a(16), Z => n2926);
   U2661 : HS65_LHS_XOR2X3 port map( A => n2640, B => a(15), Z => n2925);
   U2662 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2932, Z => n1209);
   U2663 : HS65_LH_AO22X4 port map( A => n2565, B => n2511, C => n2564, D => 
                           n2934, Z => n2932);
   U2664 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2935, Z => n1208);
   U2665 : HS65_LH_AO222X4 port map( A => n2567, B => n2511, C => n2563, D => 
                           n2515, E => n1038, F => n2513, Z => n2935);
   U2666 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2937, Z => n1207);
   U2667 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1037, D1 => n2520, S1 
                           => n2564, D2 => n2515, S2 => n2566, D3 => n2511, S3 
                           => n2568, Z => n2937);
   U2668 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2939, Z => n1206);
   U2669 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1036, D1 => n2519, S1 
                           => n2566, D2 => n2515, S2 => n2568, D3 => n2511, S3 
                           => n2570, Z => n2939);
   U2670 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2940, Z => n1205);
   U2671 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1035, D1 => n2519, S1 
                           => n2568, D2 => n2515, S2 => n2570, D3 => n2511, S3 
                           => n2572, Z => n2940);
   U2672 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2941, Z => n1204);
   U2673 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1034, D1 => n2519, S1 
                           => n2570, D2 => n2515, S2 => n2572, D3 => n2511, S3 
                           => n2574, Z => n2941);
   U2674 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2942, Z => n1203);
   U2675 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1033, D1 => n2519, S1 
                           => n2572, D2 => n2515, S2 => n2574, D3 => n2511, S3 
                           => n2576, Z => n2942);
   U2676 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2943, Z => n1202);
   U2677 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1032, D1 => n2519, S1 
                           => n2574, D2 => n2515, S2 => n2576, D3 => n2511, S3 
                           => n2578, Z => n2943);
   U2678 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2944, Z => n1201);
   U2679 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1031, D1 => n2519, S1 
                           => n2576, D2 => n2515, S2 => n2578, D3 => n2511, S3 
                           => n2580, Z => n2944);
   U2680 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2945, Z => n1200);
   U2681 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1030, D1 => n2519, S1 
                           => n2578, D2 => n2516, S2 => n2580, D3 => n2511, S3 
                           => n2582, Z => n2945);
   U2682 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2946, Z => n1199);
   U2683 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1029, D1 => n2519, S1 
                           => n2580, D2 => n2515, S2 => n2582, D3 => n2511, S3 
                           => n2584, Z => n2946);
   U2684 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2947, Z => n1198);
   U2685 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1028, D1 => n2519, S1 
                           => n2582, D2 => n2515, S2 => n2584, D3 => n2511, S3 
                           => n2586, Z => n2947);
   U2686 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2948, Z => n1197);
   U2687 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1027, D1 => n2519, S1 
                           => n2584, D2 => n2515, S2 => n2586, D3 => n2511, S3 
                           => n2589, Z => n2948);
   U2688 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2949, Z => n1196);
   U2689 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1026, D1 => n2519, S1 
                           => n2586, D2 => n2516, S2 => n2588, D3 => n2511, S3 
                           => n2591, Z => n2949);
   U2690 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2950, Z => n1195);
   U2691 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1025, D1 => n2519, S1 
                           => n2588, D2 => n2516, S2 => n2590, D3 => n2511, S3 
                           => n2592, Z => n2950);
   U2692 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2951, Z => n1194);
   U2693 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1024, D1 => n2520, S1 
                           => n2590, D2 => n2516, S2 => n2592, D3 => n2511, S3 
                           => n2594, Z => n2951);
   U2694 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2952, Z => n1193);
   U2695 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1023, D1 => n2520, S1 
                           => n2592, D2 => n2516, S2 => n2594, D3 => n2511, S3 
                           => n2596, Z => n2952);
   U2696 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2953, Z => n1192);
   U2697 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1022, D1 => n2520, S1 
                           => n2594, D2 => n2516, S2 => n2596, D3 => n2512, S3 
                           => n2598, Z => n2953);
   U2698 : HS65_LHS_XOR2X3 port map( A => n2646, B => n2954, Z => n1191);
   U2699 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1021, D1 => n2520, S1 
                           => n2596, D2 => n2516, S2 => n2598, D3 => n2512, S3 
                           => n2601, Z => n2954);
   U2700 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2955, Z => n1190);
   U2701 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1020, D1 => n2520, S1 
                           => n2598, D2 => n2516, S2 => n2600, D3 => n2512, S3 
                           => n2603, Z => n2955);
   U2702 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2956, Z => n1189);
   U2703 : HS65_LH_MX41X4 port map( D0 => n2513, S0 => n1019, D1 => n2520, S1 
                           => n2600, D2 => n2516, S2 => n2602, D3 => n2512, S3 
                           => n2605, Z => n2956);
   U2704 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2957, Z => n1188);
   U2705 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1018, D1 => n2520, S1 
                           => n2602, D2 => n2516, S2 => n2604, D3 => n2512, S3 
                           => n2606, Z => n2957);
   U2706 : HS65_LHS_XOR2X3 port map( A => a(20), B => n2958, Z => n1187);
   U2707 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1017, D1 => n2520, S1 
                           => n2604, D2 => n2516, S2 => n2606, D3 => n2512, S3 
                           => n2608, Z => n2958);
   U2708 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2959, Z => n1186);
   U2709 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1016, D1 => n2520, S1 
                           => n2606, D2 => n2516, S2 => n2608, D3 => n2512, S3 
                           => n2610, Z => n2959);
   U2710 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2960, Z => n1185);
   U2711 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1015, D1 => n2520, S1 
                           => n2608, D2 => n2516, S2 => n2610, D3 => n2512, S3 
                           => n2613, Z => n2960);
   U2712 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2961, Z => n1184);
   U2713 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1014, D1 => n2520, S1 
                           => n2610, D2 => n2516, S2 => n2612, D3 => n2512, S3 
                           => n2615, Z => n2961);
   U2714 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2962, Z => n1183);
   U2715 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1013, D1 => n2520, S1 
                           => n2612, D2 => n2517, S2 => n2614, D3 => n2512, S3 
                           => n2617, Z => n2962);
   U2716 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2963, Z => n1182);
   U2717 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1012, D1 => n2521, S1 
                           => n2614, D2 => n2517, S2 => n2616, D3 => n2512, S3 
                           => n2618, Z => n2963);
   U2718 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2964, Z => n1181);
   U2719 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1011, D1 => n2521, S1 
                           => n2616, D2 => n2517, S2 => n2618, D3 => n2512, S3 
                           => n2620, Z => n2964);
   U2720 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2965, Z => n1180);
   U2721 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1010, D1 => n2521, S1 
                           => n2618, D2 => n2517, S2 => n2620, D3 => n2512, S3 
                           => n2622, Z => n2965);
   U2722 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2966, Z => n1179);
   U2723 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1009, D1 => n2521, S1 
                           => n2620, D2 => n2517, S2 => n2622, D3 => n2512, S3 
                           => n2624, Z => n2966);
   U2724 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2967, Z => n1178);
   U2725 : HS65_LH_MX41X4 port map( D0 => n2934, S0 => n1008, D1 => n2521, S1 
                           => n2622, D2 => n2515, S2 => n2624, D3 => n2512, S3 
                           => n2626, Z => n2967);
   U2726 : HS65_LH_AND2X4 port map( A => n2968, B => n2969, Z => n2933);
   U2727 : HS65_LHS_XOR2X3 port map( A => n2647, B => n2970, Z => n1177);
   U2728 : HS65_LH_OAI12X2 port map( A => n2667, B => n2514, C => n2971, Z => 
                           n2970);
   U2729 : HS65_LH_OAI22X1 port map( A => n2625, B => n2972, C => n2519, D => 
                           n2972, Z => n2971);
   U2730 : HS65_LH_AND2X4 port map( A => n2515, B => n2626, Z => n2972);
   U2731 : HS65_LH_NOR2X2 port map( A => n2968, B => n2973, Z => n2936);
   U2732 : HS65_LHS_XOR2X3 port map( A => n2648, B => n2974, Z => n1176);
   U2733 : HS65_LH_AOI22X1 port map( A => n2934, B => n1006, C => n2521, D => 
                           n2627, Z => n2974);
   U2734 : HS65_LH_NOR3AX2 port map( A => n2973, B => n2969, C => n2968, Z => 
                           n2938);
   U2735 : HS65_LHS_XNOR2X3 port map( A => a(19), B => a(18), Z => n2973);
   U2736 : HS65_LH_NOR2AX3 port map( A => n2968, B => n2969, Z => n2934);
   U2737 : HS65_LHS_XNOR2X3 port map( A => n2647, B => a(19), Z => n2969);
   U2738 : HS65_LHS_XOR2X3 port map( A => n2643, B => a(18), Z => n2968);
   U2739 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2975, Z => n1174);
   U2740 : HS65_LH_AO22X4 port map( A => n2565, B => n2524, C => n2564, D => 
                           n2977, Z => n2975);
   U2741 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2978, Z => n1173);
   U2742 : HS65_LH_AO222X4 port map( A => n2567, B => n2524, C => n2563, D => 
                           n2528, E => n1038, F => n2526, Z => n2978);
   U2743 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2980, Z => n1172);
   U2744 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1037, D1 => n2524, S1 
                           => n2568, D2 => n2533, S2 => n2563, D3 => n2528, S3 
                           => n2566, Z => n2980);
   U2745 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2982, Z => n1171);
   U2746 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1036, D1 => n2524, S1 
                           => n2570, D2 => n2532, S2 => n2566, D3 => n2528, S3 
                           => n2568, Z => n2982);
   U2747 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2983, Z => n1170);
   U2748 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1035, D1 => n2524, S1 
                           => n2572, D2 => n2532, S2 => n2568, D3 => n2528, S3 
                           => n2570, Z => n2983);
   U2749 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2984, Z => n1169);
   U2750 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1034, D1 => n2524, S1 
                           => n2574, D2 => n2532, S2 => n2570, D3 => n2528, S3 
                           => n2572, Z => n2984);
   U2751 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2985, Z => n1168);
   U2752 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1033, D1 => n2524, S1 
                           => n2576, D2 => n2532, S2 => n2572, D3 => n2528, S3 
                           => n2574, Z => n2985);
   U2753 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2986, Z => n1167);
   U2754 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1032, D1 => n2524, S1 
                           => n2578, D2 => n2532, S2 => n2574, D3 => n2528, S3 
                           => n2576, Z => n2986);
   U2755 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2987, Z => n1166);
   U2756 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1031, D1 => n2524, S1 
                           => n2580, D2 => n2532, S2 => n2576, D3 => n2528, S3 
                           => n2578, Z => n2987);
   U2757 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2988, Z => n1165);
   U2758 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1030, D1 => n2524, S1 
                           => n2582, D2 => n2532, S2 => n2578, D3 => n2529, S3 
                           => n2580, Z => n2988);
   U2759 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2989, Z => n1164);
   U2760 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1029, D1 => n2524, S1 
                           => n2584, D2 => n2532, S2 => n2580, D3 => n2528, S3 
                           => n2582, Z => n2989);
   U2761 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2990, Z => n1163);
   U2762 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1028, D1 => n2524, S1 
                           => n2586, D2 => n2532, S2 => n2582, D3 => n2528, S3 
                           => n2584, Z => n2990);
   U2763 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2991, Z => n1162);
   U2764 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1027, D1 => n2524, S1 
                           => n2588, D2 => n2532, S2 => n2584, D3 => n2528, S3 
                           => n2586, Z => n2991);
   U2765 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2992, Z => n1161);
   U2766 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1026, D1 => n2524, S1 
                           => n2590, D2 => n2532, S2 => n2586, D3 => n2529, S3 
                           => n2588, Z => n2992);
   U2767 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2993, Z => n1160);
   U2768 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1025, D1 => n2524, S1 
                           => n2592, D2 => n2532, S2 => n2588, D3 => n2529, S3 
                           => n2590, Z => n2993);
   U2769 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2994, Z => n1159);
   U2770 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1024, D1 => n2524, S1 
                           => n2594, D2 => n2533, S2 => n2590, D3 => n2529, S3 
                           => n2592, Z => n2994);
   U2771 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2995, Z => n1158);
   U2772 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1023, D1 => n2525, S1 
                           => n2596, D2 => n2533, S2 => n2592, D3 => n2529, S3 
                           => n2594, Z => n2995);
   U2773 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2996, Z => n1157);
   U2774 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1022, D1 => n2525, S1 
                           => n2598, D2 => n2533, S2 => n2594, D3 => n2529, S3 
                           => n2596, Z => n2996);
   U2775 : HS65_LHS_XOR2X3 port map( A => n2649, B => n2997, Z => n1156);
   U2776 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1021, D1 => n2525, S1 
                           => n2600, D2 => n2533, S2 => n2596, D3 => n2529, S3 
                           => n2598, Z => n2997);
   U2777 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2998, Z => n1155);
   U2778 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1020, D1 => n2525, S1 
                           => n2602, D2 => n2533, S2 => n2598, D3 => n2529, S3 
                           => n2600, Z => n2998);
   U2779 : HS65_LHS_XOR2X3 port map( A => a(23), B => n2999, Z => n1154);
   U2780 : HS65_LH_MX41X4 port map( D0 => n2526, S0 => n1019, D1 => n2525, S1 
                           => n2604, D2 => n2533, S2 => n2600, D3 => n2529, S3 
                           => n2602, Z => n2999);
   U2781 : HS65_LHS_XOR2X3 port map( A => a(23), B => n3000, Z => n1153);
   U2782 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1018, D1 => n2525, S1 
                           => n2606, D2 => n2533, S2 => n2602, D3 => n2529, S3 
                           => n2604, Z => n3000);
   U2783 : HS65_LHS_XOR2X3 port map( A => a(23), B => n3001, Z => n1152);
   U2784 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1017, D1 => n2525, S1 
                           => n2608, D2 => n2533, S2 => n2604, D3 => n2529, S3 
                           => n2606, Z => n3001);
   U2785 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3002, Z => n1151);
   U2786 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1016, D1 => n2525, S1 
                           => n2610, D2 => n2533, S2 => n2606, D3 => n2529, S3 
                           => n2608, Z => n3002);
   U2787 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3003, Z => n1150);
   U2788 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1015, D1 => n2525, S1 
                           => n2612, D2 => n2533, S2 => n2608, D3 => n2529, S3 
                           => n2610, Z => n3003);
   U2789 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3004, Z => n1149);
   U2790 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1014, D1 => n2525, S1 
                           => n2614, D2 => n2533, S2 => n2610, D3 => n2529, S3 
                           => n2612, Z => n3004);
   U2791 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3005, Z => n1148);
   U2792 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1013, D1 => n2525, S1 
                           => n2616, D2 => n2533, S2 => n2612, D3 => n2530, S3 
                           => n2614, Z => n3005);
   U2793 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3006, Z => n1147);
   U2794 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1012, D1 => n2525, S1 
                           => n2618, D2 => n2533, S2 => n2614, D3 => n2530, S3 
                           => n2616, Z => n3006);
   U2795 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3007, Z => n1146);
   U2796 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1011, D1 => n2525, S1 
                           => n2620, D2 => n2534, S2 => n2616, D3 => n2530, S3 
                           => n2618, Z => n3007);
   U2797 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3008, Z => n1145);
   U2798 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1010, D1 => n2525, S1 
                           => n2622, D2 => n2534, S2 => n2618, D3 => n2530, S3 
                           => n2620, Z => n3008);
   U2799 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3009, Z => n1144);
   U2800 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1009, D1 => n2525, S1 
                           => n2624, D2 => n2534, S2 => n2620, D3 => n2530, S3 
                           => n2622, Z => n3009);
   U2801 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3010, Z => n1143);
   U2802 : HS65_LH_MX41X4 port map( D0 => n2977, S0 => n1008, D1 => n2525, S1 
                           => n2626, D2 => n2534, S2 => n2622, D3 => n2528, S3 
                           => n2624, Z => n3010);
   U2803 : HS65_LH_AND2X4 port map( A => n3011, B => n3012, Z => n2976);
   U2804 : HS65_LHS_XOR2X3 port map( A => n2650, B => n3013, Z => n1142);
   U2805 : HS65_LH_OAI12X2 port map( A => n2667, B => n2527, C => n3014, Z => 
                           n3013);
   U2806 : HS65_LH_OAI22X1 port map( A => n2625, B => n3015, C => n2532, D => 
                           n3015, Z => n3014);
   U2807 : HS65_LH_AND2X4 port map( A => n2528, B => n2626, Z => n3015);
   U2808 : HS65_LH_NOR2X2 port map( A => n3011, B => n3016, Z => n2979);
   U2809 : HS65_LHS_XOR2X3 port map( A => n2651, B => n3017, Z => n1141);
   U2810 : HS65_LH_AOI22X1 port map( A => n2977, B => n1006, C => n2534, D => 
                           n2627, Z => n3017);
   U2811 : HS65_LH_NOR3AX2 port map( A => n3016, B => n3012, C => n3011, Z => 
                           n2981);
   U2812 : HS65_LHS_XNOR2X3 port map( A => a(22), B => a(21), Z => n3016);
   U2813 : HS65_LH_NOR2AX3 port map( A => n3011, B => n3012, Z => n2977);
   U2814 : HS65_LHS_XNOR2X3 port map( A => n2650, B => a(22), Z => n3012);
   U2815 : HS65_LHS_XOR2X3 port map( A => n2646, B => a(21), Z => n3011);
   U2816 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3018, Z => n1139);
   U2817 : HS65_LH_AO22X4 port map( A => n2565, B => n2537, C => n2564, D => 
                           n3020, Z => n3018);
   U2818 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3021, Z => n1138);
   U2819 : HS65_LH_AO222X4 port map( A => n2567, B => n2537, C => n2563, D => 
                           n2541, E => n1038, F => n2539, Z => n3021);
   U2820 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3023, Z => n1137);
   U2821 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1037, D1 => n2546, S1 
                           => n2563, D2 => n2541, S2 => n2566, D3 => n2537, S3 
                           => n2568, Z => n3023);
   U2822 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3025, Z => n1136);
   U2823 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1036, D1 => n2545, S1 
                           => n2567, D2 => n2541, S2 => n2568, D3 => n2537, S3 
                           => n2570, Z => n3025);
   U2824 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3026, Z => n1135);
   U2825 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1035, D1 => n2545, S1 
                           => n2568, D2 => n2541, S2 => n2570, D3 => n2537, S3 
                           => n2572, Z => n3026);
   U2826 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3027, Z => n1134);
   U2827 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1034, D1 => n2545, S1 
                           => n2570, D2 => n2541, S2 => n2572, D3 => n2537, S3 
                           => n2574, Z => n3027);
   U2828 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3028, Z => n1133);
   U2829 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1033, D1 => n2545, S1 
                           => n2572, D2 => n2541, S2 => n2574, D3 => n2537, S3 
                           => n2576, Z => n3028);
   U2830 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3029, Z => n1132);
   U2831 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1032, D1 => n2545, S1 
                           => n2574, D2 => n2541, S2 => n2576, D3 => n2537, S3 
                           => n2578, Z => n3029);
   U2832 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3030, Z => n1131);
   U2833 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1031, D1 => n2545, S1 
                           => n2576, D2 => n2541, S2 => n2578, D3 => n2537, S3 
                           => n2580, Z => n3030);
   U2834 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3031, Z => n1130);
   U2835 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1030, D1 => n2545, S1 
                           => n2578, D2 => n2542, S2 => n2580, D3 => n2537, S3 
                           => n2582, Z => n3031);
   U2836 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3032, Z => n1129);
   U2837 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1029, D1 => n2545, S1 
                           => n2580, D2 => n2541, S2 => n2582, D3 => n2537, S3 
                           => n2584, Z => n3032);
   U2838 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3033, Z => n1128);
   U2839 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1028, D1 => n2545, S1 
                           => n2582, D2 => n2541, S2 => n2584, D3 => n2537, S3 
                           => n2586, Z => n3033);
   U2840 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3034, Z => n1127);
   U2841 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1027, D1 => n2545, S1 
                           => n2584, D2 => n2541, S2 => n2586, D3 => n2537, S3 
                           => n2588, Z => n3034);
   U2842 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3035, Z => n1126);
   U2843 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1026, D1 => n2545, S1 
                           => n2586, D2 => n2542, S2 => n2588, D3 => n2537, S3 
                           => n2590, Z => n3035);
   U2844 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3036, Z => n1125);
   U2845 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1025, D1 => n2545, S1 
                           => n2588, D2 => n2542, S2 => n2590, D3 => n2537, S3 
                           => n2592, Z => n3036);
   U2846 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3037, Z => n1124);
   U2847 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1024, D1 => n2546, S1 
                           => n2590, D2 => n2542, S2 => n2592, D3 => n2537, S3 
                           => n2594, Z => n3037);
   U2848 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3038, Z => n1123);
   U2849 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1023, D1 => n2546, S1 
                           => n2592, D2 => n2542, S2 => n2594, D3 => n2537, S3 
                           => n2596, Z => n3038);
   U2850 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3039, Z => n1122);
   U2851 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1022, D1 => n2546, S1 
                           => n2594, D2 => n2542, S2 => n2596, D3 => n2538, S3 
                           => n2598, Z => n3039);
   U2852 : HS65_LHS_XOR2X3 port map( A => n2652, B => n3040, Z => n1121);
   U2853 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1021, D1 => n2546, S1 
                           => n2596, D2 => n2542, S2 => n2598, D3 => n2538, S3 
                           => n2600, Z => n3040);
   U2854 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3041, Z => n1120);
   U2855 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1020, D1 => n2546, S1 
                           => n2598, D2 => n2542, S2 => n2600, D3 => n2538, S3 
                           => n2602, Z => n3041);
   U2856 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3042, Z => n1119);
   U2857 : HS65_LH_MX41X4 port map( D0 => n2539, S0 => n1019, D1 => n2546, S1 
                           => n2600, D2 => n2542, S2 => n2602, D3 => n2538, S3 
                           => n2604, Z => n3042);
   U2858 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3043, Z => n1118);
   U2859 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1018, D1 => n2546, S1 
                           => n2602, D2 => n2542, S2 => n2604, D3 => n2538, S3 
                           => n2606, Z => n3043);
   U2860 : HS65_LHS_XOR2X3 port map( A => a(26), B => n3044, Z => n1117);
   U2861 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1017, D1 => n2546, S1 
                           => n2604, D2 => n2542, S2 => n2606, D3 => n2538, S3 
                           => n2608, Z => n3044);
   U2862 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3045, Z => n1116);
   U2863 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1016, D1 => n2546, S1 
                           => n2606, D2 => n2542, S2 => n2608, D3 => n2538, S3 
                           => n2610, Z => n3045);
   U2864 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3046, Z => n1115);
   U2865 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1015, D1 => n2546, S1 
                           => n2608, D2 => n2542, S2 => n2610, D3 => n2538, S3 
                           => n2612, Z => n3046);
   U2866 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3047, Z => n1114);
   U2867 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1014, D1 => n2546, S1 
                           => n2610, D2 => n2542, S2 => n2612, D3 => n2538, S3 
                           => n2614, Z => n3047);
   U2868 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3048, Z => n1113);
   U2869 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1013, D1 => n2546, S1 
                           => n2612, D2 => n2543, S2 => n2614, D3 => n2538, S3 
                           => n2616, Z => n3048);
   U2870 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3049, Z => n1112);
   U2871 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1012, D1 => n2547, S1 
                           => n2614, D2 => n2543, S2 => n2616, D3 => n2538, S3 
                           => n2618, Z => n3049);
   U2872 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3050, Z => n1111);
   U2873 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1011, D1 => n2547, S1 
                           => n2616, D2 => n2543, S2 => n2618, D3 => n2538, S3 
                           => n2620, Z => n3050);
   U2874 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3051, Z => n1110);
   U2875 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1010, D1 => n2547, S1 
                           => n2618, D2 => n2543, S2 => n2620, D3 => n2538, S3 
                           => n2622, Z => n3051);
   U2876 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3052, Z => n1109);
   U2877 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1009, D1 => n2547, S1 
                           => n2620, D2 => n2543, S2 => n2622, D3 => n2538, S3 
                           => n2624, Z => n3052);
   U2878 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3053, Z => n1108);
   U2879 : HS65_LH_MX41X4 port map( D0 => n3020, S0 => n1008, D1 => n2547, S1 
                           => n2622, D2 => n2541, S2 => n2624, D3 => n2538, S3 
                           => n2626, Z => n3053);
   U2880 : HS65_LH_AND2X4 port map( A => n3054, B => n3055, Z => n3019);
   U2881 : HS65_LHS_XOR2X3 port map( A => n2653, B => n3056, Z => n1107);
   U2882 : HS65_LH_OAI12X2 port map( A => n2667, B => n2540, C => n3057, Z => 
                           n3056);
   U2883 : HS65_LH_OAI22X1 port map( A => n2625, B => n3058, C => n2545, D => 
                           n3058, Z => n3057);
   U2884 : HS65_LH_AND2X4 port map( A => n2541, B => n2626, Z => n3058);
   U2885 : HS65_LH_NOR2X2 port map( A => n3054, B => n3059, Z => n3022);
   U2886 : HS65_LHS_XOR2X3 port map( A => n2654, B => n3060, Z => n1106);
   U2887 : HS65_LH_AOI22X1 port map( A => n3020, B => n1006, C => n2547, D => 
                           n2627, Z => n3060);
   U2888 : HS65_LH_NOR3AX2 port map( A => n3059, B => n3055, C => n3054, Z => 
                           n3024);
   U2889 : HS65_LHS_XNOR2X3 port map( A => a(25), B => a(24), Z => n3059);
   U2890 : HS65_LH_NOR2AX3 port map( A => n3054, B => n3055, Z => n3020);
   U2891 : HS65_LHS_XNOR2X3 port map( A => n2653, B => a(25), Z => n3055);
   U2892 : HS65_LHS_XOR2X3 port map( A => n2649, B => a(24), Z => n3054);
   U2893 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3061, Z => n1104);
   U2894 : HS65_LH_AO22X4 port map( A => n2565, B => n2550, C => n2564, D => 
                           n3063, Z => n3061);
   U2895 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3064, Z => n1103);
   U2896 : HS65_LH_AO222X4 port map( A => n2567, B => n2550, C => n2563, D => 
                           n2554, E => n1038, F => n2552, Z => n3064);
   U2897 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3066, Z => n1102);
   U2898 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1037, D1 => n2559, S1 
                           => n2563, D2 => n2554, S2 => n2566, D3 => n2550, S3 
                           => n2568, Z => n3066);
   U2899 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3068, Z => n1101);
   U2900 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1036, D1 => n2558, S1 
                           => n2567, D2 => n2554, S2 => n2568, D3 => n2550, S3 
                           => n2570, Z => n3068);
   U2901 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3069, Z => n1100);
   U2902 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1035, D1 => n2558, S1 
                           => n2568, D2 => n2554, S2 => n2570, D3 => n2550, S3 
                           => n2572, Z => n3069);
   U2903 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3070, Z => n1099);
   U2904 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1034, D1 => n2558, S1 
                           => n2570, D2 => n2554, S2 => n2572, D3 => n2550, S3 
                           => n2574, Z => n3070);
   U2905 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3071, Z => n1098);
   U2906 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1033, D1 => n2558, S1 
                           => n2572, D2 => n2554, S2 => n2574, D3 => n2550, S3 
                           => n2576, Z => n3071);
   U2907 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3072, Z => n1097);
   U2908 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1032, D1 => n2558, S1 
                           => n2574, D2 => n2554, S2 => n2576, D3 => n2550, S3 
                           => n2578, Z => n3072);
   U2909 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3073, Z => n1096);
   U2910 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1031, D1 => n2558, S1 
                           => n2576, D2 => n2554, S2 => n2578, D3 => n2550, S3 
                           => n2580, Z => n3073);
   U2911 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3074, Z => n1095);
   U2912 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1030, D1 => n2558, S1 
                           => n2578, D2 => n2555, S2 => n2580, D3 => n2550, S3 
                           => n2582, Z => n3074);
   U2913 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3075, Z => n1094);
   U2914 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1029, D1 => n2558, S1 
                           => n2580, D2 => n2554, S2 => n2582, D3 => n2550, S3 
                           => n2584, Z => n3075);
   U2915 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3076, Z => n1093);
   U2916 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1028, D1 => n2558, S1 
                           => n2582, D2 => n2554, S2 => n2584, D3 => n2550, S3 
                           => n2586, Z => n3076);
   U2917 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3077, Z => n1092);
   U2918 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1027, D1 => n2558, S1 
                           => n2584, D2 => n2554, S2 => n2586, D3 => n2550, S3 
                           => n2588, Z => n3077);
   U2919 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3078, Z => n1091);
   U2920 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1026, D1 => n2558, S1 
                           => n2586, D2 => n2555, S2 => n2588, D3 => n2550, S3 
                           => n2590, Z => n3078);
   U2921 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3079, Z => n1090);
   U2922 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1025, D1 => n2558, S1 
                           => n2588, D2 => n2555, S2 => n2590, D3 => n2550, S3 
                           => n2592, Z => n3079);
   U2923 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3080, Z => n1089);
   U2924 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1024, D1 => n2559, S1 
                           => n2590, D2 => n2555, S2 => n2592, D3 => n2550, S3 
                           => n2594, Z => n3080);
   U2925 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3081, Z => n1088);
   U2926 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1023, D1 => n2559, S1 
                           => n2592, D2 => n2555, S2 => n2594, D3 => n2550, S3 
                           => n2596, Z => n3081);
   U2927 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3082, Z => n1087);
   U2928 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1022, D1 => n2559, S1 
                           => n2594, D2 => n2555, S2 => n2596, D3 => n2551, S3 
                           => n2598, Z => n3082);
   U2929 : HS65_LHS_XOR2X3 port map( A => n2655, B => n3083, Z => n1086);
   U2930 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1021, D1 => n2559, S1 
                           => n2596, D2 => n2555, S2 => n2598, D3 => n2551, S3 
                           => n2600, Z => n3083);
   U2931 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3084, Z => n1085);
   U2932 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1020, D1 => n2559, S1 
                           => n2598, D2 => n2555, S2 => n2600, D3 => n2551, S3 
                           => n2602, Z => n3084);
   U2933 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3085, Z => n1084);
   U2934 : HS65_LH_MX41X4 port map( D0 => n2552, S0 => n1019, D1 => n2559, S1 
                           => n2600, D2 => n2555, S2 => n2602, D3 => n2551, S3 
                           => n2604, Z => n3085);
   U2935 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3086, Z => n1083);
   U2936 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1018, D1 => n2559, S1 
                           => n2602, D2 => n2555, S2 => n2604, D3 => n2551, S3 
                           => n2606, Z => n3086);
   U2937 : HS65_LHS_XOR2X3 port map( A => a(29), B => n3087, Z => n1082);
   U2938 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1017, D1 => n2559, S1 
                           => n2604, D2 => n2555, S2 => n2606, D3 => n2551, S3 
                           => n2608, Z => n3087);
   U2939 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3088, Z => n1081);
   U2940 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1016, D1 => n2559, S1 
                           => n2606, D2 => n2555, S2 => n2608, D3 => n2551, S3 
                           => n2610, Z => n3088);
   U2941 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3089, Z => n1080);
   U2942 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1015, D1 => n2559, S1 
                           => n2608, D2 => n2555, S2 => n2610, D3 => n2551, S3 
                           => n2612, Z => n3089);
   U2943 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3090, Z => n1079);
   U2944 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1014, D1 => n2559, S1 
                           => n2610, D2 => n2555, S2 => n2612, D3 => n2551, S3 
                           => n2614, Z => n3090);
   U2945 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3091, Z => n1078);
   U2946 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1013, D1 => n2559, S1 
                           => n2612, D2 => n2556, S2 => n2614, D3 => n2551, S3 
                           => n2616, Z => n3091);
   U2947 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3092, Z => n1077);
   U2948 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1012, D1 => n2560, S1 
                           => n2614, D2 => n2556, S2 => n2616, D3 => n2551, S3 
                           => n2618, Z => n3092);
   U2949 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3093, Z => n1076);
   U2950 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1011, D1 => n2560, S1 
                           => n2616, D2 => n2556, S2 => n2618, D3 => n2551, S3 
                           => n2620, Z => n3093);
   U2951 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3094, Z => n1075);
   U2952 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1010, D1 => n2560, S1 
                           => n2618, D2 => n2556, S2 => n2620, D3 => n2551, S3 
                           => n2622, Z => n3094);
   U2953 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3095, Z => n1074);
   U2954 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1009, D1 => n2560, S1 
                           => n2620, D2 => n2556, S2 => n2622, D3 => n2551, S3 
                           => n2624, Z => n3095);
   U2955 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3096, Z => n1073);
   U2956 : HS65_LH_MX41X4 port map( D0 => n3063, S0 => n1008, D1 => n2560, S1 
                           => n2622, D2 => n2554, S2 => n2624, D3 => n2551, S3 
                           => n2626, Z => n3096);
   U2957 : HS65_LH_AND2X4 port map( A => n3097, B => n3098, Z => n3062);
   U2958 : HS65_LHS_XOR2X3 port map( A => n2656, B => n3099, Z => n1072);
   U2959 : HS65_LH_OAI12X2 port map( A => n2667, B => n2553, C => n3100, Z => 
                           n3099);
   U2960 : HS65_LH_OAI22X1 port map( A => n2625, B => n3101, C => n2558, D => 
                           n3101, Z => n3100);
   U2961 : HS65_LH_AND2X4 port map( A => n2554, B => n2626, Z => n3101);
   U2962 : HS65_LH_NOR2X2 port map( A => n3097, B => n3102, Z => n3065);
   U2963 : HS65_LHS_XOR2X3 port map( A => n2657, B => n3103, Z => n1071);
   U2964 : HS65_LH_AOI22X1 port map( A => n3063, B => n1006, C => n2560, D => 
                           n2627, Z => n3103);
   U2965 : HS65_LH_NOR3AX2 port map( A => n3102, B => n3098, C => n3097, Z => 
                           n3067);
   U2966 : HS65_LHS_XNOR2X3 port map( A => a(28), B => a(27), Z => n3102);
   U2967 : HS65_LH_NOR2AX3 port map( A => n3097, B => n3098, Z => n3063);
   U2968 : HS65_LHS_XNOR2X3 port map( A => n2656, B => a(28), Z => n3098);
   U2969 : HS65_LHS_XOR2X3 port map( A => n2652, B => a(27), Z => n3097);
   U2970 : HS65_LH_AO22X4 port map( A => n2428, B => n2563, C => n2419, D => 
                           n2564, Z => n1069);
   U2971 : HS65_LH_AO222X4 port map( A => n2428, B => n2566, C => n2432, D => 
                           n2563, E => n2419, F => n1038, Z => n1068);
   U2972 : HS65_LH_MX41X4 port map( D0 => n1037, S0 => n2419, D1 => n2569, S1 
                           => n2426, D2 => n2567, S2 => n2430, D3 => n2564, S3 
                           => n2423, Z => n1067);
   U2973 : HS65_LH_MX41X4 port map( D0 => n1036, S0 => n2419, D1 => n2571, S1 
                           => n2426, D2 => n2569, S2 => n2430, D3 => n2567, S3 
                           => n2423, Z => n1066);
   U2974 : HS65_LH_MX41X4 port map( D0 => n1035, S0 => n2419, D1 => n2573, S1 
                           => n2426, D2 => n2571, S2 => n2430, D3 => n2569, S3 
                           => n2423, Z => n1065);
   U2975 : HS65_LH_MX41X4 port map( D0 => n1034, S0 => n2418, D1 => n2575, S1 
                           => n2426, D2 => n2573, S2 => n2430, D3 => n2571, S3 
                           => n2423, Z => n1064);
   U2976 : HS65_LH_MX41X4 port map( D0 => n1033, S0 => n2418, D1 => n2577, S1 
                           => n2426, D2 => n2575, S2 => n2430, D3 => n2573, S3 
                           => n2423, Z => n1063);
   U2977 : HS65_LH_MX41X4 port map( D0 => n1032, S0 => n2418, D1 => n2579, S1 
                           => n2426, D2 => n2577, S2 => n2430, D3 => n2575, S3 
                           => n2423, Z => n1062);
   U2978 : HS65_LH_MX41X4 port map( D0 => n1031, S0 => n2418, D1 => n2581, S1 
                           => n2426, D2 => n2579, S2 => n2430, D3 => n2577, S3 
                           => n2423, Z => n1061);
   U2979 : HS65_LH_MX41X4 port map( D0 => n1030, S0 => n2418, D1 => n2583, S1 
                           => n2426, D2 => n2581, S2 => n2430, D3 => n2579, S3 
                           => n2423, Z => n1060);
   U2980 : HS65_LH_MX41X4 port map( D0 => n1029, S0 => n2418, D1 => n2585, S1 
                           => n2426, D2 => n2583, S2 => n2430, D3 => n2581, S3 
                           => n2423, Z => n1059);
   U2981 : HS65_LH_MX41X4 port map( D0 => n1028, S0 => n2418, D1 => n2587, S1 
                           => n2426, D2 => n2585, S2 => n2431, D3 => n2583, S3 
                           => n2424, Z => n1058);
   U2982 : HS65_LH_MX41X4 port map( D0 => n1027, S0 => n2418, D1 => n2428, S1 
                           => n2588, D2 => n2587, S2 => n2431, D3 => n2585, S3 
                           => n2424, Z => n1057);
   U2983 : HS65_LH_MX41X4 port map( D0 => n1026, S0 => n2418, D1 => n2428, S1 
                           => n2590, D2 => n2589, S2 => n2431, D3 => n2587, S3 
                           => n2424, Z => n1056);
   U2984 : HS65_LH_MX41X4 port map( D0 => n1024, S0 => n2418, D1 => n2593, S1 
                           => n2432, D2 => n2591, S2 => n2423, D3 => n2595, S3 
                           => n2426, Z => n1055);
   U2985 : HS65_LH_MX41X4 port map( D0 => n1023, S0 => n2418, D1 => n2593, S1 
                           => n2424, D2 => n2595, S2 => n2431, D3 => n2597, S3 
                           => n2427, Z => n1054);
   U2986 : HS65_LH_MX41X4 port map( D0 => n1022, S0 => n2417, D1 => n2595, S1 
                           => n2424, D2 => n2597, S2 => n2431, D3 => n2599, S3 
                           => n2427, Z => n1053);
   U2987 : HS65_LH_MX41X4 port map( D0 => n1021, S0 => n2417, D1 => n2597, S1 
                           => n2424, D2 => n2599, S2 => n2431, D3 => n2601, S3 
                           => n2427, Z => n1052);
   U2988 : HS65_LH_MX41X4 port map( D0 => n1020, S0 => n2417, D1 => n2599, S1 
                           => n2424, D2 => n2601, S2 => n2431, D3 => n2603, S3 
                           => n2427, Z => n1051);
   U2989 : HS65_LH_MX41X4 port map( D0 => n1018, S0 => n2417, D1 => n2603, S1 
                           => n2424, D2 => n2605, S2 => n2431, D3 => n2607, S3 
                           => n2427, Z => n1050);
   U2990 : HS65_LH_MX41X4 port map( D0 => n1017, S0 => n2417, D1 => n2605, S1 
                           => n2424, D2 => n2607, S2 => n2431, D3 => n2609, S3 
                           => n2427, Z => n1049);
   U2991 : HS65_LH_MX41X4 port map( D0 => n1016, S0 => n2417, D1 => n2607, S1 
                           => n2424, D2 => n2609, S2 => n2431, D3 => n2611, S3 
                           => n2427, Z => n1048);
   U2992 : HS65_LH_MX41X4 port map( D0 => n1015, S0 => n2417, D1 => n2609, S1 
                           => n2424, D2 => n2611, S2 => n2431, D3 => n2613, S3 
                           => n2427, Z => n1047);
   U2993 : HS65_LH_MX41X4 port map( D0 => n1014, S0 => n2417, D1 => n2611, S1 
                           => n2424, D2 => n2613, S2 => n2432, D3 => n2615, S3 
                           => n2427, Z => n1046);
   U2994 : HS65_LH_MX41X4 port map( D0 => n1012, S0 => n2417, D1 => n2615, S1 
                           => n2424, D2 => n2617, S2 => n2432, D3 => n2619, S3 
                           => n2427, Z => n1045);
   U2995 : HS65_LH_MX41X4 port map( D0 => n1011, S0 => n2417, D1 => n2617, S1 
                           => n2424, D2 => n2619, S2 => n2432, D3 => n2621, S3 
                           => n2427, Z => n1044);
   U2996 : HS65_LH_MX41X4 port map( D0 => n1010, S0 => n2417, D1 => n2619, S1 
                           => n2424, D2 => n2621, S2 => n2432, D3 => n2623, S3 
                           => n2427, Z => n1043);
   U2997 : HS65_LH_MX41X4 port map( D0 => n1009, S0 => n2417, D1 => n2621, S1 
                           => n2423, D2 => n2623, S2 => n2431, D3 => n2625, S3 
                           => n2428, Z => n1042);
   U2998 : HS65_LH_MX41X4 port map( D0 => n1008, S0 => n2418, D1 => n2623, S1 
                           => n2424, D2 => n2625, S2 => n2430, D3 => n2428, S3 
                           => n2626, Z => n1041);
   U2999 : HS65_LH_NOR2AX3 port map( A => n3104, B => a(31), Z => n2671);
   U3000 : HS65_LH_NOR2AX3 port map( A => n3105, B => n3104, Z => n2672);
   U3001 : HS65_LH_NOR3AX2 port map( A => a(31), B => n3105, C => n3104, Z => 
                           n2670);
   U3002 : HS65_LHS_XOR2X3 port map( A => a(31), B => a(30), Z => n3105);
   U3003 : HS65_LH_NAND2X2 port map( A => a(31), B => n3104, Z => n2673);
   U3004 : HS65_LHS_XOR2X3 port map( A => n2655, B => a(30), Z => n3104);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity if_top_DW01_inc_0 is

   port( A : in std_logic_vector (11 downto 0);  SUM : out std_logic_vector (11
         downto 0));

end if_top_DW01_inc_0;

architecture SYN_rpl of if_top_DW01_inc_0 is

   component HS65_LH_CNIVX3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_HA1X4
      port( A0, B0 : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   signal carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port : std_logic;

begin
   
   U1_1_10 : HS65_LH_HA1X4 port map( A0 => A(10), B0 => carry_10_port, CO => 
                           carry_11_port, S0 => SUM(10));
   U1_1_9 : HS65_LH_HA1X4 port map( A0 => A(9), B0 => carry_9_port, CO => 
                           carry_10_port, S0 => SUM(9));
   U1_1_8 : HS65_LH_HA1X4 port map( A0 => A(8), B0 => carry_8_port, CO => 
                           carry_9_port, S0 => SUM(8));
   U1_1_7 : HS65_LH_HA1X4 port map( A0 => A(7), B0 => carry_7_port, CO => 
                           carry_8_port, S0 => SUM(7));
   U1_1_6 : HS65_LH_HA1X4 port map( A0 => A(6), B0 => carry_6_port, CO => 
                           carry_7_port, S0 => SUM(6));
   U1_1_5 : HS65_LH_HA1X4 port map( A0 => A(5), B0 => carry_5_port, CO => 
                           carry_6_port, S0 => SUM(5));
   U1_1_4 : HS65_LH_HA1X4 port map( A0 => A(4), B0 => carry_4_port, CO => 
                           carry_5_port, S0 => SUM(4));
   U1_1_3 : HS65_LH_HA1X4 port map( A0 => A(3), B0 => carry_3_port, CO => 
                           carry_4_port, S0 => SUM(3));
   U1_1_2 : HS65_LH_HA1X4 port map( A0 => A(2), B0 => carry_2_port, CO => 
                           carry_3_port, S0 => SUM(2));
   U1_1_1 : HS65_LH_HA1X4 port map( A0 => A(1), B0 => A(0), CO => carry_2_port,
                           S0 => SUM(1));
   U1 : HS65_LHS_XOR2X3 port map( A => carry_11_port, B => A(11), Z => SUM(11))
                           ;
   U2 : HS65_LH_CNIVX3 port map( A => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_add_0;

architecture SYN_rpl of alu_DW01_add_0 is

   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1 : std_logic;

begin
   
   U1_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => B(23), CI => 
                           carry_23_port, CO => carry_24_port, S0 => SUM(23));
   U1_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => B(29), CI => 
                           carry_29_port, CO => carry_30_port, S0 => SUM(29));
   U1_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => B(26), CI => 
                           carry_26_port, CO => carry_27_port, S0 => SUM(26));
   U1_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => B(17), CI => 
                           carry_17_port, CO => carry_18_port, S0 => SUM(17));
   U1_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => B(5), CI => carry_5_port, 
                           CO => carry_6_port, S0 => SUM(5));
   U1_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => B(14), CI => 
                           carry_14_port, CO => carry_15_port, S0 => SUM(14));
   U1_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => B(8), CI => carry_8_port, 
                           CO => carry_9_port, S0 => SUM(8));
   U1_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => B(3), CI => carry_3_port, 
                           CO => carry_4_port, S0 => SUM(3));
   U1_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => B(1), CI => n1, CO => 
                           carry_2_port, S0 => SUM(1));
   U1_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => B(9), CI => carry_9_port, 
                           CO => carry_10_port, S0 => SUM(9));
   U1_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => B(7), CI => carry_7_port, 
                           CO => carry_8_port, S0 => SUM(7));
   U1_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => B(10), CI => 
                           carry_10_port, CO => carry_11_port, S0 => SUM(10));
   U1_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => B(6), CI => carry_6_port, 
                           CO => carry_7_port, S0 => SUM(6));
   U1_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => B(4), CI => carry_4_port, 
                           CO => carry_5_port, S0 => SUM(4));
   U1_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => B(30), CI => 
                           carry_30_port, CO => carry_31_port, S0 => SUM(30));
   U1_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => B(25), CI => 
                           carry_25_port, CO => carry_26_port, S0 => SUM(25));
   U1_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => B(19), CI => 
                           carry_19_port, CO => carry_20_port, S0 => SUM(19));
   U1_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => B(27), CI => 
                           carry_27_port, CO => carry_28_port, S0 => SUM(27));
   U1_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => B(24), CI => 
                           carry_24_port, CO => carry_25_port, S0 => SUM(24));
   U1_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => B(21), CI => 
                           carry_21_port, CO => carry_22_port, S0 => SUM(21));
   U1_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => B(18), CI => 
                           carry_18_port, CO => carry_19_port, S0 => SUM(18));
   U1_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => B(13), CI => 
                           carry_13_port, CO => carry_14_port, S0 => SUM(13));
   U1_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => B(12), CI => 
                           carry_12_port, CO => carry_13_port, S0 => SUM(12));
   U1_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => B(22), CI => 
                           carry_22_port, CO => carry_23_port, S0 => SUM(22));
   U1_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => B(15), CI => 
                           carry_15_port, CO => carry_16_port, S0 => SUM(15));
   U1_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => B(28), CI => 
                           carry_28_port, CO => carry_29_port, S0 => SUM(28));
   U1_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => B(16), CI => 
                           carry_16_port, CO => carry_17_port, S0 => SUM(16));
   U1_31 : HS65_LHS_XOR3X2 port map( A => A(31), B => B(31), C => carry_31_port
                           , Z => SUM(31));
   U1_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => B(2), CI => carry_2_port, 
                           CO => carry_3_port, S0 => SUM(2));
   U1_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => B(20), CI => 
                           carry_20_port, CO => carry_21_port, S0 => SUM(20));
   U1_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => B(11), CI => 
                           carry_11_port, CO => carry_12_port, S0 => SUM(11));
   U1 : HS65_LH_AND2X4 port map( A => A(0), B => B(0), Z => n1);
   U2 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => SUM(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end alu_DW01_cmp6_0;

architecture SYN_rpl of alu_DW01_cmp6_0 is

   component HS65_LH_NAND2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2AX4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND4X3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CNIVX3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal LT_port, EQ_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114 : std_logic;

begin
   LT <= LT_port;
   EQ <= EQ_port;
   
   U1 : HS65_LH_IVX9 port map( A => n114, Z => n39);
   U2 : HS65_LH_IVX9 port map( A => n53, Z => n34);
   U3 : HS65_LH_IVX9 port map( A => n101, Z => n37);
   U4 : HS65_LH_IVX9 port map( A => B(2), Z => n1);
   U5 : HS65_LH_IVX9 port map( A => A(14), Z => n21);
   U6 : HS65_LH_IVX9 port map( A => B(3), Z => n2);
   U7 : HS65_LH_IVX9 port map( A => B(11), Z => n6);
   U8 : HS65_LH_IVX9 port map( A => A(8), Z => n20);
   U9 : HS65_LH_IVX9 port map( A => A(26), Z => n22);
   U10 : HS65_LH_IVX9 port map( A => B(27), Z => n16);
   U11 : HS65_LH_IVX9 port map( A => B(20), Z => n12);
   U12 : HS65_LH_IVX9 port map( A => B(28), Z => n17);
   U13 : HS65_LH_IVX9 port map( A => B(31), Z => n19);
   U14 : HS65_LH_IVX9 port map( A => n66, Z => n26);
   U15 : HS65_LH_IVX9 port map( A => n75, Z => n23);
   U16 : HS65_LH_IVX9 port map( A => n59, Z => n24);
   U17 : HS65_LH_IVX9 port map( A => A(22), Z => n29);
   U18 : HS65_LH_IVX9 port map( A => n70, Z => n32);
   U19 : HS65_LH_IVX9 port map( A => n50, Z => n36);
   U20 : HS65_LH_IVX9 port map( A => n63, Z => n27);
   U21 : HS65_LH_IVX9 port map( A => A(6), Z => n38);
   U22 : HS65_LH_IVX9 port map( A => n69, Z => n30);
   U23 : HS65_LH_OR2X9 port map( A => B(14), B => n21, Z => n49);
   U24 : HS65_LH_IVX9 port map( A => B(12), Z => n7);
   U25 : HS65_LH_IVX9 port map( A => B(13), Z => n8);
   U26 : HS65_LH_IVX9 port map( A => B(15), Z => n9);
   U27 : HS65_LH_IVX9 port map( A => B(7), Z => n4);
   U28 : HS65_LH_IVX9 port map( A => B(5), Z => n3);
   U29 : HS65_LH_IVX9 port map( A => B(9), Z => n5);
   U30 : HS65_LH_IVX9 port map( A => A(1), Z => n41);
   U31 : HS65_LH_IVX9 port map( A => A(4), Z => n40);
   U32 : HS65_LH_IVX9 port map( A => A(10), Z => n35);
   U33 : HS65_LH_OR2X9 port map( A => B(26), B => n22, Z => n65);
   U34 : HS65_LH_IVX9 port map( A => A(16), Z => n33);
   U35 : HS65_LH_IVX9 port map( A => A(24), Z => n28);
   U36 : HS65_LH_IVX9 port map( A => A(18), Z => n31);
   U37 : HS65_LH_IVX9 port map( A => B(23), Z => n14);
   U38 : HS65_LH_IVX9 port map( A => B(19), Z => n11);
   U39 : HS65_LH_IVX9 port map( A => B(25), Z => n15);
   U40 : HS65_LH_IVX9 port map( A => B(21), Z => n13);
   U41 : HS65_LH_IVX9 port map( A => B(17), Z => n10);
   U42 : HS65_LH_IVX9 port map( A => A(30), Z => n25);
   U43 : HS65_LH_IVX9 port map( A => B(29), Z => n18);
   U44 : HS65_LH_CNIVX3 port map( A => EQ_port, Z => NE);
   U45 : HS65_LH_NOR4ABX2 port map( A => n42, B => n43, C => n44, D => n45, Z 
                           => EQ_port);
   U46 : HS65_LH_NAND4X4 port map( A => n46, B => n47, C => n48, D => n49, Z =>
                           n45);
   U47 : HS65_LH_NAND4ABX3 port map( A => n50, B => n34, C => n51, D => n52, Z 
                           => n44);
   U48 : HS65_LH_NOR4ABX2 port map( A => n54, B => n55, C => n56, D => n57, Z 
                           => n43);
   U49 : HS65_LH_NAND4ABX3 port map( A => n58, B => n59, C => n60, D => n61, Z 
                           => n57);
   U50 : HS65_LH_AOI22X1 port map( A => n41, B => n62, C => n62, D => B(1), Z 
                           => n58);
   U51 : HS65_LH_NAND2AX4 port map( A => B(0), B => A(0), Z => n62);
   U52 : HS65_LH_NAND4ABX3 port map( A => n63, B => n26, C => n64, D => n65, Z 
                           => n56);
   U53 : HS65_LH_NOR4ABX2 port map( A => n67, B => n68, C => n69, D => n70, Z 
                           => n55);
   U54 : HS65_LH_AND4X3 port map( A => n71, B => n72, C => n73, D => n74, Z => 
                           n54);
   U55 : HS65_LH_NOR4ABX2 port map( A => n75, B => n76, C => n77, D => LT_port,
                           Z => n42);
   U56 : HS65_LH_OAI22X1 port map( A => A(31), B => n19, C => n23, D => n78, Z 
                           => LT_port);
   U57 : HS65_LH_AOI32X3 port map( A => n61, B => n24, C => n79, D => B(30), E 
                           => n25, Z => n78);
   U58 : HS65_LH_OAI212X3 port map( A => A(28), B => n17, C => A(29), D => n18,
                           E => n80, Z => n79);
   U59 : HS65_LH_NAND3X2 port map( A => n60, B => n66, C => n81, Z => n80);
   U60 : HS65_LH_OAI12X2 port map( A => A(27), B => n16, C => n82, Z => n81);
   U61 : HS65_LH_AOI32X3 port map( A => n65, B => n64, C => n83, D => B(26), E 
                           => n22, Z => n82);
   U62 : HS65_LH_OAI12X2 port map( A => A(25), B => n15, C => n84, Z => n83);
   U63 : HS65_LH_AOI32X3 port map( A => n27, B => n71, C => n85, D => B(24), E 
                           => n28, Z => n84);
   U64 : HS65_LH_OAI12X2 port map( A => A(23), B => n14, C => n86, Z => n85);
   U65 : HS65_LH_AOI32X3 port map( A => n72, B => n74, C => n87, D => B(22), E 
                           => n29, Z => n86);
   U66 : HS65_LH_OAI212X3 port map( A => A(20), B => n12, C => A(21), D => n13,
                           E => n88, Z => n87);
   U67 : HS65_LH_NAND3X2 port map( A => n73, B => n67, C => n89, Z => n88);
   U68 : HS65_LH_OAI12X2 port map( A => A(19), B => n11, C => n90, Z => n89);
   U69 : HS65_LH_AOI32X3 port map( A => n30, B => n68, C => n91, D => B(18), E 
                           => n31, Z => n90);
   U70 : HS65_LH_OAI12X2 port map( A => A(17), B => n10, C => n92, Z => n91);
   U71 : HS65_LH_AOI32X3 port map( A => n32, B => n48, C => n93, D => B(16), E 
                           => n33, Z => n92);
   U72 : HS65_LH_OAI12X2 port map( A => A(15), B => n9, C => n94, Z => n93);
   U73 : HS65_LH_AOI32X3 port map( A => n49, B => n47, C => n95, D => B(14), E 
                           => n21, Z => n94);
   U74 : HS65_LH_OAI212X3 port map( A => A(12), B => n7, C => A(13), D => n8, E
                           => n96, Z => n95);
   U75 : HS65_LH_NAND3X2 port map( A => n46, B => n53, C => n97, Z => n96);
   U76 : HS65_LH_OAI12X2 port map( A => A(11), B => n6, C => n98, Z => n97);
   U77 : HS65_LH_AOI32X3 port map( A => n52, B => n51, C => n99, D => B(10), E 
                           => n35, Z => n98);
   U78 : HS65_LH_OAI12X2 port map( A => A(9), B => n5, C => n100, Z => n99);
   U79 : HS65_LH_AOI32X3 port map( A => n36, B => n101, C => n102, D => B(8), E
                           => n20, Z => n100);
   U80 : HS65_LH_OAI12X2 port map( A => A(7), B => n4, C => n103, Z => n102);
   U81 : HS65_LH_AOI32X3 port map( A => n104, B => n105, C => n106, D => B(6), 
                           E => n38, Z => n103);
   U82 : HS65_LH_OAI12X2 port map( A => A(5), B => n3, C => n107, Z => n106);
   U83 : HS65_LH_AOI32X3 port map( A => n39, B => n108, C => n109, D => B(4), E
                           => n40, Z => n107);
   U84 : HS65_LH_OAI212X3 port map( A => A(2), B => n1, C => A(3), D => n2, E 
                           => n110, Z => n109);
   U85 : HS65_LH_OAI212X3 port map( A => B(1), B => n111, C => n112, D => n41, 
                           E => n113, Z => n110);
   U86 : HS65_LH_AND2X4 port map( A => n112, B => n41, Z => n111);
   U87 : HS65_LH_NOR2AX3 port map( A => B(0), B => A(0), Z => n112);
   U88 : HS65_LH_NOR2X2 port map( A => n20, B => B(8), Z => n50);
   U89 : HS65_LH_NAND2X2 port map( A => A(9), B => n5, Z => n51);
   U90 : HS65_LH_NAND2AX4 port map( A => B(10), B => A(10), Z => n52);
   U91 : HS65_LH_NAND2X2 port map( A => A(11), B => n6, Z => n53);
   U92 : HS65_LH_NAND2X2 port map( A => A(12), B => n7, Z => n46);
   U93 : HS65_LH_NAND2X2 port map( A => A(13), B => n8, Z => n47);
   U94 : HS65_LH_NAND2X2 port map( A => A(15), B => n9, Z => n48);
   U95 : HS65_LH_NOR2X2 port map( A => n33, B => B(16), Z => n70);
   U96 : HS65_LH_NAND2X2 port map( A => A(17), B => n10, Z => n68);
   U97 : HS65_LH_NOR2X2 port map( A => B(18), B => n31, Z => n69);
   U98 : HS65_LH_NAND2X2 port map( A => A(19), B => n11, Z => n67);
   U99 : HS65_LH_NAND2X2 port map( A => A(20), B => n12, Z => n73);
   U100 : HS65_LH_NAND2X2 port map( A => A(21), B => n13, Z => n74);
   U101 : HS65_LH_NAND2AX4 port map( A => B(22), B => A(22), Z => n72);
   U102 : HS65_LH_NAND2X2 port map( A => A(23), B => n14, Z => n71);
   U103 : HS65_LH_NOR2X2 port map( A => n28, B => B(24), Z => n63);
   U104 : HS65_LH_NAND2X2 port map( A => A(25), B => n15, Z => n64);
   U105 : HS65_LH_NAND2X2 port map( A => A(27), B => n16, Z => n66);
   U106 : HS65_LH_NAND2X2 port map( A => A(28), B => n17, Z => n60);
   U107 : HS65_LH_NOR2X2 port map( A => n25, B => B(30), Z => n59);
   U108 : HS65_LH_NAND2X2 port map( A => A(29), B => n18, Z => n61);
   U109 : HS65_LH_NAND4ABX3 port map( A => n114, B => n37, C => n105, D => n104
                           , Z => n77);
   U110 : HS65_LH_NAND2AX4 port map( A => B(6), B => A(6), Z => n104);
   U111 : HS65_LH_NAND2X2 port map( A => A(5), B => n3, Z => n105);
   U112 : HS65_LH_NAND2X2 port map( A => A(7), B => n4, Z => n101);
   U113 : HS65_LH_NOR2X2 port map( A => n40, B => B(4), Z => n114);
   U114 : HS65_LH_AND2X4 port map( A => n113, B => n108, Z => n76);
   U115 : HS65_LH_NAND2X2 port map( A => A(3), B => n2, Z => n108);
   U116 : HS65_LH_NAND2X2 port map( A => A(2), B => n1, Z => n113);
   U117 : HS65_LH_NAND2X2 port map( A => A(31), B => n19, Z => n75);

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end alu_DW01_sub_0;

architecture SYN_rpl of alu_DW01_sub_0 is

   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33 : 
      std_logic;

begin
   
   U2_23 : HS65_LH_FA1X4 port map( A0 => A(23), B0 => n25, CI => carry_23_port,
                           CO => carry_24_port, S0 => DIFF(23));
   U2_29 : HS65_LH_FA1X4 port map( A0 => A(29), B0 => n31, CI => carry_29_port,
                           CO => carry_30_port, S0 => DIFF(29));
   U2_26 : HS65_LH_FA1X4 port map( A0 => A(26), B0 => n28, CI => carry_26_port,
                           CO => carry_27_port, S0 => DIFF(26));
   U2_17 : HS65_LH_FA1X4 port map( A0 => A(17), B0 => n19, CI => carry_17_port,
                           CO => carry_18_port, S0 => DIFF(17));
   U2_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => n7, CI => carry_5_port, CO 
                           => carry_6_port, S0 => DIFF(5));
   U2_14 : HS65_LH_FA1X4 port map( A0 => A(14), B0 => n16, CI => carry_14_port,
                           CO => carry_15_port, S0 => DIFF(14));
   U2_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => n10, CI => carry_8_port, CO
                           => carry_9_port, S0 => DIFF(8));
   U2_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => n5, CI => carry_3_port, CO 
                           => carry_4_port, S0 => DIFF(3));
   U2_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => n3, CI => carry_1_port, CO 
                           => carry_2_port, S0 => DIFF(1));
   U2_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => n11, CI => carry_9_port, CO
                           => carry_10_port, S0 => DIFF(9));
   U2_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => n9, CI => carry_7_port, CO 
                           => carry_8_port, S0 => DIFF(7));
   U2_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => n12, CI => carry_10_port,
                           CO => carry_11_port, S0 => DIFF(10));
   U2_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => n8, CI => carry_6_port, CO 
                           => carry_7_port, S0 => DIFF(6));
   U2_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => n6, CI => carry_4_port, CO 
                           => carry_5_port, S0 => DIFF(4));
   U2_30 : HS65_LH_FA1X4 port map( A0 => A(30), B0 => n32, CI => carry_30_port,
                           CO => carry_31_port, S0 => DIFF(30));
   U2_25 : HS65_LH_FA1X4 port map( A0 => A(25), B0 => n27, CI => carry_25_port,
                           CO => carry_26_port, S0 => DIFF(25));
   U2_19 : HS65_LH_FA1X4 port map( A0 => A(19), B0 => n21, CI => carry_19_port,
                           CO => carry_20_port, S0 => DIFF(19));
   U2_27 : HS65_LH_FA1X4 port map( A0 => A(27), B0 => n29, CI => carry_27_port,
                           CO => carry_28_port, S0 => DIFF(27));
   U2_24 : HS65_LH_FA1X4 port map( A0 => A(24), B0 => n26, CI => carry_24_port,
                           CO => carry_25_port, S0 => DIFF(24));
   U2_21 : HS65_LH_FA1X4 port map( A0 => A(21), B0 => n23, CI => carry_21_port,
                           CO => carry_22_port, S0 => DIFF(21));
   U2_18 : HS65_LH_FA1X4 port map( A0 => A(18), B0 => n20, CI => carry_18_port,
                           CO => carry_19_port, S0 => DIFF(18));
   U2_13 : HS65_LH_FA1X4 port map( A0 => A(13), B0 => n15, CI => carry_13_port,
                           CO => carry_14_port, S0 => DIFF(13));
   U2_12 : HS65_LH_FA1X4 port map( A0 => A(12), B0 => n14, CI => carry_12_port,
                           CO => carry_13_port, S0 => DIFF(12));
   U2_22 : HS65_LH_FA1X4 port map( A0 => A(22), B0 => n24, CI => carry_22_port,
                           CO => carry_23_port, S0 => DIFF(22));
   U2_15 : HS65_LH_FA1X4 port map( A0 => A(15), B0 => n17, CI => carry_15_port,
                           CO => carry_16_port, S0 => DIFF(15));
   U2_28 : HS65_LH_FA1X4 port map( A0 => A(28), B0 => n30, CI => carry_28_port,
                           CO => carry_29_port, S0 => DIFF(28));
   U2_16 : HS65_LH_FA1X4 port map( A0 => A(16), B0 => n18, CI => carry_16_port,
                           CO => carry_17_port, S0 => DIFF(16));
   U2_31 : HS65_LHS_XOR3X2 port map( A => A(31), B => n33, C => carry_31_port, 
                           Z => DIFF(31));
   U2_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => n4, CI => carry_2_port, CO 
                           => carry_3_port, S0 => DIFF(2));
   U2_20 : HS65_LH_FA1X4 port map( A0 => A(20), B0 => n22, CI => carry_20_port,
                           CO => carry_21_port, S0 => DIFF(20));
   U2_11 : HS65_LH_FA1X4 port map( A0 => A(11), B0 => n13, CI => carry_11_port,
                           CO => carry_12_port, S0 => DIFF(11));
   U1 : HS65_LH_IVX9 port map( A => B(11), Z => n13);
   U2 : HS65_LH_IVX9 port map( A => B(20), Z => n22);
   U3 : HS65_LH_IVX9 port map( A => B(2), Z => n4);
   U4 : HS65_LH_IVX9 port map( A => B(31), Z => n33);
   U5 : HS65_LH_IVX9 port map( A => B(16), Z => n18);
   U6 : HS65_LH_IVX9 port map( A => B(28), Z => n30);
   U7 : HS65_LH_IVX9 port map( A => B(15), Z => n17);
   U8 : HS65_LH_IVX9 port map( A => B(22), Z => n24);
   U9 : HS65_LH_IVX9 port map( A => B(12), Z => n14);
   U10 : HS65_LH_IVX9 port map( A => B(13), Z => n15);
   U11 : HS65_LH_IVX9 port map( A => B(18), Z => n20);
   U12 : HS65_LH_IVX9 port map( A => B(21), Z => n23);
   U13 : HS65_LH_IVX9 port map( A => B(24), Z => n26);
   U14 : HS65_LH_IVX9 port map( A => B(27), Z => n29);
   U15 : HS65_LH_IVX9 port map( A => B(19), Z => n21);
   U16 : HS65_LH_IVX9 port map( A => B(25), Z => n27);
   U17 : HS65_LH_IVX9 port map( A => B(30), Z => n32);
   U18 : HS65_LH_IVX9 port map( A => B(4), Z => n6);
   U19 : HS65_LH_IVX9 port map( A => B(6), Z => n8);
   U20 : HS65_LH_IVX9 port map( A => B(10), Z => n12);
   U21 : HS65_LH_IVX9 port map( A => B(7), Z => n9);
   U22 : HS65_LH_IVX9 port map( A => B(9), Z => n11);
   U23 : HS65_LH_IVX9 port map( A => B(1), Z => n3);
   U24 : HS65_LH_NAND2X7 port map( A => n1, B => B(0), Z => carry_1_port);
   U25 : HS65_LH_IVX9 port map( A => B(3), Z => n5);
   U26 : HS65_LH_IVX9 port map( A => B(8), Z => n10);
   U27 : HS65_LH_IVX9 port map( A => B(14), Z => n16);
   U28 : HS65_LH_IVX9 port map( A => B(5), Z => n7);
   U29 : HS65_LH_IVX9 port map( A => B(17), Z => n19);
   U30 : HS65_LH_IVX9 port map( A => B(26), Z => n28);
   U31 : HS65_LH_IVX9 port map( A => B(29), Z => n31);
   U32 : HS65_LH_IVX9 port map( A => B(23), Z => n25);
   U33 : HS65_LH_IVX9 port map( A => A(0), Z => n1);
   U34 : HS65_LH_IVX9 port map( A => B(0), Z => n2);
   U35 : HS65_LHS_XNOR2X6 port map( A => A(0), B => n2, Z => DIFF(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_DW_cmp_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in 
         std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);

end alu_DW_cmp_0;

architecture SYN_USE_DEFA_ARCH_NAME of alu_DW_cmp_0 is

   component HS65_LH_NAND2AX4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI312X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI112X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X3
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA32X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X1
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X2
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3AX3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X1
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA12X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA112X4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI32X2
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328 : std_logic;

begin
   
   U157 : HS65_LH_IVX9 port map( A => n296, Z => n247);
   U158 : HS65_LH_IVX9 port map( A => n305, Z => n256);
   U159 : HS65_LH_IVX9 port map( A => n306, Z => n260);
   U160 : HS65_LH_OR2X9 port map( A => B(11), B => n241, Z => n327);
   U161 : HS65_LH_IVX9 port map( A => n279, Z => n252);
   U162 : HS65_LH_IVX9 port map( A => n297, Z => n246);
   U163 : HS65_LH_IVX9 port map( A => n284, Z => n250);
   U164 : HS65_LH_IVX9 port map( A => n308, Z => n263);
   U165 : HS65_LH_IVX9 port map( A => B(3), Z => n228);
   U166 : HS65_LH_IVX9 port map( A => B(4), Z => n229);
   U167 : HS65_LH_IVX9 port map( A => A(11), Z => n241);
   U168 : HS65_LH_IVX9 port map( A => A(17), Z => n243);
   U169 : HS65_LH_IVX9 port map( A => B(27), Z => n237);
   U170 : HS65_LH_IVX9 port map( A => B(2), Z => n227);
   U171 : HS65_LH_IVX9 port map( A => A(8), Z => n240);
   U172 : HS65_LH_IVX9 port map( A => A(14), Z => n242);
   U173 : HS65_LH_IVX9 port map( A => A(5), Z => n239);
   U174 : HS65_LH_IVX9 port map( A => A(20), Z => n244);
   U175 : HS65_LH_IVX9 port map( A => A(29), Z => n245);
   U176 : HS65_LH_IVX9 port map( A => n321, Z => n257);
   U177 : HS65_LH_IVX9 port map( A => A(15), Z => n255);
   U178 : HS65_LH_IVX9 port map( A => A(7), Z => n264);
   U179 : HS65_LH_IVX9 port map( A => A(4), Z => n267);
   U180 : HS65_LH_IVX9 port map( A => n316, Z => n266);
   U181 : HS65_LH_IVX9 port map( A => B(25), Z => n235);
   U182 : HS65_LH_IVX9 port map( A => A(1), Z => n268);
   U183 : HS65_LH_IVX9 port map( A => n320, Z => n254);
   U184 : HS65_LH_AND2X4 port map( A => A(3), B => n228, Z => n318);
   U185 : HS65_LH_OR2X9 port map( A => B(17), B => n243, Z => n281);
   U186 : HS65_LH_IVX9 port map( A => A(9), Z => n262);
   U187 : HS65_LH_IVX9 port map( A => A(31), Z => n248);
   U188 : HS65_LH_IVX9 port map( A => A(16), Z => n253);
   U189 : HS65_LH_IVX9 port map( A => A(28), Z => n249);
   U190 : HS65_LH_IVX9 port map( A => A(21), Z => n251);
   U191 : HS65_LH_IVX9 port map( A => A(13), Z => n258);
   U192 : HS65_LH_IVX9 port map( A => A(12), Z => n259);
   U193 : HS65_LH_IVX9 port map( A => B(1), Z => n226);
   U194 : HS65_LH_IVX9 port map( A => B(23), Z => n233);
   U195 : HS65_LH_IVX9 port map( A => B(19), Z => n231);
   U196 : HS65_LH_IVX9 port map( A => B(26), Z => n236);
   U197 : HS65_LH_IVX9 port map( A => B(22), Z => n232);
   U198 : HS65_LH_IVX9 port map( A => B(18), Z => n230);
   U199 : HS65_LH_IVX9 port map( A => B(24), Z => n234);
   U200 : HS65_LH_IVX9 port map( A => B(30), Z => n238);
   U201 : HS65_LH_IVX9 port map( A => A(6), Z => n265);
   U202 : HS65_LH_IVX9 port map( A => A(10), Z => n261);
   U203 : HS65_LH_OAI12X2 port map( A => n269, B => n270, C => n271, Z => 
                           GE_LT_GT_LE);
   U204 : HS65_LH_OAI32X2 port map( A => n272, B => n273, C => n274, D => n275,
                           E => n272, Z => n271);
   U205 : HS65_LH_AOI212X2 port map( A => n276, B => n277, C => n277, D => n252
                           , E => n278, Z => n274);
   U206 : HS65_LH_OA32X4 port map( A => n230, B => A(18), C => n280, D => A(19)
                           , E => n231, Z => n277);
   U207 : HS65_LH_AOI32X3 port map( A => n281, B => n253, C => B(16), D => 
                           B(17), E => n243, Z => n276);
   U208 : HS65_LH_AOI22X1 port map( A => n282, B => n283, C => n283, D => n250,
                           Z => n273);
   U209 : HS65_LH_OA32X4 port map( A => n232, B => A(22), C => n285, D => A(23)
                           , E => n233, Z => n283);
   U210 : HS65_LH_AOI32X3 port map( A => n286, B => n244, C => B(20), D => 
                           B(21), E => n251, Z => n282);
   U211 : HS65_LH_CBI4I1X3 port map( A => n247, B => n246, C => n287, D => n288
                           , Z => n272);
   U212 : HS65_LH_OAI212X3 port map( A => n289, B => n290, C => n291, D => n289
                           , E => n292, Z => n288);
   U213 : HS65_LH_OAI32X2 port map( A => n234, B => A(24), C => n293, D => 
                           A(25), E => n235, Z => n290);
   U214 : HS65_LH_OAI32X2 port map( A => n236, B => A(26), C => n294, D => 
                           A(27), E => n237, Z => n289);
   U215 : HS65_LH_AOI312X2 port map( A => n295, B => n249, C => B(28), D => 
                           B(29), E => n245, F => n296, Z => n287);
   U216 : HS65_LH_OAI32X2 port map( A => n238, B => A(30), C => n298, D => 
                           B(31), E => n248, Z => n296);
   U217 : HS65_LH_NAND3AX3 port map( A => n278, B => n279, C => n275, Z => n270
                           );
   U218 : HS65_LH_AND3X4 port map( A => n291, B => n292, C => n299, Z => n275);
   U219 : HS65_LH_AOI12X2 port map( A => A(24), B => n234, C => n293, Z => n299
                           );
   U220 : HS65_LH_NOR2AX3 port map( A => A(25), B => B(25), Z => n293);
   U221 : HS65_LH_OA112X4 port map( A => B(28), B => n249, C => n295, D => n297
                           , Z => n292);
   U222 : HS65_LH_AOI12X2 port map( A => n238, B => A(30), C => n298, Z => n297
                           );
   U223 : HS65_LH_AND2X4 port map( A => B(31), B => n248, Z => n298);
   U224 : HS65_LH_OR2X4 port map( A => B(29), B => n245, Z => n295);
   U225 : HS65_LH_AOI12X2 port map( A => n236, B => A(26), C => n294, Z => n291
                           );
   U226 : HS65_LH_AND2X4 port map( A => A(27), B => n237, Z => n294);
   U227 : HS65_LH_AOI12X2 port map( A => n230, B => A(18), C => n280, Z => n279
                           );
   U228 : HS65_LH_AND2X4 port map( A => A(19), B => n231, Z => n280);
   U229 : HS65_LH_OAI112X1 port map( A => B(20), B => n244, C => n286, D => 
                           n284, Z => n278);
   U230 : HS65_LH_AOI12X2 port map( A => n232, B => A(22), C => n285, Z => n284
                           );
   U231 : HS65_LH_AND2X4 port map( A => A(23), B => n233, Z => n285);
   U232 : HS65_LH_OR2X4 port map( A => B(21), B => n251, Z => n286);
   U233 : HS65_LH_OAI212X3 port map( A => n300, B => n301, C => n302, D => n300
                           , E => n303, Z => n269);
   U234 : HS65_LH_OA12X4 port map( A => n253, B => B(16), C => n281, Z => n303)
                           ;
   U235 : HS65_LH_NOR3X1 port map( A => n304, B => n305, C => n306, Z => n302);
   U236 : HS65_LH_OAI12X2 port map( A => B(8), B => n240, C => n307, Z => n304)
                           ;
   U237 : HS65_LH_CBI4I1X3 port map( A => n308, B => n309, C => n310, D => n311
                           , Z => n301);
   U238 : HS65_LH_NAND3AX3 port map( A => n309, B => n312, C => n313, Z => n311
                           );
   U239 : HS65_LH_AOI212X2 port map( A => n314, B => n315, C => A(4), D => n229
                           , E => n316, Z => n313);
   U240 : HS65_LH_AOI22X1 port map( A => B(1), B => n268, C => n317, D => B(0),
                           Z => n314);
   U241 : HS65_LH_AOI12X2 port map( A => A(1), B => n226, C => A(0), Z => n317)
                           ;
   U242 : HS65_LH_CBI4I1X3 port map( A => A(2), B => n227, C => n318, D => n315
                           , Z => n312);
   U243 : HS65_LH_OA32X4 port map( A => n227, B => A(2), C => n318, D => A(3), 
                           E => n228, Z => n315);
   U244 : HS65_LH_AOI312X2 port map( A => n266, B => n267, C => B(4), D => B(5)
                           , E => n239, F => n263, Z => n310);
   U245 : HS65_LH_NOR2X2 port map( A => n239, B => B(5), Z => n316);
   U246 : HS65_LH_OAI12X2 port map( A => B(6), B => n265, C => n319, Z => n309)
                           ;
   U247 : HS65_LH_AOI32X3 port map( A => B(6), B => n265, C => n319, D => n264,
                           E => B(7), Z => n308);
   U248 : HS65_LH_NAND2AX4 port map( A => B(7), B => A(7), Z => n319);
   U249 : HS65_LH_CBI4I1X3 port map( A => n320, B => n321, C => n322, D => n323
                           , Z => n300);
   U250 : HS65_LH_OAI212X3 port map( A => n324, B => n325, C => n260, D => n324
                           , E => n256, Z => n323);
   U251 : HS65_LH_OAI112X1 port map( A => B(12), B => n259, C => n326, D => 
                           n257, Z => n305);
   U252 : HS65_LH_OAI12X2 port map( A => B(10), B => n261, C => n327, Z => n306
                           );
   U253 : HS65_LH_AO32X4 port map( A => B(8), B => n240, C => n307, D => n262, 
                           E => B(9), Z => n325);
   U254 : HS65_LH_NAND2AX4 port map( A => B(9), B => A(9), Z => n307);
   U255 : HS65_LH_AO32X4 port map( A => B(10), B => n261, C => n327, D => n241,
                           E => B(11), Z => n324);
   U256 : HS65_LH_AOI312X2 port map( A => n326, B => n259, C => B(12), D => 
                           B(13), E => n258, F => n254, Z => n322);
   U257 : HS65_LH_OR2X4 port map( A => B(13), B => n258, Z => n326);
   U258 : HS65_LH_OAI12X2 port map( A => B(14), B => n242, C => n328, Z => n321
                           );
   U259 : HS65_LH_AOI32X3 port map( A => B(14), B => n242, C => n328, D => n255
                           , E => B(15), Z => n320);
   U260 : HS65_LH_NAND2AX4 port map( A => B(15), B => A(15), Z => n328);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity exe_top_DW01_add_0 is

   port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (11 downto 0);  CO : out std_logic);

end exe_top_DW01_add_0;

architecture SYN_rpl of exe_top_DW01_add_0 is

   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR3X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_FA1X4
      port( A0, B0, CI : in std_logic;  CO, S0 : out std_logic);
   end component;
   
   signal carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1 : std_logic;

begin
   
   U1_1 : HS65_LH_FA1X4 port map( A0 => A(1), B0 => B(1), CI => n1, CO => 
                           carry_2_port, S0 => SUM(1));
   U1_10 : HS65_LH_FA1X4 port map( A0 => A(10), B0 => B(10), CI => 
                           carry_10_port, CO => carry_11_port, S0 => SUM(10));
   U1_9 : HS65_LH_FA1X4 port map( A0 => A(9), B0 => B(9), CI => carry_9_port, 
                           CO => carry_10_port, S0 => SUM(9));
   U1_8 : HS65_LH_FA1X4 port map( A0 => A(8), B0 => B(8), CI => carry_8_port, 
                           CO => carry_9_port, S0 => SUM(8));
   U1_7 : HS65_LH_FA1X4 port map( A0 => A(7), B0 => B(7), CI => carry_7_port, 
                           CO => carry_8_port, S0 => SUM(7));
   U1_6 : HS65_LH_FA1X4 port map( A0 => A(6), B0 => B(6), CI => carry_6_port, 
                           CO => carry_7_port, S0 => SUM(6));
   U1_5 : HS65_LH_FA1X4 port map( A0 => A(5), B0 => B(5), CI => carry_5_port, 
                           CO => carry_6_port, S0 => SUM(5));
   U1_4 : HS65_LH_FA1X4 port map( A0 => A(4), B0 => B(4), CI => carry_4_port, 
                           CO => carry_5_port, S0 => SUM(4));
   U1_3 : HS65_LH_FA1X4 port map( A0 => A(3), B0 => B(3), CI => carry_3_port, 
                           CO => carry_4_port, S0 => SUM(3));
   U1_2 : HS65_LH_FA1X4 port map( A0 => A(2), B0 => B(2), CI => carry_2_port, 
                           CO => carry_3_port, S0 => SUM(2));
   U1_11 : HS65_LHS_XOR3X2 port map( A => A(11), B => B(11), C => carry_11_port
                           , Z => SUM(11));
   U1 : HS65_LH_AND2X4 port map( A => A(0), B => B(0), Z => n1);
   U2 : HS65_LHS_XOR2X6 port map( A => A(0), B => B(0), Z => SUM(0));

end SYN_rpl;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu_ctrl is

   port( alu_ctrl_i : in std_logic_vector (9 downto 0);  alu_ctrl_o : out 
         std_logic_vector (6 downto 0));

end alu_ctrl;

architecture SYN_Behavioral of alu_ctrl is

   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI312X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI13X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I6X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI211X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI311X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI33X3
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO312X9
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   signal n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17 : std_logic;

begin
   
   U3 : HS65_LH_AOI12X2 port map( A => n38, B => n39, C => alu_ctrl_i(9), Z => 
                           alu_ctrl_o(2));
   U4 : HS65_LH_OAI32X5 port map( A => n41, B => alu_ctrl_i(9), C => 
                           alu_ctrl_i(7), D => n17, E => n28, Z => 
                           alu_ctrl_o(1));
   U5 : HS65_LH_IVX9 port map( A => n30, Z => n13);
   U6 : HS65_LH_NAND3X5 port map( A => n16, B => n14, C => n17, Z => n30);
   U7 : HS65_LH_AO312X9 port map( A => n11, B => n7, C => n1, D => n25, E => 
                           n12, F => n23, Z => alu_ctrl_o(4));
   U8 : HS65_LH_OAI33X3 port map( A => n29, B => n9, C => n30, D => n14, E => 
                           n17, F => n16, Z => n25);
   U9 : HS65_LH_IVX9 port map( A => n31, Z => n9);
   U10 : HS65_LH_NAND2X7 port map( A => n13, B => n12, Z => n20);
   U11 : HS65_LH_IVX9 port map( A => n35, Z => n5);
   U12 : HS65_LH_IVX9 port map( A => n27, Z => n1);
   U13 : HS65_LH_IVX9 port map( A => n41, Z => n15);
   U14 : HS65_LH_NOR2AX3 port map( A => n19, B => n20, Z => alu_ctrl_o(0));
   U15 : HS65_LH_AOI311X4 port map( A => alu_ctrl_i(0), B => n8, C => n40, D =>
                           n3, E => n15, Z => n39);
   U16 : HS65_LH_AOI12X2 port map( A => alu_ctrl_i(7), B => n17, C => n44, Z =>
                           n38);
   U17 : HS65_LH_IVX9 port map( A => n33, Z => n3);
   U18 : HS65_LH_OAI32X5 port map( A => n26, B => n7, C => n27, D => 
                           alu_ctrl_i(6), E => n28, Z => n23);
   U19 : HS65_LH_NAND2X7 port map( A => alu_ctrl_i(1), B => n11, Z => n26);
   U20 : HS65_LH_OAI211X5 port map( A => n20, B => n4, C => n2, D => n21, Z => 
                           alu_ctrl_o(5));
   U21 : HS65_LH_IVX9 port map( A => n24, Z => n4);
   U22 : HS65_LH_AOI32X5 port map( A => n1, B => alu_ctrl_i(0), C => n22, D => 
                           n5, E => n12, Z => n21);
   U23 : HS65_LH_IVX9 port map( A => n23, Z => n2);
   U24 : HS65_LH_NOR3AX2 port map( A => n45, B => n30, C => n6, Z => n40);
   U25 : HS65_LH_NOR3X4 port map( A => n10, B => alu_ctrl_i(4), C => 
                           alu_ctrl_i(2), Z => n45);
   U26 : HS65_LH_IVX9 port map( A => alu_ctrl_i(0), Z => n11);
   U27 : HS65_LH_AOI32X5 port map( A => alu_ctrl_i(4), B => alu_ctrl_i(0), C =>
                           alu_ctrl_i(3), D => n11, E => n7, Z => n37);
   U28 : HS65_LH_NOR3X4 port map( A => n7, B => alu_ctrl_i(1), C => n43, Z => 
                           n24);
   U29 : HS65_LHS_XNOR2X6 port map( A => alu_ctrl_i(0), B => n10, Z => n31);
   U30 : HS65_LH_CBI4I6X5 port map( A => n30, B => n29, C => n35, D => 
                           alu_ctrl_i(0), Z => n44);
   U31 : HS65_LH_IVX9 port map( A => alu_ctrl_i(6), Z => n17);
   U32 : HS65_LH_IVX9 port map( A => alu_ctrl_i(1), Z => n10);
   U33 : HS65_LH_IVX9 port map( A => alu_ctrl_i(4), Z => n7);
   U34 : HS65_LH_OAI21X3 port map( A => n42, B => n24, C => n13, Z => n33);
   U35 : HS65_LH_NOR3X4 port map( A => n43, B => alu_ctrl_i(4), C => n10, Z => 
                           n42);
   U36 : HS65_LH_IVX9 port map( A => alu_ctrl_i(9), Z => n12);
   U37 : HS65_LH_IVX9 port map( A => alu_ctrl_i(7), Z => n16);
   U38 : HS65_LH_NAND4ABX3 port map( A => alu_ctrl_i(3), B => alu_ctrl_i(2), C 
                           => n6, D => n11, Z => n43);
   U39 : HS65_LH_NAND4ABX3 port map( A => alu_ctrl_i(2), B => n20, C => n8, D 
                           => n6, Z => n27);
   U40 : HS65_LH_NAND2X7 port map( A => n40, B => alu_ctrl_i(3), Z => n35);
   U41 : HS65_LH_IVX9 port map( A => alu_ctrl_i(8), Z => n14);
   U42 : HS65_LH_AOI13X5 port map( A => n32, B => n33, C => n34, D => 
                           alu_ctrl_i(9), Z => alu_ctrl_o(3));
   U43 : HS65_LH_AOI22X6 port map( A => n5, B => alu_ctrl_i(0), C => n15, D => 
                           alu_ctrl_i(7), Z => n34);
   U44 : HS65_LH_NAND3X5 port map( A => n36, B => n10, C => n13, Z => n32);
   U45 : HS65_LH_OAI32X5 port map( A => n37, B => alu_ctrl_i(5), C => 
                           alu_ctrl_i(2), D => alu_ctrl_i(0), E => n29, Z => 
                           n36);
   U46 : HS65_LH_NOR2X6 port map( A => alu_ctrl_i(9), B => n18, Z => 
                           alu_ctrl_o(6));
   U47 : HS65_LH_AOI312X4 port map( A => n17, B => n16, C => n19, D => 
                           alu_ctrl_i(7), E => alu_ctrl_i(6), F => n15, Z => 
                           n18);
   U48 : HS65_LH_NAND4ABX3 port map( A => alu_ctrl_i(4), B => alu_ctrl_i(3), C 
                           => alu_ctrl_i(5), D => alu_ctrl_i(2), Z => n29);
   U49 : HS65_LH_NAND3X5 port map( A => n14, B => n12, C => alu_ctrl_i(7), Z =>
                           n28);
   U50 : HS65_LH_NOR4ABX2 port map( A => n11, B => n46, C => n8, D => n31, Z =>
                           n19);
   U51 : HS65_LH_NOR3X4 port map( A => alu_ctrl_i(2), B => alu_ctrl_i(5), C => 
                           alu_ctrl_i(4), Z => n46);
   U52 : HS65_LH_IVX9 port map( A => alu_ctrl_i(3), Z => n8);
   U53 : HS65_LH_NOR2X6 port map( A => alu_ctrl_i(4), B => n10, Z => n22);
   U54 : HS65_LH_IVX9 port map( A => alu_ctrl_i(5), Z => n6);
   U55 : HS65_LH_NAND2X7 port map( A => alu_ctrl_i(8), B => n17, Z => n41);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity alu is

   port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 0);
         alu_o : out std_logic_vector (32 downto 0));

end alu;

architecture SYN_behavioral of alu is

   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR2X9
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI222X2
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI212X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO12X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I6X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI12X2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI211X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI32X5
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO112X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component alu_DW_mult_uns_0
      port( a, b : in std_logic_vector (31 downto 0);  product : out 
            std_logic_vector (63 downto 0));
   end component;
   
   component alu_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component alu_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component alu_DW_cmp_0
      port( A, B : in std_logic_vector (31 downto 0);  TC, GE_LT, GE_GT_EQ : in
            std_logic;  GE_LT_GT_LE, EQ_NE : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal HI_LO_c_HI_31_port, HI_LO_c_HI_30_port, HI_LO_c_HI_29_port, 
      HI_LO_c_HI_28_port, HI_LO_c_HI_27_port, HI_LO_c_HI_26_port, 
      HI_LO_c_HI_25_port, HI_LO_c_HI_24_port, HI_LO_c_HI_23_port, 
      HI_LO_c_HI_22_port, HI_LO_c_HI_21_port, HI_LO_c_HI_20_port, 
      HI_LO_c_HI_19_port, HI_LO_c_HI_18_port, HI_LO_c_HI_17_port, 
      HI_LO_c_HI_16_port, HI_LO_c_HI_15_port, HI_LO_c_HI_14_port, 
      HI_LO_c_HI_13_port, HI_LO_c_HI_12_port, HI_LO_c_HI_11_port, 
      HI_LO_c_HI_10_port, HI_LO_c_HI_9_port, HI_LO_c_HI_8_port, 
      HI_LO_c_HI_7_port, HI_LO_c_HI_6_port, HI_LO_c_HI_5_port, 
      HI_LO_c_HI_4_port, HI_LO_c_HI_3_port, HI_LO_c_HI_2_port, 
      HI_LO_c_HI_1_port, HI_LO_c_HI_0_port, HI_LO_c_LO_31_port, 
      HI_LO_c_LO_30_port, HI_LO_c_LO_29_port, HI_LO_c_LO_28_port, 
      HI_LO_c_LO_27_port, HI_LO_c_LO_26_port, HI_LO_c_LO_25_port, 
      HI_LO_c_LO_24_port, HI_LO_c_LO_23_port, HI_LO_c_LO_22_port, 
      HI_LO_c_LO_21_port, HI_LO_c_LO_20_port, HI_LO_c_LO_19_port, 
      HI_LO_c_LO_18_port, HI_LO_c_LO_17_port, HI_LO_c_LO_16_port, 
      HI_LO_c_LO_15_port, HI_LO_c_LO_14_port, HI_LO_c_LO_13_port, 
      HI_LO_c_LO_12_port, HI_LO_c_LO_11_port, HI_LO_c_LO_10_port, 
      HI_LO_c_LO_9_port, HI_LO_c_LO_8_port, HI_LO_c_LO_7_port, 
      HI_LO_c_LO_6_port, HI_LO_c_LO_5_port, HI_LO_c_LO_4_port, 
      HI_LO_c_LO_3_port, HI_LO_c_LO_2_port, HI_LO_c_LO_1_port, 
      HI_LO_c_LO_0_port, N99, N100, N101, N102, N103, N104, N105, N106, N107, 
      N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, 
      N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, 
      N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, 
      N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, 
      N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, 
      N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, 
      N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, 
      N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, 
      N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, 
      N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N648, 
      N649, N714, N715, n1, n2, n3, n4, n5, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port, 
      n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113_port, n114_port, n115_port, n116_port, 
      n117_port, n118_port, n119_port, n120_port, n121_port, n122_port, 
      n123_port, n124_port, n125_port, n126_port, n127_port, n128_port, 
      n129_port, n130_port, n131_port, n132_port, n133_port, n134_port, 
      n135_port, n136_port, n137_port, n138_port, n139_port, n140_port, 
      n141_port, n142_port, n143_port, n144_port, n145_port, n146_port, 
      n147_port, n148_port, n149_port, n150_port, n151_port, n152_port, 
      n153_port, n154_port, n155_port, n156_port, n157_port, n158_port, 
      n159_port, n160_port, n161_port, n162_port, n163_port, n164_port, 
      n165_port, n166_port, n167_port, n168_port, n169_port, n170_port, 
      n171_port, n172_port, n173_port, n174_port, n175_port, n176_port, 
      n177_port, n178_port, n179_port, n180_port, n181_port, n182_port, 
      n183_port, n184_port, n185_port, n186_port, n187_port, n188_port, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204_port, n205_port, n206_port, 
      n207_port, n208_port, n209_port, n210_port, n211_port, n212_port, 
      n213_port, n214_port, n215_port, n216_port, n217_port, n218_port, 
      n219_port, n220_port, n221_port, n222_port, n223_port, n224_port, 
      n225_port, n226_port, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n300, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019 : 
      std_logic;

begin
   
   n1 <= '1';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   HI_LO_c_reg_HI_31_inst : HS65_LH_DFPRQX9 port map( D => n516, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_31_port);
   HI_LO_c_reg_HI_30_inst : HS65_LH_DFPRQX9 port map( D => n515, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_30_port);
   HI_LO_c_reg_HI_29_inst : HS65_LH_DFPRQX9 port map( D => n514, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_29_port);
   HI_LO_c_reg_HI_28_inst : HS65_LH_DFPRQX9 port map( D => n513, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_28_port);
   HI_LO_c_reg_HI_27_inst : HS65_LH_DFPRQX9 port map( D => n512, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_27_port);
   HI_LO_c_reg_HI_26_inst : HS65_LH_DFPRQX9 port map( D => n511, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_26_port);
   HI_LO_c_reg_HI_25_inst : HS65_LH_DFPRQX9 port map( D => n510, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_25_port);
   HI_LO_c_reg_HI_24_inst : HS65_LH_DFPRQX9 port map( D => n509, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_24_port);
   HI_LO_c_reg_HI_23_inst : HS65_LH_DFPRQX9 port map( D => n508, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_23_port);
   HI_LO_c_reg_HI_22_inst : HS65_LH_DFPRQX9 port map( D => n507, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_22_port);
   HI_LO_c_reg_HI_21_inst : HS65_LH_DFPRQX9 port map( D => n506, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_21_port);
   HI_LO_c_reg_HI_20_inst : HS65_LH_DFPRQX9 port map( D => n505, CP => clk, RN 
                           => n556, Q => HI_LO_c_HI_20_port);
   HI_LO_c_reg_HI_19_inst : HS65_LH_DFPRQX9 port map( D => n504, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_19_port);
   HI_LO_c_reg_HI_18_inst : HS65_LH_DFPRQX9 port map( D => n503, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_18_port);
   HI_LO_c_reg_HI_17_inst : HS65_LH_DFPRQX9 port map( D => n502, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_17_port);
   HI_LO_c_reg_HI_16_inst : HS65_LH_DFPRQX9 port map( D => n501, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_16_port);
   HI_LO_c_reg_HI_15_inst : HS65_LH_DFPRQX9 port map( D => n500, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_15_port);
   HI_LO_c_reg_HI_14_inst : HS65_LH_DFPRQX9 port map( D => n499, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_14_port);
   HI_LO_c_reg_HI_13_inst : HS65_LH_DFPRQX9 port map( D => n498, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_13_port);
   HI_LO_c_reg_HI_12_inst : HS65_LH_DFPRQX9 port map( D => n497, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_12_port);
   HI_LO_c_reg_HI_11_inst : HS65_LH_DFPRQX9 port map( D => n496, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_11_port);
   HI_LO_c_reg_HI_10_inst : HS65_LH_DFPRQX9 port map( D => n495, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_10_port);
   HI_LO_c_reg_HI_9_inst : HS65_LH_DFPRQX9 port map( D => n494, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_9_port);
   HI_LO_c_reg_HI_8_inst : HS65_LH_DFPRQX9 port map( D => n493, CP => clk, RN 
                           => n557, Q => HI_LO_c_HI_8_port);
   HI_LO_c_reg_HI_7_inst : HS65_LH_DFPRQX9 port map( D => n492, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_7_port);
   HI_LO_c_reg_HI_6_inst : HS65_LH_DFPRQX9 port map( D => n491, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_6_port);
   HI_LO_c_reg_HI_5_inst : HS65_LH_DFPRQX9 port map( D => n490, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_5_port);
   HI_LO_c_reg_HI_4_inst : HS65_LH_DFPRQX9 port map( D => n489, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_4_port);
   HI_LO_c_reg_HI_3_inst : HS65_LH_DFPRQX9 port map( D => n488, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_3_port);
   HI_LO_c_reg_HI_2_inst : HS65_LH_DFPRQX9 port map( D => n487, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_2_port);
   HI_LO_c_reg_HI_1_inst : HS65_LH_DFPRQX9 port map( D => n486, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_1_port);
   HI_LO_c_reg_HI_0_inst : HS65_LH_DFPRQX9 port map( D => n485, CP => clk, RN 
                           => n558, Q => HI_LO_c_HI_0_port);
   HI_LO_c_reg_LO_31_inst : HS65_LH_DFPRQX9 port map( D => n484, CP => clk, RN 
                           => n558, Q => HI_LO_c_LO_31_port);
   HI_LO_c_reg_LO_30_inst : HS65_LH_DFPRQX9 port map( D => n483, CP => clk, RN 
                           => n558, Q => HI_LO_c_LO_30_port);
   HI_LO_c_reg_LO_29_inst : HS65_LH_DFPRQX9 port map( D => n482, CP => clk, RN 
                           => n558, Q => HI_LO_c_LO_29_port);
   HI_LO_c_reg_LO_28_inst : HS65_LH_DFPRQX9 port map( D => n481, CP => clk, RN 
                           => n558, Q => HI_LO_c_LO_28_port);
   HI_LO_c_reg_LO_27_inst : HS65_LH_DFPRQX9 port map( D => n480, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_27_port);
   HI_LO_c_reg_LO_26_inst : HS65_LH_DFPRQX9 port map( D => n479, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_26_port);
   HI_LO_c_reg_LO_25_inst : HS65_LH_DFPRQX9 port map( D => n478, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_25_port);
   HI_LO_c_reg_LO_24_inst : HS65_LH_DFPRQX9 port map( D => n477, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_24_port);
   HI_LO_c_reg_LO_23_inst : HS65_LH_DFPRQX9 port map( D => n476, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_23_port);
   HI_LO_c_reg_LO_22_inst : HS65_LH_DFPRQX9 port map( D => n475, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_22_port);
   HI_LO_c_reg_LO_21_inst : HS65_LH_DFPRQX9 port map( D => n474, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_21_port);
   HI_LO_c_reg_LO_20_inst : HS65_LH_DFPRQX9 port map( D => n473, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_20_port);
   HI_LO_c_reg_LO_19_inst : HS65_LH_DFPRQX9 port map( D => n472, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_19_port);
   HI_LO_c_reg_LO_18_inst : HS65_LH_DFPRQX9 port map( D => n471, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_18_port);
   HI_LO_c_reg_LO_17_inst : HS65_LH_DFPRQX9 port map( D => n470, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_17_port);
   HI_LO_c_reg_LO_16_inst : HS65_LH_DFPRQX9 port map( D => n469, CP => clk, RN 
                           => n559, Q => HI_LO_c_LO_16_port);
   HI_LO_c_reg_LO_15_inst : HS65_LH_DFPRQX9 port map( D => n468, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_15_port);
   HI_LO_c_reg_LO_14_inst : HS65_LH_DFPRQX9 port map( D => n467, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_14_port);
   HI_LO_c_reg_LO_13_inst : HS65_LH_DFPRQX9 port map( D => n466, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_13_port);
   HI_LO_c_reg_LO_12_inst : HS65_LH_DFPRQX9 port map( D => n465, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_12_port);
   HI_LO_c_reg_LO_11_inst : HS65_LH_DFPRQX9 port map( D => n464, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_11_port);
   HI_LO_c_reg_LO_10_inst : HS65_LH_DFPRQX9 port map( D => n463, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_10_port);
   HI_LO_c_reg_LO_9_inst : HS65_LH_DFPRQX9 port map( D => n462, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_9_port);
   HI_LO_c_reg_LO_8_inst : HS65_LH_DFPRQX9 port map( D => n461, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_8_port);
   HI_LO_c_reg_LO_7_inst : HS65_LH_DFPRQX9 port map( D => n460, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_7_port);
   HI_LO_c_reg_LO_6_inst : HS65_LH_DFPRQX9 port map( D => n459, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_6_port);
   HI_LO_c_reg_LO_5_inst : HS65_LH_DFPRQX9 port map( D => n458, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_5_port);
   HI_LO_c_reg_LO_4_inst : HS65_LH_DFPRQX9 port map( D => n457, CP => clk, RN 
                           => n560, Q => HI_LO_c_LO_4_port);
   HI_LO_c_reg_LO_3_inst : HS65_LH_DFPRQX9 port map( D => n456, CP => clk, RN 
                           => n561, Q => HI_LO_c_LO_3_port);
   HI_LO_c_reg_LO_2_inst : HS65_LH_DFPRQX9 port map( D => n455, CP => clk, RN 
                           => n561, Q => HI_LO_c_LO_2_port);
   HI_LO_c_reg_LO_1_inst : HS65_LH_DFPRQX9 port map( D => n454, CP => clk, RN 
                           => n561, Q => HI_LO_c_LO_1_port);
   HI_LO_c_reg_LO_0_inst : HS65_LH_DFPRQX9 port map( D => n453, CP => clk, RN 
                           => n561, Q => HI_LO_c_LO_0_port);
   lt_136 : alu_DW_cmp_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => n552, A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => n550, A(25) => alu_i(67), A(24) 
                           => alu_i(66), A(23) => n548, A(22) => alu_i(64), 
                           A(21) => alu_i(63), A(20) => n546, A(19) => 
                           alu_i(61), A(18) => alu_i(60), A(17) => n544, A(16) 
                           => alu_i(58), A(15) => alu_i(57), A(14) => n542, 
                           A(13) => alu_i(55), A(12) => alu_i(54), A(11) => 
                           n540, A(10) => alu_i(52), A(9) => alu_i(51), A(8) =>
                           n538, A(7) => alu_i(49), A(6) => alu_i(48), A(5) => 
                           n536, A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           n534, A(1) => alu_i(43), A(0) => alu_i(42), B(31) =>
                           n532, B(30) => n531, B(29) => n530, B(28) => n528, 
                           B(27) => n526, B(26) => n525, B(25) => n524, B(24) 
                           => n523, B(23) => n522, B(22) => n521, B(21) => n520
                           , B(20) => n518, B(19) => n517, B(18) => n300, B(17)
                           => n90, B(16) => n89, B(15) => n88, B(14) => n87, 
                           B(13) => n86, B(12) => n85, B(11) => n83, B(10) => 
                           n82, B(9) => n81, B(8) => n80, B(7) => n79, B(6) => 
                           n78, B(5) => n77, B(4) => n75, B(3) => n73, B(2) => 
                           n71, B(1) => n70, B(0) => n69, TC => n1, GE_LT => n1
                           , GE_GT_EQ => n2, GE_LT_GT_LE => N648, EQ_NE => 
                           n_1014);
   sub_68 : alu_DW01_sub_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => n552, A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => n550, A(25) => alu_i(67), A(24) 
                           => alu_i(66), A(23) => n548, A(22) => alu_i(64), 
                           A(21) => alu_i(63), A(20) => n546, A(19) => 
                           alu_i(61), A(18) => alu_i(60), A(17) => n544, A(16) 
                           => alu_i(58), A(15) => alu_i(57), A(14) => n542, 
                           A(13) => alu_i(55), A(12) => alu_i(54), A(11) => 
                           n540, A(10) => alu_i(52), A(9) => alu_i(51), A(8) =>
                           n538, A(7) => alu_i(49), A(6) => alu_i(48), A(5) => 
                           n536, A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           n534, A(1) => alu_i(43), A(0) => alu_i(42), B(31) =>
                           n532, B(30) => n531, B(29) => n530, B(28) => n528, 
                           B(27) => n526, B(26) => n525, B(25) => n524, B(24) 
                           => n523, B(23) => n522, B(22) => n521, B(21) => n520
                           , B(20) => n518, B(19) => n517, B(18) => n300, B(17)
                           => n90, B(16) => n89, B(15) => n88, B(14) => n87, 
                           B(13) => n86, B(12) => n85, B(11) => n83, B(10) => 
                           n82, B(9) => n81, B(8) => n80, B(7) => n79, B(6) => 
                           n78, B(5) => n77, B(4) => n75, B(3) => n73, B(2) => 
                           n71, B(1) => n70, B(0) => n69, CI => n3, DIFF(31) =>
                           N162, DIFF(30) => N161, DIFF(29) => N160, DIFF(28) 
                           => N159, DIFF(27) => N158, DIFF(26) => N157, 
                           DIFF(25) => N156, DIFF(24) => N155, DIFF(23) => N154
                           , DIFF(22) => N153, DIFF(21) => N152, DIFF(20) => 
                           N151, DIFF(19) => N150, DIFF(18) => N149, DIFF(17) 
                           => N148, DIFF(16) => N147, DIFF(15) => N146, 
                           DIFF(14) => N145, DIFF(13) => N144, DIFF(12) => N143
                           , DIFF(11) => N142, DIFF(10) => N141, DIFF(9) => 
                           N140, DIFF(8) => N139, DIFF(7) => N138, DIFF(6) => 
                           N137, DIFF(5) => N136, DIFF(4) => N135, DIFF(3) => 
                           N134, DIFF(2) => N133, DIFF(1) => N132, DIFF(0) => 
                           N131, CO => n_1015);
   r325 : alu_DW01_cmp6_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => n552, A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => n550, A(25) => alu_i(67), A(24) 
                           => alu_i(66), A(23) => n548, A(22) => alu_i(64), 
                           A(21) => alu_i(63), A(20) => n546, A(19) => 
                           alu_i(61), A(18) => alu_i(60), A(17) => n544, A(16) 
                           => alu_i(58), A(15) => alu_i(57), A(14) => n542, 
                           A(13) => alu_i(55), A(12) => alu_i(54), A(11) => 
                           n540, A(10) => alu_i(52), A(9) => alu_i(51), A(8) =>
                           n538, A(7) => alu_i(49), A(6) => alu_i(48), A(5) => 
                           n536, A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           n534, A(1) => alu_i(43), A(0) => alu_i(42), B(31) =>
                           n532, B(30) => n531, B(29) => n530, B(28) => n528, 
                           B(27) => n526, B(26) => n525, B(25) => n524, B(24) 
                           => n523, B(23) => n522, B(22) => n521, B(21) => n520
                           , B(20) => n518, B(19) => n517, B(18) => n300, B(17)
                           => n90, B(16) => n89, B(15) => n88, B(14) => n87, 
                           B(13) => n86, B(12) => n85, B(11) => n83, B(10) => 
                           n82, B(9) => n81, B(8) => n80, B(7) => n79, B(6) => 
                           n78, B(5) => n77, B(4) => n75, B(3) => n73, B(2) => 
                           n71, B(1) => n70, B(0) => n69, TC => n4, LT => N649,
                           GT => n_1016, EQ => N714, LE => n_1017, GE => n_1018
                           , NE => N715);
   r321 : alu_DW01_add_0 port map( A(31) => alu_i(73), A(30) => alu_i(72), 
                           A(29) => n552, A(28) => alu_i(70), A(27) => 
                           alu_i(69), A(26) => n550, A(25) => alu_i(67), A(24) 
                           => alu_i(66), A(23) => n548, A(22) => alu_i(64), 
                           A(21) => alu_i(63), A(20) => n546, A(19) => 
                           alu_i(61), A(18) => alu_i(60), A(17) => n544, A(16) 
                           => alu_i(58), A(15) => alu_i(57), A(14) => n542, 
                           A(13) => alu_i(55), A(12) => alu_i(54), A(11) => 
                           n540, A(10) => alu_i(52), A(9) => alu_i(51), A(8) =>
                           n538, A(7) => alu_i(49), A(6) => alu_i(48), A(5) => 
                           n536, A(4) => alu_i(46), A(3) => alu_i(45), A(2) => 
                           n534, A(1) => alu_i(43), A(0) => alu_i(42), B(31) =>
                           n532, B(30) => n531, B(29) => n530, B(28) => n528, 
                           B(27) => n526, B(26) => n525, B(25) => n524, B(24) 
                           => n523, B(23) => n522, B(22) => n521, B(21) => n520
                           , B(20) => n518, B(19) => n517, B(18) => n300, B(17)
                           => n90, B(16) => n89, B(15) => n88, B(14) => n87, 
                           B(13) => n86, B(12) => n85, B(11) => n83, B(10) => 
                           n82, B(9) => n81, B(8) => n80, B(7) => n79, B(6) => 
                           n78, B(5) => n77, B(4) => n75, B(3) => n73, B(2) => 
                           n71, B(1) => n70, B(0) => n69, CI => n5, SUM(31) => 
                           N130, SUM(30) => N129, SUM(29) => N128, SUM(28) => 
                           N127, SUM(27) => N126, SUM(26) => N125, SUM(25) => 
                           N124, SUM(24) => N123, SUM(23) => N122, SUM(22) => 
                           N121, SUM(21) => N120, SUM(20) => N119, SUM(19) => 
                           N118, SUM(18) => N117, SUM(17) => N116, SUM(16) => 
                           N115, SUM(15) => N114, SUM(14) => N113, SUM(13) => 
                           N112, SUM(12) => N111, SUM(11) => N110, SUM(10) => 
                           N109, SUM(9) => N108, SUM(8) => N107, SUM(7) => N106
                           , SUM(6) => N105, SUM(5) => N104, SUM(4) => N103, 
                           SUM(3) => N102, SUM(2) => N101, SUM(1) => N100, 
                           SUM(0) => N99, CO => n_1019);
   mult_71 : alu_DW_mult_uns_0 port map( a(31) => alu_i(73), a(30) => alu_i(72)
                           , a(29) => n552, a(28) => alu_i(70), a(27) => 
                           alu_i(69), a(26) => n550, a(25) => alu_i(67), a(24) 
                           => alu_i(66), a(23) => n548, a(22) => alu_i(64), 
                           a(21) => alu_i(63), a(20) => n546, a(19) => 
                           alu_i(61), a(18) => alu_i(60), a(17) => n544, a(16) 
                           => alu_i(58), a(15) => alu_i(57), a(14) => n542, 
                           a(13) => alu_i(55), a(12) => alu_i(54), a(11) => 
                           n540, a(10) => alu_i(52), a(9) => alu_i(51), a(8) =>
                           n538, a(7) => alu_i(49), a(6) => alu_i(48), a(5) => 
                           n536, a(4) => alu_i(46), a(3) => alu_i(45), a(2) => 
                           n534, a(1) => alu_i(43), a(0) => alu_i(42), b(31) =>
                           n532, b(30) => n531, b(29) => n530, b(28) => n528, 
                           b(27) => n526, b(26) => n525, b(25) => n524, b(24) 
                           => n523, b(23) => n522, b(22) => n521, b(21) => n520
                           , b(20) => n518, b(19) => n517, b(18) => n300, b(17)
                           => n90, b(16) => n89, b(15) => n88, b(14) => n87, 
                           b(13) => n86, b(12) => n85, b(11) => n83, b(10) => 
                           n82, b(9) => n81, b(8) => n80, b(7) => n79, b(6) => 
                           n78, b(5) => n77, b(4) => n75, b(3) => n73, b(2) => 
                           n71, b(1) => n70, b(0) => n69, product(63) => N226, 
                           product(62) => N225, product(61) => N224, 
                           product(60) => N223, product(59) => N222, 
                           product(58) => N221, product(57) => N220, 
                           product(56) => N219, product(55) => N218, 
                           product(54) => N217, product(53) => N216, 
                           product(52) => N215, product(51) => N214, 
                           product(50) => N213, product(49) => N212, 
                           product(48) => N211, product(47) => N210, 
                           product(46) => N209, product(45) => N208, 
                           product(44) => N207, product(43) => N206, 
                           product(42) => N205, product(41) => N204, 
                           product(40) => N203, product(39) => N202, 
                           product(38) => N201, product(37) => N200, 
                           product(36) => N199, product(35) => N198, 
                           product(34) => N197, product(33) => N196, 
                           product(32) => N195, product(31) => N194, 
                           product(30) => N193, product(29) => N192, 
                           product(28) => N191, product(27) => N190, 
                           product(26) => N189, product(25) => N188, 
                           product(24) => N187, product(23) => N186, 
                           product(22) => N185, product(21) => N184, 
                           product(20) => N183, product(19) => N182, 
                           product(18) => N181, product(17) => N180, 
                           product(16) => N179, product(15) => N178, 
                           product(14) => N177, product(13) => N176, 
                           product(12) => N175, product(11) => N174, 
                           product(10) => N173, product(9) => N172, product(8) 
                           => N171, product(7) => N170, product(6) => N169, 
                           product(5) => N168, product(4) => N167, product(3) 
                           => N166, product(2) => N165, product(1) => N164, 
                           product(0) => N163);
   U3 : HS65_LH_NOR4ABX2 port map( A => n92, B => n93, C => n94, D => n95, Z =>
                           n91);
   U4 : HS65_LH_IVX9 port map( A => n537, Z => n536);
   U5 : HS65_LH_IVX9 port map( A => n76, Z => n75);
   U6 : HS65_LH_IVX9 port map( A => n74, Z => n73);
   U7 : HS65_LH_IVX9 port map( A => n541, Z => n540);
   U13 : HS65_LH_IVX9 port map( A => n545, Z => n544);
   U14 : HS65_LH_IVX9 port map( A => n539, Z => n538);
   U15 : HS65_LH_IVX9 port map( A => n543, Z => n542);
   U16 : HS65_LH_IVX9 port map( A => n72, Z => n71);
   U17 : HS65_LH_IVX9 port map( A => n84, Z => n83);
   U18 : HS65_LH_IVX9 port map( A => n547, Z => n546);
   U19 : HS65_LH_IVX9 port map( A => n551, Z => n550);
   U20 : HS65_LH_IVX9 port map( A => n553, Z => n552);
   U21 : HS65_LH_IVX9 port map( A => n519, Z => n518);
   U22 : HS65_LH_IVX9 port map( A => n527, Z => n526);
   U23 : HS65_LH_IVX9 port map( A => n529, Z => n528);
   U24 : HS65_LH_IVX9 port map( A => n533, Z => n532);
   U25 : HS65_LH_NOR4ABX4 port map( A => n612, B => n435, C => alu_i(8), D => 
                           alu_i(7), Z => n180_port);
   U26 : HS65_LH_BFX9 port map( A => alu_i(11), Z => n70);
   U27 : HS65_LH_BFX9 port map( A => alu_i(18), Z => n80);
   U28 : HS65_LH_BFX9 port map( A => alu_i(15), Z => n77);
   U29 : HS65_LH_BFX9 port map( A => alu_i(16), Z => n78);
   U30 : HS65_LH_BFX9 port map( A => alu_i(17), Z => n79);
   U31 : HS65_LH_BFX9 port map( A => alu_i(20), Z => n82);
   U32 : HS65_LH_BFX9 port map( A => alu_i(22), Z => n85);
   U33 : HS65_LH_BFX9 port map( A => alu_i(23), Z => n86);
   U34 : HS65_LH_BFX9 port map( A => alu_i(24), Z => n87);
   U35 : HS65_LH_BFX9 port map( A => alu_i(25), Z => n88);
   U36 : HS65_LH_BFX9 port map( A => alu_i(19), Z => n81);
   U37 : HS65_LH_BFX9 port map( A => alu_i(29), Z => n517);
   U38 : HS65_LH_BFX9 port map( A => alu_i(26), Z => n89);
   U39 : HS65_LH_BFX9 port map( A => alu_i(27), Z => n90);
   U40 : HS65_LH_BFX9 port map( A => alu_i(28), Z => n300);
   U41 : HS65_LH_BFX9 port map( A => alu_i(31), Z => n520);
   U42 : HS65_LH_BFX9 port map( A => alu_i(33), Z => n522);
   U43 : HS65_LH_BFX9 port map( A => alu_i(35), Z => n524);
   U44 : HS65_LH_BFX9 port map( A => alu_i(32), Z => n521);
   U45 : HS65_LH_BFX9 port map( A => alu_i(34), Z => n523);
   U46 : HS65_LH_BFX9 port map( A => alu_i(36), Z => n525);
   U47 : HS65_LH_BFX9 port map( A => alu_i(39), Z => n530);
   U48 : HS65_LH_BFX9 port map( A => alu_i(40), Z => n531);
   U49 : HS65_LH_NOR2X6 port map( A => n98, B => alu_i(4), Z => n284);
   U50 : HS65_LH_IVX9 port map( A => n61, Z => n60);
   U51 : HS65_LH_IVX9 port map( A => n61, Z => n59);
   U52 : HS65_LH_IVX9 port map( A => n62, Z => n58);
   U53 : HS65_LH_IVX9 port map( A => n62, Z => n57);
   U54 : HS65_LH_IVX9 port map( A => n98, Z => n605);
   U55 : HS65_LH_IVX9 port map( A => n56, Z => n55);
   U56 : HS65_LH_IVX9 port map( A => n42, Z => n41);
   U57 : HS65_LH_IVX9 port map( A => n42, Z => n40);
   U58 : HS65_LH_BFX9 port map( A => n68, Z => n61);
   U59 : HS65_LH_BFX9 port map( A => n68, Z => n62);
   U60 : HS65_LH_BFX9 port map( A => n604, Z => n12);
   U61 : HS65_LH_BFX9 port map( A => n604, Z => n11);
   U62 : HS65_LH_BFX9 port map( A => n603, Z => n8);
   U63 : HS65_LH_BFX9 port map( A => n603, Z => n9);
   U64 : HS65_LH_BFX9 port map( A => n67, Z => n65);
   U65 : HS65_LH_BFX9 port map( A => n67, Z => n64);
   U66 : HS65_LH_BFX9 port map( A => n68, Z => n63);
   U67 : HS65_LH_BFX9 port map( A => n604, Z => n13);
   U68 : HS65_LH_BFX9 port map( A => n603, Z => n10);
   U69 : HS65_LH_BFX9 port map( A => n67, Z => n66);
   U70 : HS65_LH_BFX9 port map( A => n555, Z => n560);
   U71 : HS65_LH_BFX9 port map( A => n555, Z => n559);
   U72 : HS65_LH_BFX9 port map( A => n554, Z => n558);
   U73 : HS65_LH_BFX9 port map( A => n554, Z => n557);
   U74 : HS65_LH_BFX9 port map( A => n554, Z => n556);
   U75 : HS65_LH_BFX9 port map( A => n555, Z => n561);
   U76 : HS65_LH_IVX9 port map( A => n101_port, Z => n603);
   U77 : HS65_LH_IVX9 port map( A => n100_port, Z => n604);
   U78 : HS65_LH_NAND2X7 port map( A => n442, B => n435, Z => n98);
   U79 : HS65_LH_IVX9 port map( A => n96, Z => n606);
   U80 : HS65_LH_NOR3X4 port map( A => n48, B => n45, C => n106_port, Z => n92)
                           ;
   U81 : HS65_LH_IVX9 port map( A => n176_port, Z => n597);
   U82 : HS65_LH_IVX9 port map( A => n281, Z => n598);
   U83 : HS65_LH_IVX9 port map( A => n54, Z => n56);
   U84 : HS65_LH_IVX9 port map( A => n39, Z => n42);
   U85 : HS65_LH_BFX9 port map( A => n43, Z => n44);
   U86 : HS65_LH_BFX9 port map( A => n91, Z => n68);
   U87 : HS65_LH_BFX9 port map( A => n91, Z => n67);
   U88 : HS65_LH_BFX9 port map( A => n50, Z => n52);
   U89 : HS65_LH_BFX9 port map( A => n50, Z => n51);
   U90 : HS65_LH_BFX9 port map( A => n608, Z => n15);
   U91 : HS65_LH_BFX9 port map( A => n608, Z => n14);
   U92 : HS65_LH_BFX9 port map( A => n43, Z => n45);
   U93 : HS65_LH_BFX9 port map( A => n50, Z => n53);
   U94 : HS65_LH_BFX9 port map( A => rst_n, Z => n555);
   U95 : HS65_LH_BFX9 port map( A => rst_n, Z => n554);
   U96 : HS65_LH_IVX9 port map( A => n237, Z => n592);
   U97 : HS65_LH_AO222X4 port map( A => n128_port, B => n115_port, C => 
                           n133_port, D => n118_port, E => n174_port, F => 
                           n117_port, Z => n170_port);
   U98 : HS65_LH_IVX9 port map( A => n317, Z => n582);
   U99 : HS65_LH_IVX9 port map( A => n144_port, Z => n572);
   U100 : HS65_LH_IVX9 port map( A => n130_port, Z => n579);
   U101 : HS65_LH_IVX9 port map( A => n212_port, Z => n575);
   U102 : HS65_LH_NOR4ABX2 port map( A => n100_port, B => n101_port, C => 
                           n102_port, D => n103_port, Z => n93);
   U103 : HS65_LH_NAND3X5 port map( A => n96, B => n54, C => n98, Z => n95);
   U104 : HS65_LH_NAND4ABX3 port map( A => n42, B => n53, C => n612, D => n15, 
                           Z => n94);
   U105 : HS65_LH_NOR2X6 port map( A => n96, B => n189_port, Z => n279);
   U106 : HS65_LH_IVX9 port map( A => n180_port, Z => n608);
   U107 : HS65_LH_NAND2X7 port map( A => n436, B => n442, Z => n96);
   U108 : HS65_LH_NOR2X6 port map( A => n189_port, B => n98, Z => n115_port);
   U109 : HS65_LH_NOR2X6 port map( A => n611, B => n609, Z => n435);
   U110 : HS65_LH_IVX9 port map( A => n208_port, Z => n600);
   U111 : HS65_LH_AND2X4 port map( A => n390, B => n391, Z => n106_port);
   U112 : HS65_LH_IVX9 port map( A => n186_port, Z => n599);
   U113 : HS65_LH_NAND2X7 port map( A => n195_port, B => n605, Z => n176_port);
   U114 : HS65_LH_AND2X4 port map( A => n445, B => n607, Z => n442);
   U115 : HS65_LH_NAND2X7 port map( A => n606, B => n195_port, Z => n281);
   U116 : HS65_LH_IVX9 port map( A => n189_port, Z => n595);
   U117 : HS65_LH_NAND2X7 port map( A => n434, B => n438, Z => n101_port);
   U118 : HS65_LH_AND2X4 port map( A => n275, B => n16, Z => n368);
   U119 : HS65_LH_AND2X4 port map( A => n117_port, B => n16, Z => n397);
   U120 : HS65_LH_NAND2X7 port map( A => n434, B => n435, Z => n100_port);
   U121 : HS65_LH_BFX9 port map( A => n123_port, Z => n39);
   U122 : HS65_LH_NAND2X7 port map( A => n438, B => n442, Z => n123_port);
   U123 : HS65_LH_BFX9 port map( A => n97, Z => n54);
   U124 : HS65_LH_NAND2X7 port map( A => n391, B => n442, Z => n97);
   U125 : HS65_LH_IVX9 port map( A => n438, Z => n610);
   U126 : HS65_LH_BFX9 port map( A => n105_port, Z => n43);
   U127 : HS65_LH_NOR2AX3 port map( A => n390, B => n610, Z => n105_port);
   U128 : HS65_LH_BFX9 port map( A => n99_port, Z => n50);
   U129 : HS65_LH_NOR2X6 port map( A => n609, B => n437, Z => n99_port);
   U130 : HS65_LH_IVX9 port map( A => n38, Z => n36);
   U131 : HS65_LH_BFX9 port map( A => n46, Z => n48);
   U132 : HS65_LH_BFX9 port map( A => n46, Z => n47);
   U133 : HS65_LH_AND2X4 port map( A => n434, B => n391, Z => n102_port);
   U134 : HS65_LH_BFX9 port map( A => n29, Z => n31);
   U135 : HS65_LH_BFX9 port map( A => n29, Z => n32);
   U136 : HS65_LH_BFX9 port map( A => n30, Z => n33);
   U137 : HS65_LH_IVX9 port map( A => n38, Z => n37);
   U138 : HS65_LH_AND2X4 port map( A => n434, B => n436, Z => n103_port);
   U139 : HS65_LH_BFX9 port map( A => n18, Z => n20);
   U140 : HS65_LH_BFX9 port map( A => n18, Z => n22);
   U141 : HS65_LH_BFX9 port map( A => n18, Z => n21);
   U142 : HS65_LH_BFX9 port map( A => n19, Z => n23);
   U143 : HS65_LH_BFX9 port map( A => n19, Z => n24);
   U144 : HS65_LH_BFX9 port map( A => n46, Z => n49);
   U145 : HS65_LH_BFX9 port map( A => n30, Z => n34);
   U146 : HS65_LH_IVX9 port map( A => n535, Z => n534);
   U147 : HS65_LH_IVX9 port map( A => n549, Z => n548);
   U148 : HS65_LH_AO112X9 port map( A => N714, B => n450, C => n451, D => n452,
                           Z => alu_o(32));
   U149 : HS65_LH_AO222X4 port map( A => n391, B => n450, C => n438, D => n450,
                           E => n436, F => n450, Z => n452);
   U150 : HS65_LH_NOR3X4 port map( A => alu_i(7), B => alu_i(8), C => n612, Z 
                           => n450);
   U151 : HS65_LH_NOR4ABX2 port map( A => N715, B => n607, C => n612, D => n610
                           , Z => n451);
   U152 : HS65_LH_AOI222X2 port map( A => n31, B => n70, C => n26, D => n69, E 
                           => n35, F => n71, Z => n237);
   U153 : HS65_LH_AOI212X4 port map( A => alu_i(46), B => n180_port, C => n56, 
                           D => n589, E => n42, Z => n175_port);
   U154 : HS65_LH_IVX9 port map( A => alu_i(46), Z => n589);
   U155 : HS65_LH_AOI212X4 port map( A => n540, B => n180_port, C => n56, D => 
                           n541, E => n42, Z => n421);
   U156 : HS65_LH_AOI212X4 port map( A => n546, B => n180_port, C => n56, D => 
                           n547, E => n42, Z => n350);
   U157 : HS65_LH_AOI212X4 port map( A => alu_i(69), B => n180_port, C => n56, 
                           D => n567, E => n42, Z => n280);
   U158 : HS65_LH_IVX9 port map( A => alu_i(69), Z => n567);
   U159 : HS65_LH_OAI212X5 port map( A => n585, B => n189_port, C => n190_port,
                           D => n596, E => n191_port, Z => n183_port);
   U160 : HS65_LH_IVX9 port map( A => n140_port, Z => n585);
   U161 : HS65_LH_AOI222X2 port map( A => n192_port, B => n145_port, C => 
                           n193_port, D => n194_port, E => n195_port, F => 
                           n142_port, Z => n191_port);
   U162 : HS65_LH_MX41X7 port map( D0 => n73, S0 => n36, D1 => n75, S1 => n32, 
                           D2 => n77, S2 => n27, D3 => n78, S3 => n22, Z => 
                           n194_port);
   U163 : HS65_LH_OAI212X5 port map( A => n570, B => n189_port, C => n264, D =>
                           n596, E => n265, Z => n259);
   U164 : HS65_LH_IVX9 port map( A => n269, Z => n570);
   U165 : HS65_LH_AOI222X2 port map( A => n192_port, B => n266, C => n193_port,
                           D => n267, E => n195_port, F => n268, Z => n265);
   U166 : HS65_LH_MX41X7 port map( D0 => n528, S0 => n196_port, D1 => n526, S1 
                           => n31, D2 => n525, S2 => n26, D3 => n524, S3 => n20
                           , Z => n267);
   U167 : HS65_LH_OAI212X5 port map( A => n236, B => n72, C => n237, D => 
                           n186_port, E => n238, Z => n235);
   U168 : HS65_LH_CBI4I1X5 port map( A => n56, B => n72, C => n42, D => n534, Z
                           => n238);
   U169 : HS65_LH_AOI212X4 port map( A => n534, B => n180_port, C => n56, D => 
                           n535, E => n42, Z => n236);
   U170 : HS65_LH_OAI212X5 port map( A => n185_port, B => n74, C => n591, D => 
                           n186_port, E => n187_port, Z => n184_port);
   U171 : HS65_LH_CBI4I1X5 port map( A => n56, B => n74, C => n42, D => 
                           alu_i(45), Z => n187_port);
   U172 : HS65_LH_AOI212X4 port map( A => alu_i(45), B => n180_port, C => n56, 
                           D => n590, E => n42, Z => n185_port);
   U173 : HS65_LH_IVX9 port map( A => n188_port, Z => n591);
   U174 : HS65_LH_OAI212X5 port map( A => n261, B => n529, C => n564, D => 
                           n208_port, E => n262, Z => n260);
   U175 : HS65_LH_CBI4I1X5 port map( A => n56, B => n529, C => n42, D => 
                           alu_i(70), Z => n262);
   U176 : HS65_LH_AOI212X4 port map( A => alu_i(70), B => n180_port, C => n56, 
                           D => n566, E => n42, Z => n261);
   U177 : HS65_LH_IVX9 port map( A => n263, Z => n564);
   U178 : HS65_LH_OAI212X5 port map( A => n552, B => n97, C => n14, D => n553, 
                           E => n41, Z => n248);
   U179 : HS65_LH_AOI32X5 port map( A => n283, B => n601, C => n284, D => 
                           alu_i(69), E => n285, Z => n282);
   U180 : HS65_LH_OAI21X3 port map( A => n526, B => n55, C => n41, Z => n285);
   U181 : HS65_LH_OAI212X5 port map( A => alu_i(58), B => n55, C => n15, D => 
                           n577, E => n41, Z => n388);
   U182 : HS65_LH_IVX9 port map( A => alu_i(58), Z => n577);
   U183 : HS65_LH_OAI212X5 port map( A => alu_i(57), B => n55, C => n15, D => 
                           n578, E => n40, Z => n396);
   U184 : HS65_LH_IVX9 port map( A => alu_i(57), Z => n578);
   U185 : HS65_LH_OAI212X5 port map( A => alu_i(54), B => n55, C => n15, D => 
                           n581, E => n40, Z => n415);
   U186 : HS65_LH_IVX9 port map( A => alu_i(54), Z => n581);
   U187 : HS65_LH_OAI212X5 port map( A => alu_i(55), B => n55, C => n15, D => 
                           n580, E => n40, Z => n409);
   U188 : HS65_LH_IVX9 port map( A => alu_i(55), Z => n580);
   U189 : HS65_LH_OAI212X5 port map( A => n542, B => n55, C => n15, D => n543, 
                           E => n40, Z => n403);
   U190 : HS65_LH_OAI212X5 port map( A => n544, B => n55, C => n15, D => n545, 
                           E => n123_port, Z => n381);
   U191 : HS65_LH_OAI212X5 port map( A => alu_i(61), B => n55, C => n15, D => 
                           n574, E => n40, Z => n367);
   U192 : HS65_LH_IVX9 port map( A => alu_i(61), Z => n574);
   U193 : HS65_LH_OAI212X5 port map( A => alu_i(64), B => n55, C => n14, D => 
                           n571, E => n41, Z => n338);
   U194 : HS65_LH_IVX9 port map( A => alu_i(64), Z => n571);
   U195 : HS65_LH_OAI212X5 port map( A => n536, B => n54, C => n14, D => n537, 
                           E => n41, Z => n167_port);
   U196 : HS65_LH_OAI212X5 port map( A => alu_i(49), B => n54, C => n14, D => 
                           n587, E => n41, Z => n146_port);
   U197 : HS65_LH_IVX9 port map( A => alu_i(49), Z => n587);
   U198 : HS65_LH_OAI212X5 port map( A => n538, B => n54, C => n14, D => n539, 
                           E => n41, Z => n134_port);
   U199 : HS65_LH_OAI212X5 port map( A => alu_i(51), B => n54, C => n586, D => 
                           n15, E => n41, Z => n121_port);
   U200 : HS65_LH_IVX9 port map( A => alu_i(51), Z => n586);
   U201 : HS65_LH_OAI212X5 port map( A => n548, B => n54, C => n14, D => n549, 
                           E => n41, Z => n328);
   U202 : HS65_LH_OAI212X5 port map( A => n550, B => n54, C => n14, D => n551, 
                           E => n41, Z => n293);
   U203 : HS65_LH_OAI212X5 port map( A => alu_i(52), B => n55, C => n15, D => 
                           n584, E => n41, Z => n428);
   U204 : HS65_LH_IVX9 port map( A => alu_i(52), Z => n584);
   U205 : HS65_LH_OAI212X5 port map( A => alu_i(67), B => n55, C => n14, D => 
                           n568, E => n41, Z => n307);
   U206 : HS65_LH_IVX9 port map( A => alu_i(67), Z => n568);
   U207 : HS65_LH_AOI32X5 port map( A => n178_port, B => n601, C => n275, D => 
                           n546, E => n352, Z => n351);
   U208 : HS65_LH_OAI21X3 port map( A => n518, B => n55, C => n123_port, Z => 
                           n352);
   U209 : HS65_LH_AOI32X5 port map( A => n178_port, B => n601, C => n113_port, 
                           D => alu_i(46), E => n179_port, Z => n177_port);
   U210 : HS65_LH_OAI21X3 port map( A => n75, B => n55, C => n39, Z => 
                           n179_port);
   U211 : HS65_LH_AOI32X5 port map( A => n283, B => n601, C => n117_port, D => 
                           n540, E => n423, Z => n422);
   U212 : HS65_LH_OAI21X3 port map( A => n83, B => n55, C => n40, Z => n423);
   U213 : HS65_LH_MX41X7 port map( D0 => n85, S0 => n37, D1 => n83, S1 => n33, 
                           D2 => n82, S2 => n28, D3 => n20, S3 => n81, Z => 
                           n317);
   U214 : HS65_LH_MX41X7 port map( D0 => n80, S0 => n37, D1 => n79, S1 => n33, 
                           D2 => n78, S2 => n27, D3 => n77, S3 => n22, Z => 
                           n316);
   U215 : HS65_LH_MX41X7 port map( D0 => n88, S0 => n37, D1 => n89, S1 => n33, 
                           D2 => n90, S2 => n28, D3 => n300, S3 => n23, Z => 
                           n145_port);
   U216 : HS65_LH_MX41X7 port map( D0 => n89, S0 => n36, D1 => n88, S1 => n32, 
                           D2 => n87, S2 => n27, D3 => n86, S3 => n21, Z => 
                           n266);
   U217 : HS65_LH_MX41X7 port map( D0 => n88, S0 => n36, D1 => n87, S1 => n32, 
                           D2 => n86, S2 => n27, D3 => n85, S3 => n21, Z => 
                           n278);
   U218 : HS65_LH_NOR2AX3 port map( A => n69, B => n38, Z => n315);
   U219 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n517, D1 => n31, S1 
                           => n518, D2 => n520, S2 => n28, D3 => n521, S3 => 
                           n23, Z => n144_port);
   U220 : HS65_LH_MX41X7 port map( D0 => n528, S0 => n37, D1 => n530, S1 => n33
                           , D2 => n531, S2 => n28, D3 => n532, S3 => n24, Z =>
                           n263);
   U221 : HS65_LH_MX41X7 port map( D0 => n73, S0 => n37, D1 => n71, S1 => n33, 
                           D2 => n70, S2 => n28, D3 => n69, S3 => n23, Z => 
                           n188_port);
   U222 : HS65_LH_MX41X7 port map( D0 => n85, S0 => n37, D1 => n86, S1 => n33, 
                           D2 => n87, S2 => n28, D3 => n88, S3 => n24, Z => 
                           n130_port);
   U223 : HS65_LH_MX41X7 port map( D0 => n35, S0 => n517, D1 => n300, S1 => n32
                           , D2 => n90, S2 => n27, D3 => n89, S3 => n21, Z => 
                           n212_port);
   U224 : HS65_LH_MX41X7 port map( D0 => n522, S0 => n37, D1 => n523, S1 => n33
                           , D2 => n524, S2 => n28, D3 => n525, S3 => n23, Z =>
                           n325);
   U225 : HS65_LH_MX41X7 port map( D0 => n87, S0 => n37, D1 => n88, S1 => n33, 
                           D2 => n89, S2 => n28, D3 => n90, S3 => n23, Z => 
                           n157_port);
   U226 : HS65_LH_MX41X7 port map( D0 => n86, S0 => n36, D1 => n87, S1 => n32, 
                           D2 => n88, S2 => n27, D3 => n89, S3 => n22, Z => 
                           n114_port);
   U227 : HS65_LH_MX41X7 port map( D0 => n83, S0 => n37, D1 => n85, S1 => n33, 
                           D2 => n86, S2 => n28, D3 => n87, S3 => n22, Z => 
                           n142_port);
   U228 : HS65_LH_MX41X7 port map( D0 => n77, S0 => n36, D1 => n75, S1 => n32, 
                           D2 => n73, S2 => n27, D3 => n71, S3 => n22, Z => 
                           n302);
   U229 : HS65_LH_MX41X7 port map( D0 => n78, S0 => n37, D1 => n77, S1 => n33, 
                           D2 => n75, S2 => n28, D3 => n73, S3 => n23, Z => 
                           n336);
   U230 : HS65_LH_MX41X7 port map( D0 => n79, S0 => n37, D1 => n78, S1 => n33, 
                           D2 => n77, S2 => n28, D3 => n75, S3 => n23, Z => 
                           n326);
   U231 : HS65_LH_MX41X7 port map( D0 => n35, S0 => n300, D1 => n90, S1 => n32,
                           D2 => n89, S2 => n27, D3 => n88, S3 => n21, Z => 
                           n229);
   U232 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n518, D1 => n31, S1 
                           => n517, D2 => n300, S2 => n27, D3 => n90, S3 => n21
                           , Z => n268);
   U233 : HS65_LH_MX41X7 port map( D0 => n90, S0 => n36, D1 => n89, S1 => n32, 
                           D2 => n88, S2 => n27, D3 => n87, S3 => n21, Z => 
                           n254);
   U234 : HS65_LH_MX41X7 port map( D0 => n87, S0 => n36, D1 => n86, S1 => n32, 
                           D2 => n85, S2 => n27, D3 => n83, S3 => n22, Z => 
                           n292);
   U235 : HS65_LH_MX41X7 port map( D0 => n86, S0 => n36, D1 => n85, S1 => n32, 
                           D2 => n83, S2 => n27, D3 => n82, S3 => n22, Z => 
                           n306);
   U236 : HS65_LH_CBI4I6X5 port map( A => n530, B => n54, C => n40, D => n553, 
                           Z => n249);
   U237 : HS65_LH_AO222X4 port map( A => n33, B => n531, C => n26, D => n532, E
                           => n35, F => n530, Z => n247);
   U238 : HS65_LH_NOR2X6 port map( A => n533, B => n38, Z => n216_port);
   U239 : HS65_LH_MX41X7 port map( D0 => n523, S0 => n37, D1 => n524, S1 => n33
                           , D2 => n525, S2 => n28, D3 => n526, S3 => n24, Z =>
                           n313);
   U240 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n81, D1 => n82, S1 =>
                           n32, D2 => n83, S2 => n27, D3 => n85, S3 => n21, Z 
                           => n111_port);
   U241 : HS65_LH_MX41X7 port map( D0 => n82, S0 => n37, D1 => n83, S1 => n33, 
                           D2 => n85, S2 => n28, D3 => n86, S3 => n23, Z => 
                           n154_port);
   U242 : HS65_LH_MX41X7 port map( D0 => n524, S0 => n36, D1 => n525, S1 => n32
                           , D2 => n526, S2 => n27, D3 => n528, S3 => n22, Z =>
                           n299);
   U243 : HS65_LH_MX41X7 port map( D0 => n525, S0 => n37, D1 => n526, S1 => n33
                           , D2 => n528, S2 => n28, D3 => n530, S3 => n23, Z =>
                           n334);
   U244 : HS65_LH_MX41X7 port map( D0 => n89, S0 => n35, D1 => n90, S1 => n33, 
                           D2 => n300, S2 => n28, D3 => n517, S3 => n24, Z => 
                           n133_port);
   U245 : HS65_LH_MX41X7 port map( D0 => n35, S0 => n518, D1 => n520, S1 => n33
                           , D2 => n521, S2 => n28, D3 => n522, S3 => n24, Z =>
                           n132_port);
   U246 : HS65_LH_MX41X7 port map( D0 => n521, S0 => n36, D1 => n520, S1 => n32
                           , D2 => n26, S2 => n518, D3 => n517, S3 => n21, Z =>
                           n231);
   U247 : HS65_LH_MX41X7 port map( D0 => n521, S0 => n37, D1 => n522, S1 => n33
                           , D2 => n523, S2 => n28, D3 => n524, S3 => n23, Z =>
                           n335);
   U248 : HS65_LH_MX41X7 port map( D0 => n82, S0 => n37, D1 => n31, S1 => n81, 
                           D2 => n80, S2 => n28, D3 => n79, S3 => n23, Z => 
                           n337);
   U249 : HS65_LH_MX41X7 port map( D0 => n520, S0 => n36, D1 => n521, S1 => n32
                           , D2 => n522, S2 => n27, D3 => n523, S3 => n22, Z =>
                           n119_port);
   U250 : HS65_LH_MX41X7 port map( D0 => n520, S0 => n36, D1 => n31, S1 => n518
                           , D2 => n517, S2 => n26, D3 => n300, S3 => n21, Z =>
                           n256);
   U251 : HS65_LH_MX41X7 port map( D0 => n35, S0 => n81, D1 => n80, S1 => n32, 
                           D2 => n79, S2 => n27, D3 => n78, S3 => n22, Z => 
                           n305);
   U252 : HS65_LH_MX41X7 port map( D0 => n83, S0 => n37, D1 => n82, S1 => n33, 
                           D2 => n26, S2 => n81, D3 => n80, S3 => n22, Z => 
                           n327);
   U253 : HS65_LH_MX41X7 port map( D0 => n75, S0 => n37, D1 => n73, S1 => n32, 
                           D2 => n71, S2 => n27, D3 => n70, S3 => n22, Z => 
                           n314);
   U254 : HS65_LH_MX41X7 port map( D0 => n90, S0 => n36, D1 => n300, S1 => n32,
                           D2 => n517, S2 => n27, D3 => n518, S3 => n22, Z => 
                           n120_port);
   U255 : HS65_LH_MX41X7 port map( D0 => n196_port, S0 => n300, D1 => n31, S1 
                           => n517, D2 => n26, S2 => n518, D3 => n520, S3 => 
                           n23, Z => n156_port);
   U256 : HS65_LH_MX41X7 port map( D0 => n80, S0 => n37, D1 => n31, S1 => n81, 
                           D2 => n82, S2 => n28, D3 => n83, S3 => n24, Z => 
                           n128_port);
   U257 : HS65_LH_MX41X7 port map( D0 => n522, S0 => n36, D1 => n521, S1 => n31
                           , D2 => n520, S2 => n26, D3 => n518, S3 => n21, Z =>
                           n214_port);
   U258 : HS65_LH_MX41X7 port map( D0 => n79, S0 => n36, D1 => n80, S1 => n31, 
                           D2 => n26, S2 => n81, D3 => n82, S3 => n20, Z => 
                           n140_port);
   U259 : HS65_LH_AO22X9 port map( A => n35, B => n70, C => n31, D => n69, Z =>
                           n303);
   U260 : HS65_LH_AO22X9 port map( A => n35, B => n531, C => n31, D => n532, Z 
                           => n222_port);
   U261 : HS65_LH_MX41X7 port map( D0 => n526, S0 => n37, D1 => n528, S1 => n33
                           , D2 => n530, S2 => n28, D3 => n531, S3 => n23, Z =>
                           n324);
   U262 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n133_port, D1 => n7, S1 => 
                           n132_port, D2 => n304, S2 => n313, D3 => n374, S3 =>
                           n263, Z => n387);
   U263 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n120_port, D1 => n7, S1 => 
                           n119_port, D2 => n304, S2 => n299, D3 => n374, S3 =>
                           n247, Z => n360);
   U264 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n156_port, D1 => n301, S1 
                           => n335, D2 => n304, S2 => n334, D3 => n374, S3 => 
                           n222_port, Z => n239);
   U265 : HS65_LH_MX41X7 port map( D0 => n75, S0 => n196_port, D1 => n77, S1 =>
                           n31, D2 => n78, S2 => n26, D3 => n79, S3 => n20, Z 
                           => n173_port);
   U266 : HS65_LH_MX41X7 port map( D0 => n77, S0 => n36, D1 => n78, S1 => n32, 
                           D2 => n79, S2 => n27, D3 => n80, S3 => n21, Z => 
                           n164_port);
   U267 : HS65_LH_MX41X7 port map( D0 => n78, S0 => n36, D1 => n79, S1 => n31, 
                           D2 => n80, S2 => n26, D3 => n20, S3 => n81, Z => 
                           n152_port);
   U268 : HS65_LH_OAI21X3 port map( A => n205_port, B => n533, C => n206_port, 
                           Z => n204_port);
   U269 : HS65_LH_AOI212X4 port map( A => n56, B => n562, C => alu_i(73), D => 
                           n180_port, E => n207_port, Z => n205_port);
   U270 : HS65_LH_CBI4I1X5 port map( A => n56, B => n533, C => n42, D => 
                           alu_i(73), Z => n206_port);
   U271 : HS65_LH_OAI211X5 port map( A => n38, B => n208_port, C => n101_port, 
                           D => n39, Z => n207_port);
   U272 : HS65_LH_AO222X4 port map( A => n313, B => n7, C => n263, D => n304, E
                           => n132_port, F => n16, Z => n174_port);
   U273 : HS65_LH_AO222X4 port map( A => n326, B => n301, C => n188_port, D => 
                           n304, E => n327, F => n16, Z => n276);
   U274 : HS65_LH_AO222X4 port map( A => n314, B => n7, C => n304, D => n315, E
                           => n316, F => n17, Z => n129_port);
   U275 : HS65_LH_AO222X4 port map( A => n302, B => n301, C => n303, D => n304,
                           E => n305, F => n17, Z => n112_port);
   U276 : HS65_LH_AO222X4 port map( A => n336, B => n301, C => n592, D => n304,
                           E => n337, F => n16, Z => n290);
   U277 : HS65_LH_MX41X7 port map( D0 => n523, S0 => n196_port, D1 => n522, S1 
                           => n32, D2 => n521, S2 => n26, D3 => n520, S3 => n20
                           , Z => n269);
   U278 : HS65_LH_AO222X4 port map( A => n324, B => n301, C => n304, D => 
                           n216_port, E => n325, F => n17, Z => n143_port);
   U279 : HS65_LH_AO222X4 port map( A => n299, B => n301, C => n247, D => n304,
                           E => n119_port, F => n16, Z => n166_port);
   U280 : HS65_LH_AO222X4 port map( A => n334, B => n7, C => n222_port, D => 
                           n304, E => n335, F => n17, Z => n155_port);
   U281 : HS65_LH_MX41X7 port map( D0 => n525, S0 => n196_port, D1 => n524, S1 
                           => n31, D2 => n523, S2 => n26, D3 => n522, S3 => n20
                           , Z => n226_port);
   U282 : HS65_LH_MX41X7 port map( D0 => n526, S0 => n196_port, D1 => n525, S1 
                           => n31, D2 => n524, S2 => n26, D3 => n523, S3 => n20
                           , Z => n209_port);
   U283 : HS65_LH_MX41X7 port map( D0 => n524, S0 => n36, D1 => n523, S1 => n31
                           , D2 => n522, S2 => n26, D3 => n521, S3 => n21, Z =>
                           n251);
   U284 : HS65_LH_OAI21X3 port map( A => n77, B => n97, C => n123_port, Z => 
                           n168_port);
   U285 : HS65_LH_OAI21X3 port map( A => n79, B => n97, C => n40, Z => 
                           n147_port);
   U286 : HS65_LH_OAI21X3 port map( A => n85, B => n54, C => n40, Z => n416);
   U287 : HS65_LH_OAI21X3 port map( A => n86, B => n54, C => n40, Z => n410);
   U288 : HS65_LH_OAI21X3 port map( A => n88, B => n54, C => n40, Z => n398);
   U289 : HS65_LH_OAI21X3 port map( A => n90, B => n97, C => n123_port, Z => 
                           n382);
   U290 : HS65_LH_OAI21X3 port map( A => n517, B => n97, C => n123_port, Z => 
                           n369);
   U291 : HS65_LH_OAI21X3 port map( A => n523, B => n97, C => n123_port, Z => 
                           n319);
   U292 : HS65_LH_OAI21X3 port map( A => n524, B => n97, C => n123_port, Z => 
                           n308);
   U293 : HS65_LH_OAI21X3 port map( A => n525, B => n97, C => n123_port, Z => 
                           n294);
   U294 : HS65_LH_OAI21X3 port map( A => n520, B => n55, C => n123_port, Z => 
                           n345);
   U295 : HS65_LH_OAI21X3 port map( A => n521, B => n55, C => n123_port, Z => 
                           n339);
   U296 : HS65_LH_OAI21X3 port map( A => n522, B => n55, C => n123_port, Z => 
                           n329);
   U297 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n306, D1 => n301, S1 => 
                           n305, D2 => n304, S2 => n302, D3 => n374, S3 => n303
                           , Z => n252);
   U298 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n292, D1 => n7, S1 => n337,
                           D2 => n304, S2 => n336, D3 => n374, S3 => n592, Z =>
                           n227);
   U299 : HS65_LH_MX41X7 port map( D0 => n16, S0 => n278, D1 => n301, S1 => 
                           n327, D2 => n304, S2 => n326, D3 => n374, S3 => 
                           n188_port, Z => n210_port);
   U300 : HS65_LH_OAI21X3 port map( A => n81, B => n97, C => n40, Z => 
                           n122_port);
   U301 : HS65_LH_OAI21X3 port map( A => n300, B => n97, C => n123_port, Z => 
                           n376);
   U302 : HS65_LH_IVX9 port map( A => alu_i(73), Z => n562);
   U303 : HS65_LH_AO22X9 port map( A => n302, B => n16, C => n303, D => n301, Z
                           => n165_port);
   U304 : HS65_LH_AO22X9 port map( A => n326, B => n16, C => n188_port, D => 
                           n301, Z => n141_port);
   U305 : HS65_LH_AO22X9 port map( A => n336, B => n16, C => n592, D => n7, Z 
                           => n153_port);
   U306 : HS65_LH_IVX9 port map( A => alu_i(70), Z => n566);
   U307 : HS65_LH_AO22X9 port map( A => n299, B => n16, C => n247, D => n301, Z
                           => n116_port);
   U308 : HS65_LH_AO22X9 port map( A => n313, B => n16, C => n263, D => n7, Z 
                           => n131_port);
   U309 : HS65_LH_AO22X9 port map( A => n334, B => n16, C => n222_port, D => n7
                           , Z => n291);
   U310 : HS65_LH_OAI212X5 port map( A => alu_i(66), B => n54, C => n14, D => 
                           n569, E => n41, Z => n318);
   U311 : HS65_LH_IVX9 port map( A => alu_i(66), Z => n569);
   U312 : HS65_LH_OAI212X5 port map( A => alu_i(63), B => n55, C => n15, D => 
                           n573, E => n41, Z => n344);
   U313 : HS65_LH_IVX9 port map( A => alu_i(63), Z => n573);
   U314 : HS65_LH_IVX9 port map( A => n190_port, Z => n563);
   U315 : HS65_LH_OAI212X5 port map( A => alu_i(60), B => n55, C => n15, D => 
                           n576, E => n40, Z => n375);
   U316 : HS65_LH_IVX9 port map( A => alu_i(60), Z => n576);
   U317 : HS65_LH_IVX9 port map( A => n264, Z => n583);
   U318 : HS65_LH_OAI212X5 port map( A => alu_i(48), B => n54, C => n14, D => 
                           n588, E => n41, Z => n158_port);
   U319 : HS65_LH_IVX9 port map( A => alu_i(48), Z => n588);
   U320 : HS65_LH_OAI212X5 port map( A => alu_i(42), B => n97, C => n14, D => 
                           n594, E => n441, Z => n439);
   U321 : HS65_LH_AOI12X2 port map( A => n599, B => n196_port, C => n42, Z => 
                           n441);
   U322 : HS65_LH_OAI212X5 port map( A => alu_i(72), B => n54, C => n14, D => 
                           n565, E => n41, Z => n223_port);
   U323 : HS65_LH_OAI212X5 port map( A => alu_i(43), B => n55, C => n15, D => 
                           n593, E => n41, Z => n357);
   U324 : HS65_LH_CBI4I6X5 port map( A => n531, B => n54, C => n40, D => n565, 
                           Z => n224_port);
   U325 : HS65_LH_CBI4I6X5 port map( A => n69, B => n54, C => n40, D => n594, Z
                           => n440);
   U326 : HS65_LH_CBI4I6X5 port map( A => n70, B => n54, C => n40, D => n593, Z
                           => n358);
   U327 : HS65_LH_IVX9 port map( A => alu_i(72), Z => n565);
   U328 : HS65_LH_OAI21X3 port map( A => n78, B => n97, C => n40, Z => 
                           n159_port);
   U329 : HS65_LH_OAI21X3 port map( A => n80, B => n54, C => n40, Z => 
                           n135_port);
   U330 : HS65_LH_OAI21X3 port map( A => n82, B => n97, C => n40, Z => n429);
   U331 : HS65_LH_OAI21X3 port map( A => n87, B => n54, C => n40, Z => n404);
   U332 : HS65_LH_OAI21X3 port map( A => n89, B => n97, C => n123_port, Z => 
                           n389);
   U333 : HS65_LH_IVX9 port map( A => alu_i(42), Z => n594);
   U334 : HS65_LH_IVX9 port map( A => alu_i(43), Z => n593);
   U335 : HS65_LH_IVX9 port map( A => alu_i(45), Z => n590);
   U336 : HS65_LH_NOR3X4 port map( A => alu_i(7), B => alu_i(9), C => n607, Z 
                           => n434);
   U337 : HS65_LH_BFX9 port map( A => n104_port, Z => n46);
   U338 : HS65_LH_OAI21X3 port map( A => alu_i(5), B => n437, C => n443, Z => 
                           n104_port);
   U339 : HS65_LH_OAI21X3 port map( A => n436, B => n435, C => n390, Z => n443)
                           ;
   U340 : HS65_LH_NOR2X6 port map( A => n596, B => n96, Z => n275);
   U341 : HS65_LH_NAND2X7 port map( A => n7, B => n596, Z => n189_port);
   U342 : HS65_LH_NOR2X6 port map( A => n602, B => n601, Z => n374);
   U343 : HS65_LH_NOR2X6 port map( A => n596, B => n98, Z => n117_port);
   U344 : HS65_LH_NOR2X6 port map( A => n609, B => alu_i(6), Z => n391);
   U345 : HS65_LH_NOR2X6 port map( A => alu_i(6), B => alu_i(5), Z => n438);
   U346 : HS65_LH_NOR2X6 port map( A => n611, B => alu_i(5), Z => n436);
   U347 : HS65_LH_AND2X4 port map( A => n192_port, B => n606, Z => n277);
   U348 : HS65_LH_NAND2X7 port map( A => n193_port, B => n605, Z => n208_port);
   U349 : HS65_LH_NAND2X7 port map( A => n193_port, B => n606, Z => n186_port);
   U350 : HS65_LH_NAND4ABX3 port map( A => alu_i(9), B => alu_i(7), C => n611, 
                           D => n607, Z => n437);
   U351 : HS65_LH_IVX9 port map( A => alu_i(5), Z => n609);
   U352 : HS65_LH_NOR2AX3 port map( A => alu_i(7), B => alu_i(9), Z => n445);
   U353 : HS65_LH_IVX9 port map( A => alu_i(9), Z => n612);
   U354 : HS65_LH_AND2X4 port map( A => n448, B => n602, Z => n195_port);
   U355 : HS65_LH_IVX9 port map( A => alu_i(8), Z => n607);
   U356 : HS65_LH_IVX9 port map( A => alu_i(6), Z => n611);
   U357 : HS65_LH_AND2X4 port map( A => n192_port, B => n605, Z => n118_port);
   U358 : HS65_LH_AND2X4 port map( A => n445, B => alu_i(8), Z => n390);
   U359 : HS65_LH_IVX9 port map( A => n35, Z => n38);
   U360 : HS65_LH_IVX9 port map( A => n6, Z => n16);
   U361 : HS65_LH_BFX9 port map( A => n199_port, Z => n18);
   U362 : HS65_LH_BFX9 port map( A => n197_port, Z => n30);
   U363 : HS65_LH_BFX9 port map( A => n197_port, Z => n29);
   U364 : HS65_LH_BFX9 port map( A => n25, Z => n26);
   U365 : HS65_LH_BFX9 port map( A => n25, Z => n28);
   U366 : HS65_LH_BFX9 port map( A => n25, Z => n27);
   U367 : HS65_LH_BFX9 port map( A => n199_port, Z => n19);
   U368 : HS65_LH_IVX9 port map( A => n6, Z => n17);
   U369 : HS65_LH_AO22X9 port map( A => N226, B => n61, C => HI_LO_c_HI_31_port
                           , D => n57, Z => n516);
   U370 : HS65_LH_IVX9 port map( A => alu_i(44), Z => n535);
   U371 : HS65_LH_IVX9 port map( A => alu_i(47), Z => n537);
   U372 : HS65_LH_IVX9 port map( A => alu_i(50), Z => n539);
   U373 : HS65_LH_IVX9 port map( A => alu_i(12), Z => n72);
   U374 : HS65_LH_BFX9 port map( A => alu_i(10), Z => n69);
   U375 : HS65_LH_AO22X9 port map( A => N224, B => n63, C => HI_LO_c_HI_29_port
                           , D => n57, Z => n514);
   U376 : HS65_LH_AO22X9 port map( A => N225, B => n62, C => HI_LO_c_HI_30_port
                           , D => n57, Z => n515);
   U377 : HS65_LH_IVX9 port map( A => alu_i(14), Z => n76);
   U378 : HS65_LH_IVX9 port map( A => alu_i(53), Z => n541);
   U379 : HS65_LH_IVX9 port map( A => alu_i(56), Z => n543);
   U380 : HS65_LH_IVX9 port map( A => alu_i(59), Z => n545);
   U381 : HS65_LH_IVX9 port map( A => alu_i(62), Z => n547);
   U382 : HS65_LH_IVX9 port map( A => alu_i(13), Z => n74);
   U383 : HS65_LH_AO22X9 port map( A => N217, B => n63, C => HI_LO_c_HI_22_port
                           , D => n57, Z => n507);
   U384 : HS65_LH_AO22X9 port map( A => N218, B => n63, C => HI_LO_c_HI_23_port
                           , D => n57, Z => n508);
   U385 : HS65_LH_AO22X9 port map( A => N219, B => n63, C => HI_LO_c_HI_24_port
                           , D => n57, Z => n509);
   U386 : HS65_LH_AO22X9 port map( A => N220, B => n63, C => HI_LO_c_HI_25_port
                           , D => n57, Z => n510);
   U387 : HS65_LH_AO22X9 port map( A => N221, B => n63, C => HI_LO_c_HI_26_port
                           , D => n57, Z => n511);
   U388 : HS65_LH_AO22X9 port map( A => N222, B => n63, C => HI_LO_c_HI_27_port
                           , D => n57, Z => n512);
   U389 : HS65_LH_AO22X9 port map( A => N223, B => n63, C => HI_LO_c_HI_28_port
                           , D => n57, Z => n513);
   U390 : HS65_LH_IVX9 port map( A => alu_i(21), Z => n84);
   U391 : HS65_LH_IVX9 port map( A => alu_i(65), Z => n549);
   U392 : HS65_LH_IVX9 port map( A => alu_i(68), Z => n551);
   U393 : HS65_LH_IVX9 port map( A => alu_i(71), Z => n553);
   U394 : HS65_LH_AO22X9 port map( A => N210, B => n63, C => HI_LO_c_HI_15_port
                           , D => n58, Z => n500);
   U395 : HS65_LH_AO22X9 port map( A => N211, B => n63, C => HI_LO_c_HI_16_port
                           , D => n58, Z => n501);
   U396 : HS65_LH_AO22X9 port map( A => N212, B => n63, C => HI_LO_c_HI_17_port
                           , D => n58, Z => n502);
   U397 : HS65_LH_AO22X9 port map( A => N213, B => n63, C => HI_LO_c_HI_18_port
                           , D => n58, Z => n503);
   U398 : HS65_LH_AO22X9 port map( A => N214, B => n63, C => HI_LO_c_HI_19_port
                           , D => n58, Z => n504);
   U399 : HS65_LH_AO22X9 port map( A => N215, B => n63, C => HI_LO_c_HI_20_port
                           , D => n57, Z => n505);
   U400 : HS65_LH_AO22X9 port map( A => N216, B => n63, C => HI_LO_c_HI_21_port
                           , D => n57, Z => n506);
   U401 : HS65_LH_IVX9 port map( A => alu_i(30), Z => n519);
   U402 : HS65_LH_AO22X9 port map( A => N204, B => n64, C => HI_LO_c_HI_9_port,
                           D => n58, Z => n494);
   U403 : HS65_LH_AO22X9 port map( A => N205, B => n63, C => HI_LO_c_HI_10_port
                           , D => n58, Z => n495);
   U404 : HS65_LH_AO22X9 port map( A => N206, B => n63, C => HI_LO_c_HI_11_port
                           , D => n58, Z => n496);
   U405 : HS65_LH_AO22X9 port map( A => N207, B => n63, C => HI_LO_c_HI_12_port
                           , D => n58, Z => n497);
   U406 : HS65_LH_AO22X9 port map( A => N208, B => n63, C => HI_LO_c_HI_13_port
                           , D => n58, Z => n498);
   U407 : HS65_LH_AO22X9 port map( A => N209, B => n63, C => HI_LO_c_HI_14_port
                           , D => n58, Z => n499);
   U408 : HS65_LH_IVX9 port map( A => alu_i(38), Z => n529);
   U409 : HS65_LH_IVX9 port map( A => alu_i(37), Z => n527);
   U410 : HS65_LH_AO22X9 port map( A => N199, B => n64, C => HI_LO_c_HI_4_port,
                           D => n58, Z => n489);
   U411 : HS65_LH_AO22X9 port map( A => N200, B => n64, C => HI_LO_c_HI_5_port,
                           D => n57, Z => n490);
   U412 : HS65_LH_AO22X9 port map( A => N201, B => n64, C => HI_LO_c_HI_6_port,
                           D => n58, Z => n491);
   U413 : HS65_LH_AO22X9 port map( A => N202, B => n64, C => HI_LO_c_HI_7_port,
                           D => n57, Z => n492);
   U414 : HS65_LH_AO22X9 port map( A => N203, B => n64, C => HI_LO_c_HI_8_port,
                           D => n58, Z => n493);
   U415 : HS65_LH_AO22X9 port map( A => N197, B => n64, C => HI_LO_c_HI_2_port,
                           D => n58, Z => n487);
   U416 : HS65_LH_AO22X9 port map( A => N198, B => n64, C => HI_LO_c_HI_3_port,
                           D => n57, Z => n488);
   U417 : HS65_LH_IVX9 port map( A => alu_i(41), Z => n533);
   U418 : HS65_LH_AO22X9 port map( A => N194, B => n64, C => HI_LO_c_LO_31_port
                           , D => n58, Z => n484);
   U419 : HS65_LH_AO22X9 port map( A => N196, B => n64, C => HI_LO_c_HI_1_port,
                           D => n57, Z => n486);
   U420 : HS65_LH_AO22X9 port map( A => N191, B => n64, C => HI_LO_c_LO_28_port
                           , D => n59, Z => n481);
   U421 : HS65_LH_AO22X9 port map( A => N192, B => n64, C => HI_LO_c_LO_29_port
                           , D => n58, Z => n482);
   U422 : HS65_LH_AO22X9 port map( A => N193, B => n64, C => HI_LO_c_LO_30_port
                           , D => n57, Z => n483);
   U423 : HS65_LH_AO22X9 port map( A => N195, B => n64, C => HI_LO_c_HI_0_port,
                           D => n60, Z => n485);
   U424 : HS65_LH_AO22X9 port map( A => N184, B => n65, C => HI_LO_c_LO_21_port
                           , D => n59, Z => n474);
   U425 : HS65_LH_AO22X9 port map( A => N185, B => n64, C => HI_LO_c_LO_22_port
                           , D => n59, Z => n475);
   U426 : HS65_LH_AO22X9 port map( A => N186, B => n64, C => HI_LO_c_LO_23_port
                           , D => n59, Z => n476);
   U427 : HS65_LH_AO22X9 port map( A => N187, B => n64, C => HI_LO_c_LO_24_port
                           , D => n59, Z => n477);
   U428 : HS65_LH_AO22X9 port map( A => N188, B => n64, C => HI_LO_c_LO_25_port
                           , D => n59, Z => n478);
   U429 : HS65_LH_AO22X9 port map( A => N189, B => n64, C => HI_LO_c_LO_26_port
                           , D => n59, Z => n479);
   U430 : HS65_LH_AO22X9 port map( A => N190, B => n64, C => HI_LO_c_LO_27_port
                           , D => n59, Z => n480);
   U431 : HS65_LH_AOI222X2 port map( A => N157, B => n51, C => n11, D => 
                           HI_LO_c_HI_26_port, E => n8, F => n526, Z => n288);
   U432 : HS65_LH_AOI222X2 port map( A => N158, B => n51, C => n11, D => 
                           HI_LO_c_HI_27_port, E => n8, F => n528, Z => n273);
   U433 : HS65_LH_AOI22X6 port map( A => N128, B => n48, C => n606, D => n250, 
                           Z => n243);
   U434 : HS65_LH_AO212X4 port map( A => n251, B => n595, C => n252, D => 
                           alu_i(4), E => n253, Z => n250);
   U435 : HS65_LH_AO222X4 port map( A => n192_port, B => n254, C => n193_port, 
                           D => n255, E => n195_port, F => n256, Z => n253);
   U436 : HS65_LH_MX41X7 port map( D0 => n530, S0 => n196_port, D1 => n528, S1 
                           => n31, D2 => n526, S2 => n26, D3 => n525, S3 => n20
                           , Z => n255);
   U437 : HS65_LH_AOI22X6 port map( A => N129, B => n48, C => n606, D => 
                           n225_port, Z => n218_port);
   U438 : HS65_LH_AO212X4 port map( A => n226_port, B => n595, C => n227, D => 
                           alu_i(4), E => n228, Z => n225_port);
   U439 : HS65_LH_AO222X4 port map( A => n192_port, B => n229, C => n193_port, 
                           D => n230, E => n195_port, F => n231, Z => n228);
   U440 : HS65_LH_MX41X7 port map( D0 => n531, S0 => n36, D1 => n530, S1 => n31
                           , D2 => n528, S2 => n26, D3 => n526, S3 => n20, Z =>
                           n230);
   U441 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_25_port, D1 => 
                           n106_port, S1 => n81, D2 => N124, S2 => n48, D3 => 
                           n599, S3 => n251, Z => n295);
   U442 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_26_port, D1 => 
                           n106_port, S1 => n82, D2 => N125, S2 => n48, D3 => 
                           n599, S3 => n226_port, Z => n286);
   U443 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_27_port, D1 => 
                           n106_port, S1 => n83, D2 => N126, S2 => n48, D3 => 
                           n599, S3 => n209_port, Z => n271);
   U444 : HS65_LH_AO22X9 port map( A => N177, B => n65, C => HI_LO_c_LO_14_port
                           , D => n60, Z => n467);
   U445 : HS65_LH_AO22X9 port map( A => N178, B => n65, C => HI_LO_c_LO_15_port
                           , D => n60, Z => n468);
   U446 : HS65_LH_AO22X9 port map( A => N179, B => n65, C => HI_LO_c_LO_16_port
                           , D => n59, Z => n469);
   U447 : HS65_LH_AO22X9 port map( A => N180, B => n65, C => HI_LO_c_LO_17_port
                           , D => n59, Z => n470);
   U448 : HS65_LH_AO22X9 port map( A => N181, B => n65, C => HI_LO_c_LO_18_port
                           , D => n59, Z => n471);
   U449 : HS65_LH_AO22X9 port map( A => N182, B => n65, C => HI_LO_c_LO_19_port
                           , D => n59, Z => n472);
   U450 : HS65_LH_AO22X9 port map( A => N183, B => n65, C => HI_LO_c_LO_20_port
                           , D => n59, Z => n473);
   U451 : HS65_LH_NAND4ABX3 port map( A => n295, B => n296, C => n297, D => 
                           n298, Z => alu_o(25));
   U452 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n306, D1 => n598, S1 => 
                           n254, D2 => n524, S2 => n307, D3 => alu_i(67), S3 =>
                           n308, Z => n296);
   U453 : HS65_LH_AOI222X2 port map( A => n275, B => n112_port, C => n279, D =>
                           n256, E => n284, F => n116_port, Z => n298);
   U454 : HS65_LH_NAND4ABX3 port map( A => n286, B => n287, C => n288, D => 
                           n289, Z => alu_o(26));
   U455 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n292, D1 => n598, S1 => 
                           n229, D2 => n525, S2 => n293, D3 => n550, S3 => n294
                           , Z => n287);
   U456 : HS65_LH_AOI222X2 port map( A => n275, B => n290, C => n279, D => n231
                           , E => n284, F => n291, Z => n289);
   U457 : HS65_LH_NAND4ABX3 port map( A => n271, B => n272, C => n273, D => 
                           n274, Z => alu_o(27));
   U458 : HS65_LH_AOI222X2 port map( A => n275, B => n276, C => n277, D => n278
                           , E => n279, F => n214_port, Z => n274);
   U459 : HS65_LH_OAI212X5 port map( A => n280, B => n527, C => n575, D => n281
                           , E => n282, Z => n272);
   U460 : HS65_LH_NAND3X5 port map( A => n243, B => n244, C => n245, Z => 
                           alu_o(29));
   U461 : HS65_LH_AOI212X4 port map( A => n600, B => n247, C => n530, D => n248
                           , E => n249, Z => n244);
   U462 : HS65_LH_AOI212X4 port map( A => n10, B => n531, C => N160, D => n53, 
                           E => n246, Z => n245);
   U463 : HS65_LH_NAND3X5 port map( A => n218_port, B => n219_port, C => 
                           n220_port, Z => alu_o(30));
   U464 : HS65_LH_AOI212X4 port map( A => n600, B => n222_port, C => n531, D =>
                           n223_port, E => n224_port, Z => n219_port);
   U465 : HS65_LH_AOI212X4 port map( A => n10, B => n532, C => N161, D => n53, 
                           E => n221_port, Z => n220_port);
   U466 : HS65_LH_NAND2X7 port map( A => n257, B => n258, Z => alu_o(28));
   U467 : HS65_LH_AOI212X4 port map( A => n9, B => n530, C => N159, D => n53, E
                           => n270, Z => n257);
   U468 : HS65_LH_AOI212X4 port map( A => N127, B => n48, C => n606, D => n259,
                           E => n260, Z => n258);
   U469 : HS65_LH_NAND2X7 port map( A => n201_port, B => n202_port, Z => 
                           alu_o(31));
   U470 : HS65_LH_AOI212X4 port map( A => n13, B => HI_LO_c_HI_31_port, C => 
                           N162, D => n53, E => n217_port, Z => n201_port);
   U471 : HS65_LH_AOI212X4 port map( A => N130, B => n48, C => n606, D => 
                           n203_port, E => n204_port, Z => n202_port);
   U472 : HS65_LH_AOI222X2 port map( A => N152, B => n52, C => n11, D => 
                           HI_LO_c_HI_21_port, E => n8, F => n521, Z => n342);
   U473 : HS65_LH_AOI222X2 port map( A => N153, B => n51, C => n11, D => 
                           HI_LO_c_HI_22_port, E => n8, F => n522, Z => n332);
   U474 : HS65_LH_AOI222X2 port map( A => N154, B => n51, C => n11, D => 
                           HI_LO_c_HI_23_port, E => n8, F => n523, Z => n322);
   U475 : HS65_LH_AOI222X2 port map( A => N155, B => n51, C => n11, D => 
                           HI_LO_c_HI_24_port, E => n8, F => n524, Z => n311);
   U476 : HS65_LH_AOI222X2 port map( A => N156, B => n51, C => n11, D => 
                           HI_LO_c_HI_25_port, E => n8, F => n525, Z => n297);
   U477 : HS65_LH_AOI222X2 port map( A => N149, B => n52, C => n12, D => 
                           HI_LO_c_HI_18_port, E => n9, F => n517, Z => n372);
   U478 : HS65_LH_AOI222X2 port map( A => N150, B => n52, C => n12, D => 
                           HI_LO_c_HI_19_port, E => n9, F => n518, Z => n365);
   U479 : HS65_LH_AOI222X2 port map( A => N151, B => n52, C => n12, D => 
                           HI_LO_c_HI_20_port, E => n9, F => n520, Z => n348);
   U480 : HS65_LH_AOI212X4 port map( A => n10, B => n70, C => N131, D => n53, E
                           => n433, Z => n432);
   U481 : HS65_LH_AO222X4 port map( A => N649, B => n103_port, C => n13, D => 
                           HI_LO_c_HI_0_port, E => N648, F => n102_port, Z => 
                           n433);
   U482 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_17_port, D1 => 
                           n106_port, S1 => n70, D2 => N116, S2 => n49, D3 => 
                           n599, S3 => n254, Z => n377);
   U483 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_18_port, D1 => 
                           n106_port, S1 => n71, D2 => N117, S2 => n49, D3 => 
                           n599, S3 => n229, Z => n370);
   U484 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_19_port, D1 => 
                           n106_port, S1 => n73, D2 => N118, S2 => n48, D3 => 
                           n599, S3 => n212_port, Z => n363);
   U485 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_20_port, D1 => 
                           n106_port, S1 => n75, D2 => N119, S2 => n48, D3 => 
                           n599, S3 => n268, Z => n346);
   U486 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_21_port, D1 => 
                           n106_port, S1 => n77, D2 => N120, S2 => n48, D3 => 
                           n599, S3 => n256, Z => n340);
   U487 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_22_port, D1 => 
                           n106_port, S1 => n78, D2 => N121, S2 => n48, D3 => 
                           n599, S3 => n231, Z => n330);
   U488 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_23_port, D1 => 
                           n106_port, S1 => n79, D2 => N122, S2 => n48, D3 => 
                           n599, S3 => n214_port, Z => n320);
   U489 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_24_port, D1 => 
                           n106_port, S1 => n80, D2 => N123, S2 => n48, D3 => 
                           n599, S3 => n269, Z => n309);
   U490 : HS65_LH_AO22X9 port map( A => N171, B => n65, C => HI_LO_c_LO_8_port,
                           D => n60, Z => n461);
   U491 : HS65_LH_AO22X9 port map( A => N172, B => n65, C => HI_LO_c_LO_9_port,
                           D => n60, Z => n462);
   U492 : HS65_LH_AO22X9 port map( A => N173, B => n65, C => HI_LO_c_LO_10_port
                           , D => n60, Z => n463);
   U493 : HS65_LH_AO22X9 port map( A => N174, B => n65, C => HI_LO_c_LO_11_port
                           , D => n60, Z => n464);
   U494 : HS65_LH_AO22X9 port map( A => N175, B => n65, C => HI_LO_c_LO_12_port
                           , D => n60, Z => n465);
   U495 : HS65_LH_AO22X9 port map( A => N176, B => n65, C => HI_LO_c_LO_13_port
                           , D => n60, Z => n466);
   U496 : HS65_LH_NAND4ABX3 port map( A => n340, B => n341, C => n342, D => 
                           n343, Z => alu_o(21));
   U497 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n305, D1 => n598, S1 => 
                           n306, D2 => n520, S2 => n344, D3 => alu_i(63), S3 =>
                           n345, Z => n341);
   U498 : HS65_LH_AOI222X2 port map( A => n275, B => n165_port, C => n279, D =>
                           n254, E => n284, F => n166_port, Z => n343);
   U499 : HS65_LH_NAND4ABX3 port map( A => n330, B => n331, C => n332, D => 
                           n333, Z => alu_o(22));
   U500 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n337, D1 => n598, S1 => 
                           n292, D2 => n521, S2 => n338, D3 => alu_i(64), S3 =>
                           n339, Z => n331);
   U501 : HS65_LH_AOI222X2 port map( A => n275, B => n153_port, C => n279, D =>
                           n229, E => n284, F => n155_port, Z => n333);
   U502 : HS65_LH_NAND4ABX3 port map( A => n320, B => n321, C => n322, D => 
                           n323, Z => alu_o(23));
   U503 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n327, D1 => n598, S1 => 
                           n278, D2 => n522, S2 => n328, D3 => n548, S3 => n329
                           , Z => n321);
   U504 : HS65_LH_AOI222X2 port map( A => n275, B => n141_port, C => n279, D =>
                           n212_port, E => n284, F => n143_port, Z => n323);
   U505 : HS65_LH_NAND4ABX3 port map( A => n309, B => n310, C => n311, D => 
                           n312, Z => alu_o(24));
   U506 : HS65_LH_MX41X7 port map( D0 => n277, S0 => n317, D1 => n598, S1 => 
                           n266, D2 => n523, S2 => n318, D3 => alu_i(66), S3 =>
                           n319, Z => n310);
   U507 : HS65_LH_AOI222X2 port map( A => n275, B => n129_port, C => n279, D =>
                           n268, E => n284, F => n131_port, Z => n312);
   U508 : HS65_LH_NAND4ABX3 port map( A => n377, B => n378, C => n379, D => 
                           n380, Z => alu_o(17));
   U509 : HS65_LH_MX41X7 port map( D0 => n598, S0 => n305, D1 => n90, S1 => 
                           n381, D2 => n368, S2 => n303, D3 => n544, S3 => n382
                           , Z => n378);
   U510 : HS65_LH_AOI222X2 port map( A => n284, B => n360, C => n277, D => n302
                           , E => n279, F => n306, Z => n380);
   U511 : HS65_LH_NAND4ABX3 port map( A => n370, B => n371, C => n372, D => 
                           n373, Z => alu_o(18));
   U512 : HS65_LH_MX41X7 port map( D0 => n598, S0 => n337, D1 => n300, S1 => 
                           n375, D2 => n368, S2 => n592, D3 => alu_i(60), S3 =>
                           n376, Z => n371);
   U513 : HS65_LH_AOI222X2 port map( A => n284, B => n239, C => n277, D => n336
                           , E => n279, F => n292, Z => n373);
   U514 : HS65_LH_NAND4ABX3 port map( A => n363, B => n364, C => n365, D => 
                           n366, Z => alu_o(19));
   U515 : HS65_LH_MX41X7 port map( D0 => n598, S0 => n327, D1 => n517, S1 => 
                           n367, D2 => n368, S2 => n188_port, D3 => alu_i(61), 
                           S3 => n369, Z => n364);
   U516 : HS65_LH_AOI222X2 port map( A => n284, B => n563, C => n277, D => n326
                           , E => n279, F => n278, Z => n366);
   U517 : HS65_LH_NAND4ABX3 port map( A => n346, B => n347, C => n348, D => 
                           n349, Z => alu_o(20));
   U518 : HS65_LH_AOI222X2 port map( A => n284, B => n174_port, C => n277, D =>
                           n316, E => n279, F => n266, Z => n349);
   U519 : HS65_LH_OAI212X5 port map( A => n350, B => n519, C => n582, D => n281
                           , E => n351, Z => n347);
   U520 : HS65_LH_NAND3X5 port map( A => n430, B => n431, C => n432, Z => 
                           alu_o(0));
   U521 : HS65_LH_AOI212X4 port map( A => N99, B => n48, C => n69, D => n439, E
                           => n440, Z => n431);
   U522 : HS65_LH_AOI22X6 port map( A => n605, B => n444, C => n45, D => 
                           HI_LO_c_LO_0_port, Z => n430);
   U523 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_9_port, C => 
                           n600, D => n111_port, E => N108, F => n47, Z => 
                           n110_port);
   U524 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_10_port, C => 
                           n600, D => n154_port, E => N109, F => n47, Z => n427
                           );
   U525 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_11_port, C => 
                           n600, D => n142_port, E => N110, F => n47, Z => n420
                           );
   U526 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_12_port, C => 
                           n600, D => n130_port, E => N111, F => n47, Z => n414
                           );
   U527 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_13_port, C => 
                           n600, D => n114_port, E => N112, F => n47, Z => n408
                           );
   U528 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_14_port, C => 
                           n600, D => n157_port, E => N113, F => n47, Z => n402
                           );
   U529 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_15_port, C => 
                           n600, D => n145_port, E => N114, F => n47, Z => n395
                           );
   U530 : HS65_LH_AOI222X2 port map( A => N140, B => n51, C => n11, D => 
                           HI_LO_c_HI_9_port, E => n8, F => n82, Z => n109_port
                           );
   U531 : HS65_LH_AOI222X2 port map( A => N141, B => n52, C => n12, D => 
                           HI_LO_c_HI_10_port, E => n9, F => n83, Z => n426);
   U532 : HS65_LH_AOI222X2 port map( A => N142, B => n52, C => n12, D => 
                           HI_LO_c_HI_11_port, E => n9, F => n85, Z => n419);
   U533 : HS65_LH_AOI222X2 port map( A => N143, B => n52, C => n12, D => 
                           HI_LO_c_HI_12_port, E => n9, F => n86, Z => n413);
   U534 : HS65_LH_AOI222X2 port map( A => N144, B => n52, C => n12, D => 
                           HI_LO_c_HI_13_port, E => n9, F => n87, Z => n407);
   U535 : HS65_LH_AOI222X2 port map( A => N145, B => n52, C => n12, D => 
                           HI_LO_c_HI_14_port, E => n9, F => n88, Z => n401);
   U536 : HS65_LH_AOI222X2 port map( A => N146, B => n52, C => n12, D => 
                           HI_LO_c_HI_15_port, E => n9, F => n89, Z => n394);
   U537 : HS65_LH_AOI222X2 port map( A => N147, B => n52, C => n12, D => 
                           HI_LO_c_HI_16_port, E => n9, F => n90, Z => n385);
   U538 : HS65_LH_AOI222X2 port map( A => N148, B => n52, C => n12, D => 
                           HI_LO_c_HI_17_port, E => n9, F => n300, Z => n379);
   U539 : HS65_LH_MX41X7 port map( D0 => n45, S0 => HI_LO_c_LO_16_port, D1 => 
                           n106_port, S1 => n69, D2 => N115, S2 => n49, D3 => 
                           n599, S3 => n266, Z => n383);
   U540 : HS65_LH_AO22X9 port map( A => N167, B => n65, C => HI_LO_c_LO_4_port,
                           D => n60, Z => n457);
   U541 : HS65_LH_AO22X9 port map( A => N168, B => n65, C => HI_LO_c_LO_5_port,
                           D => n60, Z => n458);
   U542 : HS65_LH_AO22X9 port map( A => N169, B => n65, C => HI_LO_c_LO_6_port,
                           D => n60, Z => n459);
   U543 : HS65_LH_AO22X9 port map( A => N170, B => n65, C => HI_LO_c_LO_7_port,
                           D => n60, Z => n460);
   U544 : HS65_LH_AO22X9 port map( A => N163, B => n66, C => HI_LO_c_LO_0_port,
                           D => n60, Z => n453);
   U545 : HS65_LH_AO22X9 port map( A => N164, B => n66, C => HI_LO_c_LO_1_port,
                           D => n59, Z => n454);
   U546 : HS65_LH_AO22X9 port map( A => N165, B => n65, C => HI_LO_c_LO_2_port,
                           D => n60, Z => n455);
   U547 : HS65_LH_AO22X9 port map( A => N166, B => n65, C => HI_LO_c_LO_3_port,
                           D => n59, Z => n456);
   U548 : HS65_LH_NAND4ABX3 port map( A => n383, B => n384, C => n385, D => 
                           n386, Z => alu_o(16));
   U549 : HS65_LH_MX41X7 port map( D0 => n598, S0 => n316, D1 => n89, S1 => 
                           n388, D2 => n368, S2 => n315, D3 => alu_i(58), S3 =>
                           n389, Z => n384);
   U550 : HS65_LH_AOI222X2 port map( A => n284, B => n387, C => n277, D => n314
                           , E => n279, F => n317, Z => n386);
   U551 : HS65_LH_NAND4ABX3 port map( A => n107_port, B => n108_port, C => 
                           n109_port, D => n110_port, Z => alu_o(9));
   U552 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n119_port, D1 => n597
                           , S1 => n120_port, D2 => n81, S2 => n121_port, D3 =>
                           alu_i(51), S3 => n122_port, Z => n107_port);
   U553 : HS65_LH_AO222X4 port map( A => n112_port, B => n113_port, C => 
                           n114_port, D => n115_port, E => n116_port, F => 
                           n117_port, Z => n108_port);
   U554 : HS65_LH_NAND4ABX3 port map( A => n424, B => n425, C => n426, D => 
                           n427, Z => alu_o(10));
   U555 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n335, D1 => n597, S1 
                           => n156_port, D2 => n82, S2 => n428, D3 => alu_i(52)
                           , S3 => n429, Z => n424);
   U556 : HS65_LH_AO222X4 port map( A => n290, B => n113_port, C => n157_port, 
                           D => n115_port, E => n291, F => n117_port, Z => n425
                           );
   U557 : HS65_LH_NAND4ABX3 port map( A => n417, B => n418, C => n419, D => 
                           n420, Z => alu_o(11));
   U558 : HS65_LH_OAI212X5 port map( A => n421, B => n84, C => n572, D => 
                           n176_port, E => n422, Z => n417);
   U559 : HS65_LH_AO222X4 port map( A => n145_port, B => n115_port, C => n325, 
                           D => n118_port, E => n276, F => n113_port, Z => n418
                           );
   U560 : HS65_LH_NAND4ABX3 port map( A => n411, B => n412, C => n413, D => 
                           n414, Z => alu_o(12));
   U561 : HS65_LH_MX41X7 port map( D0 => n597, S0 => n132_port, D1 => n85, S1 
                           => n415, D2 => n397, S2 => n263, D3 => alu_i(54), S3
                           => n416, Z => n411);
   U562 : HS65_LH_AO222X4 port map( A => n133_port, B => n115_port, C => n313, 
                           D => n118_port, E => n583, F => n113_port, Z => n412
                           );
   U563 : HS65_LH_NAND4ABX3 port map( A => n405, B => n406, C => n407, D => 
                           n408, Z => alu_o(13));
   U564 : HS65_LH_MX41X7 port map( D0 => n597, S0 => n119_port, D1 => n86, S1 
                           => n409, D2 => n397, S2 => n247, D3 => alu_i(55), S3
                           => n410, Z => n405);
   U565 : HS65_LH_AO222X4 port map( A => n120_port, B => n115_port, C => n299, 
                           D => n118_port, E => n252, F => n113_port, Z => n406
                           );
   U566 : HS65_LH_NAND4ABX3 port map( A => n399, B => n400, C => n401, D => 
                           n402, Z => alu_o(14));
   U567 : HS65_LH_MX41X7 port map( D0 => n597, S0 => n335, D1 => n87, S1 => 
                           n403, D2 => n397, S2 => n222_port, D3 => n542, S3 =>
                           n404, Z => n399);
   U568 : HS65_LH_AO222X4 port map( A => n156_port, B => n115_port, C => n334, 
                           D => n118_port, E => n227, F => n113_port, Z => n400
                           );
   U569 : HS65_LH_NAND4ABX3 port map( A => n392, B => n393, C => n394, D => 
                           n395, Z => alu_o(15));
   U570 : HS65_LH_MX41X7 port map( D0 => n597, S0 => n325, D1 => n88, S1 => 
                           n396, D2 => n397, S2 => n216_port, D3 => alu_i(57), 
                           S3 => n398, Z => n392);
   U571 : HS65_LH_AO222X4 port map( A => n144_port, B => n115_port, C => n324, 
                           D => n118_port, E => n210_port, F => n113_port, Z =>
                           n393);
   U572 : HS65_LH_AOI222X2 port map( A => n317, B => n16, C => n316, D => n301,
                           E => n178_port, F => alu_i(3), Z => n264);
   U573 : HS65_LH_AOI222X2 port map( A => n144_port, B => n16, C => n325, D => 
                           n7, E => n283, F => alu_i(3), Z => n190_port);
   U574 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_5_port, C => 
                           n600, D => n164_port, E => N104, F => n47, Z => 
                           n163_port);
   U575 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_6_port, C => 
                           n600, D => n152_port, E => N105, F => n47, Z => 
                           n151_port);
   U576 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_7_port, C => 
                           n600, D => n140_port, E => N106, F => n47, Z => 
                           n139_port);
   U577 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_8_port, C => 
                           n600, D => n128_port, E => N107, F => n47, Z => 
                           n127_port);
   U578 : HS65_LH_AOI222X2 port map( A => N135, B => n51, C => n11, D => 
                           HI_LO_c_HI_4_port, E => n8, F => n77, Z => n171_port
                           );
   U579 : HS65_LH_AOI222X2 port map( A => N136, B => n51, C => n12, D => 
                           HI_LO_c_HI_5_port, E => n8, F => n78, Z => n162_port
                           );
   U580 : HS65_LH_AOI222X2 port map( A => N137, B => n51, C => n11, D => 
                           HI_LO_c_HI_6_port, E => n8, F => n79, Z => n150_port
                           );
   U581 : HS65_LH_AOI222X2 port map( A => N138, B => n51, C => n11, D => 
                           HI_LO_c_HI_7_port, E => n8, F => n80, Z => n138_port
                           );
   U582 : HS65_LH_AOI222X2 port map( A => N139, B => n51, C => n11, D => 
                           HI_LO_c_HI_8_port, E => n8, F => n81, Z => n126_port
                           );
   U583 : HS65_LH_AOI22X6 port map( A => N100, B => n48, C => n605, D => n359, 
                           Z => n353);
   U584 : HS65_LH_AO212X4 port map( A => n164_port, B => n595, C => n360, D => 
                           alu_i(4), E => n361, Z => n359);
   U585 : HS65_LH_AO222X4 port map( A => n192_port, B => n114_port, C => 
                           n193_port, D => n362, E => n195_port, F => n111_port
                           , Z => n361);
   U586 : HS65_LH_MX41X7 port map( D0 => n70, S0 => n36, D1 => n71, S1 => n32, 
                           D2 => n73, S2 => n27, D3 => n75, S3 => n21, Z => 
                           n362);
   U587 : HS65_LH_AO22X9 port map( A => n602, B => n314, C => alu_i(2), D => 
                           n315, Z => n178_port);
   U588 : HS65_LH_AO22X9 port map( A => n602, B => n324, C => alu_i(2), D => 
                           n216_port, Z => n283);
   U589 : HS65_LH_NAND3X5 port map( A => n353, B => n354, C => n355, Z => 
                           alu_o(1));
   U590 : HS65_LH_AOI212X4 port map( A => n599, B => n303, C => n70, D => n357,
                           E => n358, Z => n354);
   U591 : HS65_LH_AOI212X4 port map( A => n9, B => n71, C => N132, D => n53, E 
                           => n356, Z => n355);
   U592 : HS65_LH_AO212X4 port map( A => n152_port, B => n595, C => n239, D => 
                           alu_i(4), E => n240, Z => n234);
   U593 : HS65_LH_AO222X4 port map( A => n192_port, B => n157_port, C => 
                           n193_port, D => n241, E => n195_port, F => n154_port
                           , Z => n240);
   U594 : HS65_LH_MX41X7 port map( D0 => n71, S0 => n196_port, D1 => n73, S1 =>
                           n31, D2 => n75, S2 => n26, D3 => n77, S3 => n20, Z 
                           => n241);
   U595 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_28_port, B => n45, C => n85
                           , D => n106_port, E => HI_LO_c_HI_28_port, F => n13,
                           Z => n270);
   U596 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_29_port, B => n45, C => n86
                           , D => n106_port, E => HI_LO_c_HI_29_port, F => n13,
                           Z => n246);
   U597 : HS65_LH_AO222X4 port map( A => HI_LO_c_LO_30_port, B => n44, C => n87
                           , D => n106_port, E => HI_LO_c_HI_30_port, F => n13,
                           Z => n221_port);
   U598 : HS65_LH_AO212X4 port map( A => n173_port, B => n595, C => n387, D => 
                           alu_i(4), E => n446, Z => n444);
   U599 : HS65_LH_AO222X4 port map( A => n192_port, B => n130_port, C => 
                           n193_port, D => n447, E => n195_port, F => n128_port
                           , Z => n446);
   U600 : HS65_LH_AO212X4 port map( A => n26, B => n71, C => n34, D => n70, E 
                           => n449, Z => n447);
   U601 : HS65_LH_AO12X9 port map( A => n73, B => n20, C => n315, Z => n449);
   U602 : HS65_LH_AO22X9 port map( A => HI_LO_c_LO_31_port, B => n45, C => n88,
                           D => n106_port, Z => n217_port);
   U603 : HS65_LH_AO212X4 port map( A => n209_port, B => n595, C => n210_port, 
                           D => alu_i(4), E => n211_port, Z => n203_port);
   U604 : HS65_LH_AO222X4 port map( A => n192_port, B => n212_port, C => 
                           n193_port, D => n213_port, E => n195_port, F => 
                           n214_port, Z => n211_port);
   U605 : HS65_LH_AO212X4 port map( A => n26, B => n530, C => n34, D => n531, E
                           => n215_port, Z => n213_port);
   U606 : HS65_LH_AO12X9 port map( A => n528, B => n20, C => n216_port, Z => 
                           n215_port);
   U607 : HS65_LH_NAND4ABX3 port map( A => n169_port, B => n170_port, C => 
                           n171_port, D => n172_port, Z => alu_o(4));
   U608 : HS65_LH_OAI212X5 port map( A => n175_port, B => n76, C => n579, D => 
                           n176_port, E => n177_port, Z => n169_port);
   U609 : HS65_LH_AOI222X2 port map( A => n44, B => HI_LO_c_LO_4_port, C => 
                           n600, D => n173_port, E => N103, F => n47, Z => 
                           n172_port);
   U610 : HS65_LH_NAND4ABX3 port map( A => n160_port, B => n161_port, C => 
                           n162_port, D => n163_port, Z => alu_o(5));
   U611 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n120_port, D1 => n597
                           , S1 => n114_port, D2 => n77, S2 => n167_port, D3 =>
                           n536, S3 => n168_port, Z => n160_port);
   U612 : HS65_LH_AO222X4 port map( A => n165_port, B => n113_port, C => 
                           n111_port, D => n115_port, E => n166_port, F => 
                           n117_port, Z => n161_port);
   U613 : HS65_LH_NAND4ABX3 port map( A => n148_port, B => n149_port, C => 
                           n150_port, D => n151_port, Z => alu_o(6));
   U614 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n156_port, D1 => n597
                           , S1 => n157_port, D2 => n78, S2 => n158_port, D3 =>
                           alu_i(48), S3 => n159_port, Z => n148_port);
   U615 : HS65_LH_AO222X4 port map( A => n153_port, B => n113_port, C => 
                           n154_port, D => n115_port, E => n155_port, F => 
                           n117_port, Z => n149_port);
   U616 : HS65_LH_NAND4ABX3 port map( A => n136_port, B => n137_port, C => 
                           n138_port, D => n139_port, Z => alu_o(7));
   U617 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n144_port, D1 => n597
                           , S1 => n145_port, D2 => n79, S2 => n146_port, D3 =>
                           alu_i(49), S3 => n147_port, Z => n136_port);
   U618 : HS65_LH_AO222X4 port map( A => n141_port, B => n113_port, C => 
                           n142_port, D => n115_port, E => n143_port, F => 
                           n117_port, Z => n137_port);
   U619 : HS65_LH_NAND4ABX3 port map( A => n124_port, B => n125_port, C => 
                           n126_port, D => n127_port, Z => alu_o(8));
   U620 : HS65_LH_MX41X7 port map( D0 => n118_port, S0 => n132_port, D1 => n597
                           , S1 => n133_port, D2 => n80, S2 => n134_port, D3 =>
                           n538, S3 => n135_port, Z => n124_port);
   U621 : HS65_LH_AO222X4 port map( A => n129_port, B => n113_port, C => 
                           n130_port, D => n115_port, E => n131_port, F => 
                           n117_port, Z => n125_port);
   U622 : HS65_LH_NAND2X7 port map( A => n232, B => n233, Z => alu_o(2));
   U623 : HS65_LH_AOI212X4 port map( A => n10, B => n73, C => N133, D => n53, E
                           => n242, Z => n232);
   U624 : HS65_LH_AOI212X4 port map( A => N101, B => n48, C => n605, D => n234,
                           E => n235, Z => n233);
   U625 : HS65_LH_NAND2X7 port map( A => n181_port, B => n182_port, Z => 
                           alu_o(3));
   U626 : HS65_LH_AOI212X4 port map( A => n10, B => n75, C => N134, D => n53, E
                           => n200_port, Z => n181_port);
   U627 : HS65_LH_AOI212X4 port map( A => N102, B => n48, C => n605, D => 
                           n183_port, E => n184_port, Z => n182_port);
   U628 : HS65_LH_OR2X9 port map( A => alu_i(2), B => alu_i(3), Z => n6);
   U629 : HS65_LH_NOR2X6 port map( A => n602, B => alu_i(3), Z => n301);
   U630 : HS65_LH_NOR2X6 port map( A => n602, B => alu_i(3), Z => n7);
   U631 : HS65_LH_IVX9 port map( A => alu_i(4), Z => n596);
   U632 : HS65_LH_AND2X4 port map( A => alu_i(1), B => alu_i(0), Z => n199_port
                           );
   U633 : HS65_LH_NOR2X6 port map( A => n6, B => alu_i(4), Z => n193_port);
   U634 : HS65_LH_NOR2X6 port map( A => n601, B => alu_i(2), Z => n304);
   U635 : HS65_LH_NOR2X6 port map( A => n96, B => alu_i(4), Z => n113_port);
   U636 : HS65_LH_NOR2AX3 port map( A => alu_i(0), B => alu_i(1), Z => 
                           n197_port);
   U637 : HS65_LH_IVX9 port map( A => alu_i(3), Z => n601);
   U638 : HS65_LH_NOR2X6 port map( A => n601, B => alu_i(4), Z => n448);
   U639 : HS65_LH_IVX9 port map( A => alu_i(2), Z => n602);
   U640 : HS65_LH_AND2X4 port map( A => n448, B => alu_i(2), Z => n192_port);
   U641 : HS65_LH_BFX9 port map( A => n196_port, Z => n35);
   U642 : HS65_LH_NOR2X6 port map( A => alu_i(0), B => alu_i(1), Z => n196_port
                           );
   U643 : HS65_LH_BFX9 port map( A => n198_port, Z => n25);
   U644 : HS65_LH_NOR2AX3 port map( A => alu_i(1), B => alu_i(0), Z => 
                           n198_port);
   U645 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_1_port, B => n13, C => 
                           HI_LO_c_LO_1_port, D => n45, Z => n356);
   U646 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_2_port, B => n13, C => 
                           HI_LO_c_LO_2_port, D => n45, Z => n242);
   U647 : HS65_LH_AO22X9 port map( A => HI_LO_c_HI_3_port, B => n13, C => 
                           HI_LO_c_LO_3_port, D => n45, Z => n200_port);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity regfile is

   port( clk, rst_n : in std_logic;  regfile_i : in std_logic_vector (49 downto
         0);  regfile_o : out std_logic_vector (63 downto 0));

end regfile;

architecture SYN_Behavioral of regfile is

   component HS65_LH_AND3X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI22X6
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AOI212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_MX41X7
      port( D0, S0, D1, S1, D2, S2, D3, S3 : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPRQNX9
      port( D, CP, RN : in std_logic;  QN : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal registers_13_31_port, registers_13_30_port, registers_13_29_port, 
      registers_13_28_port, registers_13_27_port, registers_13_26_port, 
      registers_13_25_port, registers_13_24_port, registers_13_23_port, 
      registers_13_22_port, registers_13_21_port, registers_13_20_port, 
      registers_13_19_port, registers_13_18_port, registers_13_17_port, 
      registers_13_16_port, registers_13_15_port, registers_13_14_port, 
      registers_13_13_port, registers_13_12_port, registers_13_11_port, 
      registers_13_10_port, registers_13_9_port, registers_13_8_port, 
      registers_13_7_port, registers_13_6_port, registers_13_5_port, 
      registers_13_4_port, registers_13_3_port, registers_13_2_port, 
      registers_13_1_port, registers_13_0_port, registers_12_31_port, 
      registers_12_30_port, registers_12_29_port, registers_12_28_port, 
      registers_12_27_port, registers_12_26_port, registers_12_25_port, 
      registers_12_24_port, registers_12_23_port, registers_12_22_port, 
      registers_12_21_port, registers_12_20_port, registers_12_19_port, 
      registers_12_18_port, registers_12_17_port, registers_12_16_port, 
      registers_12_15_port, registers_12_14_port, registers_12_13_port, 
      registers_12_12_port, registers_12_11_port, registers_12_10_port, 
      registers_12_9_port, registers_12_8_port, registers_12_7_port, 
      registers_12_6_port, registers_12_5_port, registers_12_4_port, 
      registers_12_3_port, registers_12_2_port, registers_12_1_port, 
      registers_12_0_port, registers_11_31_port, registers_11_30_port, 
      registers_11_29_port, registers_11_28_port, registers_11_27_port, 
      registers_11_26_port, registers_11_25_port, registers_11_24_port, 
      registers_11_23_port, registers_11_22_port, registers_11_21_port, 
      registers_11_20_port, registers_11_19_port, registers_11_18_port, 
      registers_11_17_port, registers_11_16_port, registers_11_15_port, 
      registers_11_14_port, registers_11_13_port, registers_11_12_port, 
      registers_11_11_port, registers_11_10_port, registers_11_9_port, 
      registers_11_8_port, registers_11_7_port, registers_11_6_port, 
      registers_11_5_port, registers_11_4_port, registers_11_3_port, 
      registers_11_2_port, registers_11_1_port, registers_11_0_port, 
      registers_10_31_port, registers_10_30_port, registers_10_29_port, 
      registers_10_28_port, registers_10_27_port, registers_10_26_port, 
      registers_10_25_port, registers_10_24_port, registers_10_23_port, 
      registers_10_22_port, registers_10_21_port, registers_10_20_port, 
      registers_10_19_port, registers_10_18_port, registers_10_17_port, 
      registers_10_16_port, registers_10_15_port, registers_10_14_port, 
      registers_10_13_port, registers_10_12_port, registers_10_11_port, 
      registers_10_10_port, registers_10_9_port, registers_10_8_port, 
      registers_10_7_port, registers_10_6_port, registers_10_5_port, 
      registers_10_4_port, registers_10_3_port, registers_10_2_port, 
      registers_10_1_port, registers_10_0_port, registers_7_31_port, 
      registers_7_30_port, registers_7_29_port, registers_7_28_port, 
      registers_7_27_port, registers_7_26_port, registers_7_25_port, 
      registers_7_24_port, registers_7_23_port, registers_7_22_port, 
      registers_7_21_port, registers_7_20_port, registers_7_19_port, 
      registers_7_18_port, registers_7_17_port, registers_7_16_port, 
      registers_7_15_port, registers_7_14_port, registers_7_13_port, 
      registers_7_12_port, registers_7_11_port, registers_7_10_port, 
      registers_7_9_port, registers_7_8_port, registers_7_7_port, 
      registers_7_6_port, registers_7_5_port, registers_7_4_port, 
      registers_7_3_port, registers_7_2_port, registers_7_1_port, 
      registers_7_0_port, registers_6_31_port, registers_6_30_port, 
      registers_6_29_port, registers_6_28_port, registers_6_27_port, 
      registers_6_26_port, registers_6_25_port, registers_6_24_port, 
      registers_6_23_port, registers_6_22_port, registers_6_21_port, 
      registers_6_20_port, registers_6_19_port, registers_6_18_port, 
      registers_6_17_port, registers_6_16_port, registers_6_15_port, 
      registers_6_14_port, registers_6_13_port, registers_6_12_port, 
      registers_6_11_port, registers_6_10_port, registers_6_9_port, 
      registers_6_8_port, registers_6_7_port, registers_6_6_port, 
      registers_6_5_port, registers_6_4_port, registers_6_3_port, 
      registers_6_2_port, registers_6_1_port, registers_6_0_port, 
      registers_5_31_port, registers_5_30_port, registers_5_29_port, 
      registers_5_28_port, registers_5_27_port, registers_5_26_port, 
      registers_5_25_port, registers_5_24_port, registers_5_23_port, 
      registers_5_22_port, registers_5_21_port, registers_5_20_port, 
      registers_5_19_port, registers_5_18_port, registers_5_17_port, 
      registers_5_16_port, registers_5_15_port, registers_5_14_port, 
      registers_5_13_port, registers_5_12_port, registers_5_11_port, 
      registers_5_10_port, registers_5_9_port, registers_5_8_port, 
      registers_5_7_port, registers_5_6_port, registers_5_5_port, 
      registers_5_4_port, registers_5_3_port, registers_5_2_port, 
      registers_5_1_port, registers_5_0_port, registers_4_31_port, 
      registers_4_30_port, registers_4_29_port, registers_4_28_port, 
      registers_4_27_port, registers_4_26_port, registers_4_25_port, 
      registers_4_24_port, registers_4_23_port, registers_4_22_port, 
      registers_4_21_port, registers_4_20_port, registers_4_19_port, 
      registers_4_18_port, registers_4_17_port, registers_4_16_port, 
      registers_4_15_port, registers_4_14_port, registers_4_13_port, 
      registers_4_12_port, registers_4_11_port, registers_4_10_port, 
      registers_4_9_port, registers_4_8_port, registers_4_7_port, 
      registers_4_6_port, registers_4_5_port, registers_4_4_port, 
      registers_4_3_port, registers_4_2_port, registers_4_1_port, 
      registers_4_0_port, registers_3_31_port, registers_3_30_port, 
      registers_3_29_port, registers_3_28_port, registers_3_27_port, 
      registers_3_26_port, registers_3_25_port, registers_3_24_port, 
      registers_3_23_port, registers_3_22_port, registers_3_21_port, 
      registers_3_20_port, registers_3_19_port, registers_3_18_port, 
      registers_3_17_port, registers_3_16_port, registers_3_15_port, 
      registers_3_14_port, registers_3_13_port, registers_3_12_port, 
      registers_3_11_port, registers_3_10_port, registers_3_9_port, 
      registers_3_8_port, registers_3_7_port, registers_3_6_port, 
      registers_3_5_port, registers_3_4_port, registers_3_3_port, 
      registers_3_2_port, registers_3_1_port, registers_3_0_port, 
      registers_2_31_port, registers_2_30_port, registers_2_29_port, 
      registers_2_28_port, registers_2_27_port, registers_2_26_port, 
      registers_2_25_port, registers_2_24_port, registers_2_23_port, 
      registers_2_22_port, registers_2_21_port, registers_2_20_port, 
      registers_2_19_port, registers_2_18_port, registers_2_17_port, 
      registers_2_16_port, registers_2_15_port, registers_2_14_port, 
      registers_2_13_port, registers_2_12_port, registers_2_11_port, 
      registers_2_10_port, registers_2_9_port, registers_2_8_port, 
      registers_2_7_port, registers_2_6_port, registers_2_5_port, 
      registers_2_4_port, registers_2_3_port, registers_2_2_port, 
      registers_2_1_port, registers_2_0_port, registers_1_31_port, 
      registers_1_30_port, registers_1_29_port, registers_1_28_port, 
      registers_1_27_port, registers_1_26_port, registers_1_25_port, 
      registers_1_24_port, registers_1_23_port, registers_1_22_port, 
      registers_1_21_port, registers_1_20_port, registers_1_19_port, 
      registers_1_18_port, registers_1_17_port, registers_1_16_port, 
      registers_1_15_port, registers_1_14_port, registers_1_13_port, 
      registers_1_12_port, registers_1_11_port, registers_1_10_port, 
      registers_1_9_port, registers_1_8_port, registers_1_7_port, 
      registers_1_6_port, registers_1_5_port, registers_1_4_port, 
      registers_1_3_port, registers_1_2_port, registers_1_1_port, 
      registers_1_0_port, registers_31_31_port, registers_31_30_port, 
      registers_31_29_port, registers_31_28_port, registers_31_27_port, 
      registers_31_26_port, registers_31_25_port, registers_31_24_port, 
      registers_31_23_port, registers_31_22_port, registers_31_21_port, 
      registers_31_20_port, registers_31_19_port, registers_31_18_port, 
      registers_31_17_port, registers_31_16_port, registers_31_15_port, 
      registers_31_14_port, registers_31_13_port, registers_31_12_port, 
      registers_31_11_port, registers_31_10_port, registers_31_9_port, 
      registers_31_8_port, registers_31_7_port, registers_31_6_port, 
      registers_31_5_port, registers_31_4_port, registers_31_3_port, 
      registers_31_2_port, registers_31_1_port, registers_31_0_port, 
      registers_30_31_port, registers_30_30_port, registers_30_29_port, 
      registers_30_28_port, registers_30_27_port, registers_30_26_port, 
      registers_30_25_port, registers_30_24_port, registers_30_23_port, 
      registers_30_22_port, registers_30_21_port, registers_30_20_port, 
      registers_30_19_port, registers_30_18_port, registers_30_17_port, 
      registers_30_16_port, registers_30_15_port, registers_30_14_port, 
      registers_30_13_port, registers_30_12_port, registers_30_11_port, 
      registers_30_10_port, registers_30_9_port, registers_30_8_port, 
      registers_30_7_port, registers_30_6_port, registers_30_5_port, 
      registers_30_4_port, registers_30_3_port, registers_30_2_port, 
      registers_30_1_port, registers_30_0_port, registers_25_31_port, 
      registers_25_30_port, registers_25_29_port, registers_25_28_port, 
      registers_25_27_port, registers_25_26_port, registers_25_25_port, 
      registers_25_24_port, registers_25_23_port, registers_25_22_port, 
      registers_25_21_port, registers_25_20_port, registers_25_19_port, 
      registers_25_18_port, registers_25_17_port, registers_25_16_port, 
      registers_25_15_port, registers_25_14_port, registers_25_13_port, 
      registers_25_12_port, registers_25_11_port, registers_25_10_port, 
      registers_25_9_port, registers_25_8_port, registers_25_7_port, 
      registers_25_6_port, registers_25_5_port, registers_25_4_port, 
      registers_25_3_port, registers_25_2_port, registers_25_1_port, 
      registers_25_0_port, registers_24_31_port, registers_24_30_port, 
      registers_24_29_port, registers_24_28_port, registers_24_27_port, 
      registers_24_26_port, registers_24_25_port, registers_24_24_port, 
      registers_24_23_port, registers_24_22_port, registers_24_21_port, 
      registers_24_20_port, registers_24_19_port, registers_24_18_port, 
      registers_24_17_port, registers_24_16_port, registers_24_15_port, 
      registers_24_14_port, registers_24_13_port, registers_24_12_port, 
      registers_24_11_port, registers_24_10_port, registers_24_9_port, 
      registers_24_8_port, registers_24_7_port, registers_24_6_port, 
      registers_24_5_port, registers_24_4_port, registers_24_3_port, 
      registers_24_2_port, registers_24_1_port, registers_24_0_port, 
      registers_23_31_port, registers_23_30_port, registers_23_29_port, 
      registers_23_28_port, registers_23_27_port, registers_23_26_port, 
      registers_23_25_port, registers_23_24_port, registers_23_23_port, 
      registers_23_22_port, registers_23_21_port, registers_23_20_port, 
      registers_23_19_port, registers_23_18_port, registers_23_17_port, 
      registers_23_16_port, registers_23_15_port, registers_23_14_port, 
      registers_23_13_port, registers_23_12_port, registers_23_11_port, 
      registers_23_10_port, registers_23_9_port, registers_23_8_port, 
      registers_23_7_port, registers_23_6_port, registers_23_5_port, 
      registers_23_4_port, registers_23_3_port, registers_23_2_port, 
      registers_23_1_port, registers_23_0_port, registers_22_31_port, 
      registers_22_30_port, registers_22_29_port, registers_22_28_port, 
      registers_22_27_port, registers_22_26_port, registers_22_25_port, 
      registers_22_24_port, registers_22_23_port, registers_22_22_port, 
      registers_22_21_port, registers_22_20_port, registers_22_19_port, 
      registers_22_18_port, registers_22_17_port, registers_22_16_port, 
      registers_22_15_port, registers_22_14_port, registers_22_13_port, 
      registers_22_12_port, registers_22_11_port, registers_22_10_port, 
      registers_22_9_port, registers_22_8_port, registers_22_7_port, 
      registers_22_6_port, registers_22_5_port, registers_22_4_port, 
      registers_22_3_port, registers_22_2_port, registers_22_1_port, 
      registers_22_0_port, registers_21_31_port, registers_21_30_port, 
      registers_21_29_port, registers_21_28_port, registers_21_27_port, 
      registers_21_26_port, registers_21_25_port, registers_21_24_port, 
      registers_21_23_port, registers_21_22_port, registers_21_21_port, 
      registers_21_20_port, registers_21_19_port, registers_21_18_port, 
      registers_21_17_port, registers_21_16_port, registers_21_15_port, 
      registers_21_14_port, registers_21_13_port, registers_21_12_port, 
      registers_21_11_port, registers_21_10_port, registers_21_9_port, 
      registers_21_8_port, registers_21_7_port, registers_21_6_port, 
      registers_21_5_port, registers_21_4_port, registers_21_3_port, 
      registers_21_2_port, registers_21_1_port, registers_21_0_port, 
      registers_20_31_port, registers_20_30_port, registers_20_29_port, 
      registers_20_28_port, registers_20_27_port, registers_20_26_port, 
      registers_20_25_port, registers_20_24_port, registers_20_23_port, 
      registers_20_22_port, registers_20_21_port, registers_20_20_port, 
      registers_20_19_port, registers_20_18_port, registers_20_17_port, 
      registers_20_16_port, registers_20_15_port, registers_20_14_port, 
      registers_20_13_port, registers_20_12_port, registers_20_11_port, 
      registers_20_10_port, registers_20_9_port, registers_20_8_port, 
      registers_20_7_port, registers_20_6_port, registers_20_5_port, 
      registers_20_4_port, registers_20_3_port, registers_20_2_port, 
      registers_20_1_port, registers_20_0_port, registers_19_31_port, 
      registers_19_30_port, registers_19_29_port, registers_19_28_port, 
      registers_19_27_port, registers_19_26_port, registers_19_25_port, 
      registers_19_24_port, registers_19_23_port, registers_19_22_port, 
      registers_19_21_port, registers_19_20_port, registers_19_19_port, 
      registers_19_18_port, registers_19_17_port, registers_19_16_port, 
      registers_19_15_port, registers_19_14_port, registers_19_13_port, 
      registers_19_12_port, registers_19_11_port, registers_19_10_port, 
      registers_19_9_port, registers_19_8_port, registers_19_7_port, 
      registers_19_6_port, registers_19_5_port, registers_19_4_port, 
      registers_19_3_port, registers_19_2_port, registers_19_1_port, 
      registers_19_0_port, registers_18_31_port, registers_18_30_port, 
      registers_18_29_port, registers_18_28_port, registers_18_27_port, 
      registers_18_26_port, registers_18_25_port, registers_18_24_port, 
      registers_18_23_port, registers_18_22_port, registers_18_21_port, 
      registers_18_20_port, registers_18_19_port, registers_18_18_port, 
      registers_18_17_port, registers_18_16_port, registers_18_15_port, 
      registers_18_14_port, registers_18_13_port, registers_18_12_port, 
      registers_18_11_port, registers_18_10_port, registers_18_9_port, 
      registers_18_8_port, registers_18_7_port, registers_18_6_port, 
      registers_18_5_port, registers_18_4_port, registers_18_3_port, 
      registers_18_2_port, registers_18_1_port, registers_18_0_port, 
      registers_17_31_port, registers_17_30_port, registers_17_29_port, 
      registers_17_28_port, registers_17_27_port, registers_17_26_port, 
      registers_17_25_port, registers_17_24_port, registers_17_23_port, 
      registers_17_22_port, registers_17_21_port, registers_17_20_port, 
      registers_17_19_port, registers_17_18_port, registers_17_17_port, 
      registers_17_16_port, registers_17_15_port, registers_17_14_port, 
      registers_17_13_port, registers_17_12_port, registers_17_11_port, 
      registers_17_10_port, registers_17_9_port, registers_17_8_port, 
      registers_17_7_port, registers_17_6_port, registers_17_5_port, 
      registers_17_4_port, registers_17_3_port, registers_17_2_port, 
      registers_17_1_port, registers_17_0_port, registers_16_31_port, 
      registers_16_30_port, registers_16_29_port, registers_16_28_port, 
      registers_16_27_port, registers_16_26_port, registers_16_25_port, 
      registers_16_24_port, registers_16_23_port, registers_16_22_port, 
      registers_16_21_port, registers_16_20_port, registers_16_19_port, 
      registers_16_18_port, registers_16_17_port, registers_16_16_port, 
      registers_16_15_port, registers_16_14_port, registers_16_13_port, 
      registers_16_12_port, registers_16_11_port, registers_16_10_port, 
      registers_16_9_port, registers_16_8_port, registers_16_7_port, 
      registers_16_6_port, registers_16_5_port, registers_16_4_port, 
      registers_16_3_port, registers_16_2_port, registers_16_1_port, 
      registers_16_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
      n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
      n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n877, n878, n879, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1393, n1394, n1396, n1398, n1400, 
      n1402, n1404, n1406, n1407, n1408, n1409, n1414, n1415, n1416, n1417, 
      n1425, n1426, n1428, n1429, n1430, n1431, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
      n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
      n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, 
      n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
      n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
      n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
      n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, 
      n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, 
      n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, 
      n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, 
      n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, 
      n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, 
      n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
      n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
      n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, 
      n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
      n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, 
      n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, 
      n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, 
      n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, 
      n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, 
      n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, 
      n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
      n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, 
      n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, 
      n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n257, n258, n259,
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n352, n880, n1392, n1395, n1397, n1399, n1401, n1403, 
      n1405, n1410, n1411, n1412, n1413, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1427, n1432, n1433, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
      n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
      n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
      n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
      n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
      n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
      n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, 
      n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, 
      n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
      n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
      n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
      n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
      n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
      n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
      n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
      n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
      n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
      n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
      n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
      n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
      n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
      n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
      n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
      n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
      n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
      n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
      n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, 
      n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
      n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
      n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
      n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
      n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
      n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
      n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, 
      n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, 
      n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
      n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
      n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, 
      n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
      n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099 : std_logic
      ;

begin
   
   registers_reg_31_31_inst : HS65_LH_DFPRQX9 port map( D => n2425, CP => clk, 
                           RN => n2765, Q => registers_31_31_port);
   registers_reg_31_30_inst : HS65_LH_DFPRQX9 port map( D => n2424, CP => clk, 
                           RN => n2817, Q => registers_31_30_port);
   registers_reg_31_29_inst : HS65_LH_DFPRQX9 port map( D => n2423, CP => clk, 
                           RN => n2816, Q => registers_31_29_port);
   registers_reg_31_28_inst : HS65_LH_DFPRQX9 port map( D => n2422, CP => clk, 
                           RN => n2816, Q => registers_31_28_port);
   registers_reg_31_27_inst : HS65_LH_DFPRQX9 port map( D => n2421, CP => clk, 
                           RN => n2816, Q => registers_31_27_port);
   registers_reg_31_26_inst : HS65_LH_DFPRQX9 port map( D => n2420, CP => clk, 
                           RN => n2816, Q => registers_31_26_port);
   registers_reg_31_25_inst : HS65_LH_DFPRQX9 port map( D => n2419, CP => clk, 
                           RN => n2815, Q => registers_31_25_port);
   registers_reg_31_24_inst : HS65_LH_DFPRQX9 port map( D => n2418, CP => clk, 
                           RN => n2815, Q => registers_31_24_port);
   registers_reg_31_23_inst : HS65_LH_DFPRQX9 port map( D => n2417, CP => clk, 
                           RN => n2815, Q => registers_31_23_port);
   registers_reg_31_22_inst : HS65_LH_DFPRQX9 port map( D => n2416, CP => clk, 
                           RN => n2815, Q => registers_31_22_port);
   registers_reg_31_21_inst : HS65_LH_DFPRQX9 port map( D => n2415, CP => clk, 
                           RN => n2815, Q => registers_31_21_port);
   registers_reg_31_20_inst : HS65_LH_DFPRQX9 port map( D => n2414, CP => clk, 
                           RN => n2815, Q => registers_31_20_port);
   registers_reg_31_19_inst : HS65_LH_DFPRQX9 port map( D => n2413, CP => clk, 
                           RN => n2815, Q => registers_31_19_port);
   registers_reg_31_18_inst : HS65_LH_DFPRQX9 port map( D => n2412, CP => clk, 
                           RN => n2815, Q => registers_31_18_port);
   registers_reg_31_17_inst : HS65_LH_DFPRQX9 port map( D => n2411, CP => clk, 
                           RN => n2815, Q => registers_31_17_port);
   registers_reg_31_16_inst : HS65_LH_DFPRQX9 port map( D => n2410, CP => clk, 
                           RN => n2815, Q => registers_31_16_port);
   registers_reg_31_15_inst : HS65_LH_DFPRQX9 port map( D => n2409, CP => clk, 
                           RN => n2815, Q => registers_31_15_port);
   registers_reg_31_14_inst : HS65_LH_DFPRQX9 port map( D => n2408, CP => clk, 
                           RN => n2815, Q => registers_31_14_port);
   registers_reg_31_13_inst : HS65_LH_DFPRQX9 port map( D => n2407, CP => clk, 
                           RN => n2814, Q => registers_31_13_port);
   registers_reg_31_12_inst : HS65_LH_DFPRQX9 port map( D => n2406, CP => clk, 
                           RN => n2814, Q => registers_31_12_port);
   registers_reg_31_11_inst : HS65_LH_DFPRQX9 port map( D => n2405, CP => clk, 
                           RN => n2814, Q => registers_31_11_port);
   registers_reg_31_10_inst : HS65_LH_DFPRQX9 port map( D => n2404, CP => clk, 
                           RN => n2814, Q => registers_31_10_port);
   registers_reg_31_9_inst : HS65_LH_DFPRQX9 port map( D => n2403, CP => clk, 
                           RN => n2814, Q => registers_31_9_port);
   registers_reg_31_8_inst : HS65_LH_DFPRQX9 port map( D => n2402, CP => clk, 
                           RN => n2814, Q => registers_31_8_port);
   registers_reg_31_7_inst : HS65_LH_DFPRQX9 port map( D => n2401, CP => clk, 
                           RN => n2814, Q => registers_31_7_port);
   registers_reg_31_6_inst : HS65_LH_DFPRQX9 port map( D => n2400, CP => clk, 
                           RN => n2814, Q => registers_31_6_port);
   registers_reg_31_5_inst : HS65_LH_DFPRQX9 port map( D => n2399, CP => clk, 
                           RN => n2814, Q => registers_31_5_port);
   registers_reg_31_4_inst : HS65_LH_DFPRQX9 port map( D => n2398, CP => clk, 
                           RN => n2814, Q => registers_31_4_port);
   registers_reg_31_3_inst : HS65_LH_DFPRQX9 port map( D => n2397, CP => clk, 
                           RN => n2814, Q => registers_31_3_port);
   registers_reg_31_2_inst : HS65_LH_DFPRQX9 port map( D => n2396, CP => clk, 
                           RN => n2814, Q => registers_31_2_port);
   registers_reg_31_1_inst : HS65_LH_DFPRQX9 port map( D => n2395, CP => clk, 
                           RN => n2813, Q => registers_31_1_port);
   registers_reg_31_0_inst : HS65_LH_DFPRQX9 port map( D => n2394, CP => clk, 
                           RN => n2813, Q => registers_31_0_port);
   registers_reg_30_31_inst : HS65_LH_DFPRQX9 port map( D => n2393, CP => clk, 
                           RN => n2813, Q => registers_30_31_port);
   registers_reg_30_30_inst : HS65_LH_DFPRQX9 port map( D => n2392, CP => clk, 
                           RN => n2813, Q => registers_30_30_port);
   registers_reg_30_29_inst : HS65_LH_DFPRQX9 port map( D => n2391, CP => clk, 
                           RN => n2813, Q => registers_30_29_port);
   registers_reg_30_28_inst : HS65_LH_DFPRQX9 port map( D => n2390, CP => clk, 
                           RN => n2813, Q => registers_30_28_port);
   registers_reg_30_27_inst : HS65_LH_DFPRQX9 port map( D => n2389, CP => clk, 
                           RN => n2813, Q => registers_30_27_port);
   registers_reg_30_26_inst : HS65_LH_DFPRQX9 port map( D => n2388, CP => clk, 
                           RN => n2813, Q => registers_30_26_port);
   registers_reg_30_25_inst : HS65_LH_DFPRQX9 port map( D => n2387, CP => clk, 
                           RN => n2813, Q => registers_30_25_port);
   registers_reg_30_24_inst : HS65_LH_DFPRQX9 port map( D => n2386, CP => clk, 
                           RN => n2813, Q => registers_30_24_port);
   registers_reg_30_23_inst : HS65_LH_DFPRQX9 port map( D => n2385, CP => clk, 
                           RN => n2813, Q => registers_30_23_port);
   registers_reg_30_22_inst : HS65_LH_DFPRQX9 port map( D => n2384, CP => clk, 
                           RN => n2813, Q => registers_30_22_port);
   registers_reg_30_21_inst : HS65_LH_DFPRQX9 port map( D => n2383, CP => clk, 
                           RN => n2812, Q => registers_30_21_port);
   registers_reg_30_20_inst : HS65_LH_DFPRQX9 port map( D => n2382, CP => clk, 
                           RN => n2812, Q => registers_30_20_port);
   registers_reg_30_19_inst : HS65_LH_DFPRQX9 port map( D => n2381, CP => clk, 
                           RN => n2812, Q => registers_30_19_port);
   registers_reg_30_18_inst : HS65_LH_DFPRQX9 port map( D => n2380, CP => clk, 
                           RN => n2812, Q => registers_30_18_port);
   registers_reg_30_17_inst : HS65_LH_DFPRQX9 port map( D => n2379, CP => clk, 
                           RN => n2812, Q => registers_30_17_port);
   registers_reg_30_16_inst : HS65_LH_DFPRQX9 port map( D => n2378, CP => clk, 
                           RN => n2812, Q => registers_30_16_port);
   registers_reg_30_15_inst : HS65_LH_DFPRQX9 port map( D => n2377, CP => clk, 
                           RN => n2812, Q => registers_30_15_port);
   registers_reg_30_14_inst : HS65_LH_DFPRQX9 port map( D => n2376, CP => clk, 
                           RN => n2812, Q => registers_30_14_port);
   registers_reg_30_13_inst : HS65_LH_DFPRQX9 port map( D => n2375, CP => clk, 
                           RN => n2812, Q => registers_30_13_port);
   registers_reg_30_12_inst : HS65_LH_DFPRQX9 port map( D => n2374, CP => clk, 
                           RN => n2812, Q => registers_30_12_port);
   registers_reg_30_11_inst : HS65_LH_DFPRQX9 port map( D => n2373, CP => clk, 
                           RN => n2812, Q => registers_30_11_port);
   registers_reg_30_10_inst : HS65_LH_DFPRQX9 port map( D => n2372, CP => clk, 
                           RN => n2812, Q => registers_30_10_port);
   registers_reg_30_9_inst : HS65_LH_DFPRQX9 port map( D => n2371, CP => clk, 
                           RN => n2811, Q => registers_30_9_port);
   registers_reg_30_8_inst : HS65_LH_DFPRQX9 port map( D => n2370, CP => clk, 
                           RN => n2811, Q => registers_30_8_port);
   registers_reg_30_7_inst : HS65_LH_DFPRQX9 port map( D => n2369, CP => clk, 
                           RN => n2811, Q => registers_30_7_port);
   registers_reg_30_6_inst : HS65_LH_DFPRQX9 port map( D => n2368, CP => clk, 
                           RN => n2811, Q => registers_30_6_port);
   registers_reg_30_5_inst : HS65_LH_DFPRQX9 port map( D => n2367, CP => clk, 
                           RN => n2811, Q => registers_30_5_port);
   registers_reg_30_4_inst : HS65_LH_DFPRQX9 port map( D => n2366, CP => clk, 
                           RN => n2811, Q => registers_30_4_port);
   registers_reg_30_3_inst : HS65_LH_DFPRQX9 port map( D => n2365, CP => clk, 
                           RN => n2811, Q => registers_30_3_port);
   registers_reg_30_2_inst : HS65_LH_DFPRQX9 port map( D => n2364, CP => clk, 
                           RN => n2811, Q => registers_30_2_port);
   registers_reg_30_1_inst : HS65_LH_DFPRQX9 port map( D => n2363, CP => clk, 
                           RN => n2811, Q => registers_30_1_port);
   registers_reg_30_0_inst : HS65_LH_DFPRQX9 port map( D => n2362, CP => clk, 
                           RN => n2811, Q => registers_30_0_port);
   registers_reg_25_31_inst : HS65_LH_DFPRQX9 port map( D => n2233, CP => clk, 
                           RN => n2811, Q => registers_25_31_port);
   registers_reg_25_30_inst : HS65_LH_DFPRQX9 port map( D => n2232, CP => clk, 
                           RN => n2811, Q => registers_25_30_port);
   registers_reg_25_29_inst : HS65_LH_DFPRQX9 port map( D => n2231, CP => clk, 
                           RN => n2810, Q => registers_25_29_port);
   registers_reg_25_28_inst : HS65_LH_DFPRQX9 port map( D => n2230, CP => clk, 
                           RN => n2810, Q => registers_25_28_port);
   registers_reg_25_27_inst : HS65_LH_DFPRQX9 port map( D => n2229, CP => clk, 
                           RN => n2810, Q => registers_25_27_port);
   registers_reg_25_26_inst : HS65_LH_DFPRQX9 port map( D => n2228, CP => clk, 
                           RN => n2810, Q => registers_25_26_port);
   registers_reg_25_25_inst : HS65_LH_DFPRQX9 port map( D => n2227, CP => clk, 
                           RN => n2810, Q => registers_25_25_port);
   registers_reg_25_24_inst : HS65_LH_DFPRQX9 port map( D => n2226, CP => clk, 
                           RN => n2810, Q => registers_25_24_port);
   registers_reg_25_23_inst : HS65_LH_DFPRQX9 port map( D => n2225, CP => clk, 
                           RN => n2810, Q => registers_25_23_port);
   registers_reg_25_22_inst : HS65_LH_DFPRQX9 port map( D => n2224, CP => clk, 
                           RN => n2810, Q => registers_25_22_port);
   registers_reg_25_21_inst : HS65_LH_DFPRQX9 port map( D => n2223, CP => clk, 
                           RN => n2810, Q => registers_25_21_port);
   registers_reg_25_20_inst : HS65_LH_DFPRQX9 port map( D => n2222, CP => clk, 
                           RN => n2810, Q => registers_25_20_port);
   registers_reg_25_19_inst : HS65_LH_DFPRQX9 port map( D => n2221, CP => clk, 
                           RN => n2810, Q => registers_25_19_port);
   registers_reg_25_18_inst : HS65_LH_DFPRQX9 port map( D => n2220, CP => clk, 
                           RN => n2810, Q => registers_25_18_port);
   registers_reg_25_17_inst : HS65_LH_DFPRQX9 port map( D => n2219, CP => clk, 
                           RN => n2809, Q => registers_25_17_port);
   registers_reg_25_16_inst : HS65_LH_DFPRQX9 port map( D => n2218, CP => clk, 
                           RN => n2809, Q => registers_25_16_port);
   registers_reg_25_15_inst : HS65_LH_DFPRQX9 port map( D => n2217, CP => clk, 
                           RN => n2809, Q => registers_25_15_port);
   registers_reg_25_14_inst : HS65_LH_DFPRQX9 port map( D => n2216, CP => clk, 
                           RN => n2809, Q => registers_25_14_port);
   registers_reg_25_13_inst : HS65_LH_DFPRQX9 port map( D => n2215, CP => clk, 
                           RN => n2809, Q => registers_25_13_port);
   registers_reg_25_12_inst : HS65_LH_DFPRQX9 port map( D => n2214, CP => clk, 
                           RN => n2809, Q => registers_25_12_port);
   registers_reg_25_11_inst : HS65_LH_DFPRQX9 port map( D => n2213, CP => clk, 
                           RN => n2809, Q => registers_25_11_port);
   registers_reg_25_10_inst : HS65_LH_DFPRQX9 port map( D => n2212, CP => clk, 
                           RN => n2809, Q => registers_25_10_port);
   registers_reg_25_9_inst : HS65_LH_DFPRQX9 port map( D => n2211, CP => clk, 
                           RN => n2809, Q => registers_25_9_port);
   registers_reg_25_8_inst : HS65_LH_DFPRQX9 port map( D => n2210, CP => clk, 
                           RN => n2809, Q => registers_25_8_port);
   registers_reg_25_7_inst : HS65_LH_DFPRQX9 port map( D => n2209, CP => clk, 
                           RN => n2809, Q => registers_25_7_port);
   registers_reg_25_6_inst : HS65_LH_DFPRQX9 port map( D => n2208, CP => clk, 
                           RN => n2809, Q => registers_25_6_port);
   registers_reg_25_5_inst : HS65_LH_DFPRQX9 port map( D => n2207, CP => clk, 
                           RN => n2808, Q => registers_25_5_port);
   registers_reg_25_4_inst : HS65_LH_DFPRQX9 port map( D => n2206, CP => clk, 
                           RN => n2808, Q => registers_25_4_port);
   registers_reg_25_3_inst : HS65_LH_DFPRQX9 port map( D => n2205, CP => clk, 
                           RN => n2808, Q => registers_25_3_port);
   registers_reg_25_2_inst : HS65_LH_DFPRQX9 port map( D => n2204, CP => clk, 
                           RN => n2808, Q => registers_25_2_port);
   registers_reg_25_1_inst : HS65_LH_DFPRQX9 port map( D => n2203, CP => clk, 
                           RN => n2808, Q => registers_25_1_port);
   registers_reg_25_0_inst : HS65_LH_DFPRQX9 port map( D => n2202, CP => clk, 
                           RN => n2808, Q => registers_25_0_port);
   registers_reg_24_31_inst : HS65_LH_DFPRQX9 port map( D => n2201, CP => clk, 
                           RN => n2808, Q => registers_24_31_port);
   registers_reg_24_30_inst : HS65_LH_DFPRQX9 port map( D => n2200, CP => clk, 
                           RN => n2808, Q => registers_24_30_port);
   registers_reg_24_29_inst : HS65_LH_DFPRQX9 port map( D => n2199, CP => clk, 
                           RN => n2808, Q => registers_24_29_port);
   registers_reg_24_28_inst : HS65_LH_DFPRQX9 port map( D => n2198, CP => clk, 
                           RN => n2808, Q => registers_24_28_port);
   registers_reg_24_27_inst : HS65_LH_DFPRQX9 port map( D => n2197, CP => clk, 
                           RN => n2808, Q => registers_24_27_port);
   registers_reg_24_26_inst : HS65_LH_DFPRQX9 port map( D => n2196, CP => clk, 
                           RN => n2807, Q => registers_24_26_port);
   registers_reg_24_25_inst : HS65_LH_DFPRQX9 port map( D => n2195, CP => clk, 
                           RN => n2807, Q => registers_24_25_port);
   registers_reg_24_24_inst : HS65_LH_DFPRQX9 port map( D => n2194, CP => clk, 
                           RN => n2807, Q => registers_24_24_port);
   registers_reg_24_23_inst : HS65_LH_DFPRQX9 port map( D => n2193, CP => clk, 
                           RN => n2807, Q => registers_24_23_port);
   registers_reg_24_22_inst : HS65_LH_DFPRQX9 port map( D => n2192, CP => clk, 
                           RN => n2807, Q => registers_24_22_port);
   registers_reg_24_21_inst : HS65_LH_DFPRQX9 port map( D => n2191, CP => clk, 
                           RN => n2807, Q => registers_24_21_port);
   registers_reg_24_20_inst : HS65_LH_DFPRQX9 port map( D => n2190, CP => clk, 
                           RN => n2807, Q => registers_24_20_port);
   registers_reg_24_19_inst : HS65_LH_DFPRQX9 port map( D => n2189, CP => clk, 
                           RN => n2807, Q => registers_24_19_port);
   registers_reg_24_18_inst : HS65_LH_DFPRQX9 port map( D => n2188, CP => clk, 
                           RN => n2807, Q => registers_24_18_port);
   registers_reg_24_17_inst : HS65_LH_DFPRQX9 port map( D => n2187, CP => clk, 
                           RN => n2807, Q => registers_24_17_port);
   registers_reg_24_16_inst : HS65_LH_DFPRQX9 port map( D => n2186, CP => clk, 
                           RN => n2807, Q => registers_24_16_port);
   registers_reg_24_15_inst : HS65_LH_DFPRQX9 port map( D => n2185, CP => clk, 
                           RN => n2807, Q => registers_24_15_port);
   registers_reg_24_14_inst : HS65_LH_DFPRQX9 port map( D => n2184, CP => clk, 
                           RN => n2806, Q => registers_24_14_port);
   registers_reg_24_13_inst : HS65_LH_DFPRQX9 port map( D => n2183, CP => clk, 
                           RN => n2806, Q => registers_24_13_port);
   registers_reg_24_12_inst : HS65_LH_DFPRQX9 port map( D => n2182, CP => clk, 
                           RN => n2806, Q => registers_24_12_port);
   registers_reg_24_11_inst : HS65_LH_DFPRQX9 port map( D => n2181, CP => clk, 
                           RN => n2806, Q => registers_24_11_port);
   registers_reg_24_10_inst : HS65_LH_DFPRQX9 port map( D => n2180, CP => clk, 
                           RN => n2806, Q => registers_24_10_port);
   registers_reg_24_9_inst : HS65_LH_DFPRQX9 port map( D => n2179, CP => clk, 
                           RN => n2806, Q => registers_24_9_port);
   registers_reg_24_8_inst : HS65_LH_DFPRQX9 port map( D => n2178, CP => clk, 
                           RN => n2806, Q => registers_24_8_port);
   registers_reg_24_7_inst : HS65_LH_DFPRQX9 port map( D => n2177, CP => clk, 
                           RN => n2806, Q => registers_24_7_port);
   registers_reg_24_6_inst : HS65_LH_DFPRQX9 port map( D => n2176, CP => clk, 
                           RN => n2806, Q => registers_24_6_port);
   registers_reg_24_5_inst : HS65_LH_DFPRQX9 port map( D => n2175, CP => clk, 
                           RN => n2806, Q => registers_24_5_port);
   registers_reg_24_4_inst : HS65_LH_DFPRQX9 port map( D => n2174, CP => clk, 
                           RN => n2806, Q => registers_24_4_port);
   registers_reg_24_3_inst : HS65_LH_DFPRQX9 port map( D => n2173, CP => clk, 
                           RN => n2806, Q => registers_24_3_port);
   registers_reg_24_2_inst : HS65_LH_DFPRQX9 port map( D => n2172, CP => clk, 
                           RN => n2805, Q => registers_24_2_port);
   registers_reg_24_1_inst : HS65_LH_DFPRQX9 port map( D => n2171, CP => clk, 
                           RN => n2805, Q => registers_24_1_port);
   registers_reg_24_0_inst : HS65_LH_DFPRQX9 port map( D => n2170, CP => clk, 
                           RN => n2805, Q => registers_24_0_port);
   registers_reg_23_31_inst : HS65_LH_DFPRQX9 port map( D => n2169, CP => clk, 
                           RN => n2805, Q => registers_23_31_port);
   registers_reg_23_30_inst : HS65_LH_DFPRQX9 port map( D => n2168, CP => clk, 
                           RN => n2805, Q => registers_23_30_port);
   registers_reg_23_29_inst : HS65_LH_DFPRQX9 port map( D => n2167, CP => clk, 
                           RN => n2805, Q => registers_23_29_port);
   registers_reg_23_28_inst : HS65_LH_DFPRQX9 port map( D => n2166, CP => clk, 
                           RN => n2805, Q => registers_23_28_port);
   registers_reg_23_27_inst : HS65_LH_DFPRQX9 port map( D => n2165, CP => clk, 
                           RN => n2805, Q => registers_23_27_port);
   registers_reg_23_26_inst : HS65_LH_DFPRQX9 port map( D => n2164, CP => clk, 
                           RN => n2805, Q => registers_23_26_port);
   registers_reg_23_25_inst : HS65_LH_DFPRQX9 port map( D => n2163, CP => clk, 
                           RN => n2805, Q => registers_23_25_port);
   registers_reg_23_24_inst : HS65_LH_DFPRQX9 port map( D => n2162, CP => clk, 
                           RN => n2805, Q => registers_23_24_port);
   registers_reg_23_23_inst : HS65_LH_DFPRQX9 port map( D => n2161, CP => clk, 
                           RN => n2805, Q => registers_23_23_port);
   registers_reg_23_22_inst : HS65_LH_DFPRQX9 port map( D => n2160, CP => clk, 
                           RN => n2804, Q => registers_23_22_port);
   registers_reg_23_21_inst : HS65_LH_DFPRQX9 port map( D => n2159, CP => clk, 
                           RN => n2804, Q => registers_23_21_port);
   registers_reg_23_20_inst : HS65_LH_DFPRQX9 port map( D => n2158, CP => clk, 
                           RN => n2804, Q => registers_23_20_port);
   registers_reg_23_19_inst : HS65_LH_DFPRQX9 port map( D => n2157, CP => clk, 
                           RN => n2804, Q => registers_23_19_port);
   registers_reg_23_18_inst : HS65_LH_DFPRQX9 port map( D => n2156, CP => clk, 
                           RN => n2804, Q => registers_23_18_port);
   registers_reg_23_17_inst : HS65_LH_DFPRQX9 port map( D => n2155, CP => clk, 
                           RN => n2804, Q => registers_23_17_port);
   registers_reg_23_16_inst : HS65_LH_DFPRQX9 port map( D => n2154, CP => clk, 
                           RN => n2804, Q => registers_23_16_port);
   registers_reg_23_15_inst : HS65_LH_DFPRQX9 port map( D => n2153, CP => clk, 
                           RN => n2804, Q => registers_23_15_port);
   registers_reg_23_14_inst : HS65_LH_DFPRQX9 port map( D => n2152, CP => clk, 
                           RN => n2804, Q => registers_23_14_port);
   registers_reg_23_13_inst : HS65_LH_DFPRQX9 port map( D => n2151, CP => clk, 
                           RN => n2804, Q => registers_23_13_port);
   registers_reg_23_12_inst : HS65_LH_DFPRQX9 port map( D => n2150, CP => clk, 
                           RN => n2804, Q => registers_23_12_port);
   registers_reg_23_11_inst : HS65_LH_DFPRQX9 port map( D => n2149, CP => clk, 
                           RN => n2804, Q => registers_23_11_port);
   registers_reg_23_10_inst : HS65_LH_DFPRQX9 port map( D => n2148, CP => clk, 
                           RN => n2803, Q => registers_23_10_port);
   registers_reg_23_9_inst : HS65_LH_DFPRQX9 port map( D => n2147, CP => clk, 
                           RN => n2803, Q => registers_23_9_port);
   registers_reg_23_8_inst : HS65_LH_DFPRQX9 port map( D => n2146, CP => clk, 
                           RN => n2803, Q => registers_23_8_port);
   registers_reg_23_7_inst : HS65_LH_DFPRQX9 port map( D => n2145, CP => clk, 
                           RN => n2803, Q => registers_23_7_port);
   registers_reg_23_6_inst : HS65_LH_DFPRQX9 port map( D => n2144, CP => clk, 
                           RN => n2803, Q => registers_23_6_port);
   registers_reg_23_5_inst : HS65_LH_DFPRQX9 port map( D => n2143, CP => clk, 
                           RN => n2803, Q => registers_23_5_port);
   registers_reg_23_4_inst : HS65_LH_DFPRQX9 port map( D => n2142, CP => clk, 
                           RN => n2803, Q => registers_23_4_port);
   registers_reg_23_3_inst : HS65_LH_DFPRQX9 port map( D => n2141, CP => clk, 
                           RN => n2803, Q => registers_23_3_port);
   registers_reg_23_2_inst : HS65_LH_DFPRQX9 port map( D => n2140, CP => clk, 
                           RN => n2803, Q => registers_23_2_port);
   registers_reg_23_1_inst : HS65_LH_DFPRQX9 port map( D => n2139, CP => clk, 
                           RN => n2803, Q => registers_23_1_port);
   registers_reg_23_0_inst : HS65_LH_DFPRQX9 port map( D => n2138, CP => clk, 
                           RN => n2803, Q => registers_23_0_port);
   registers_reg_22_31_inst : HS65_LH_DFPRQX9 port map( D => n2137, CP => clk, 
                           RN => n2803, Q => registers_22_31_port);
   registers_reg_22_30_inst : HS65_LH_DFPRQX9 port map( D => n2136, CP => clk, 
                           RN => n2802, Q => registers_22_30_port);
   registers_reg_22_29_inst : HS65_LH_DFPRQX9 port map( D => n2135, CP => clk, 
                           RN => n2802, Q => registers_22_29_port);
   registers_reg_22_28_inst : HS65_LH_DFPRQX9 port map( D => n2134, CP => clk, 
                           RN => n2802, Q => registers_22_28_port);
   registers_reg_22_27_inst : HS65_LH_DFPRQX9 port map( D => n2133, CP => clk, 
                           RN => n2802, Q => registers_22_27_port);
   registers_reg_22_26_inst : HS65_LH_DFPRQX9 port map( D => n2132, CP => clk, 
                           RN => n2802, Q => registers_22_26_port);
   registers_reg_22_25_inst : HS65_LH_DFPRQX9 port map( D => n2131, CP => clk, 
                           RN => n2802, Q => registers_22_25_port);
   registers_reg_22_24_inst : HS65_LH_DFPRQX9 port map( D => n2130, CP => clk, 
                           RN => n2802, Q => registers_22_24_port);
   registers_reg_22_23_inst : HS65_LH_DFPRQX9 port map( D => n2129, CP => clk, 
                           RN => n2802, Q => registers_22_23_port);
   registers_reg_22_22_inst : HS65_LH_DFPRQX9 port map( D => n2128, CP => clk, 
                           RN => n2802, Q => registers_22_22_port);
   registers_reg_22_21_inst : HS65_LH_DFPRQX9 port map( D => n2127, CP => clk, 
                           RN => n2802, Q => registers_22_21_port);
   registers_reg_22_20_inst : HS65_LH_DFPRQX9 port map( D => n2126, CP => clk, 
                           RN => n2802, Q => registers_22_20_port);
   registers_reg_22_19_inst : HS65_LH_DFPRQX9 port map( D => n2125, CP => clk, 
                           RN => n2802, Q => registers_22_19_port);
   registers_reg_22_18_inst : HS65_LH_DFPRQX9 port map( D => n2124, CP => clk, 
                           RN => n2801, Q => registers_22_18_port);
   registers_reg_22_17_inst : HS65_LH_DFPRQX9 port map( D => n2123, CP => clk, 
                           RN => n2801, Q => registers_22_17_port);
   registers_reg_22_16_inst : HS65_LH_DFPRQX9 port map( D => n2122, CP => clk, 
                           RN => n2801, Q => registers_22_16_port);
   registers_reg_22_15_inst : HS65_LH_DFPRQX9 port map( D => n2121, CP => clk, 
                           RN => n2801, Q => registers_22_15_port);
   registers_reg_22_14_inst : HS65_LH_DFPRQX9 port map( D => n2120, CP => clk, 
                           RN => n2801, Q => registers_22_14_port);
   registers_reg_22_13_inst : HS65_LH_DFPRQX9 port map( D => n2119, CP => clk, 
                           RN => n2801, Q => registers_22_13_port);
   registers_reg_22_12_inst : HS65_LH_DFPRQX9 port map( D => n2118, CP => clk, 
                           RN => n2801, Q => registers_22_12_port);
   registers_reg_22_11_inst : HS65_LH_DFPRQX9 port map( D => n2117, CP => clk, 
                           RN => n2801, Q => registers_22_11_port);
   registers_reg_22_10_inst : HS65_LH_DFPRQX9 port map( D => n2116, CP => clk, 
                           RN => n2801, Q => registers_22_10_port);
   registers_reg_22_9_inst : HS65_LH_DFPRQX9 port map( D => n2115, CP => clk, 
                           RN => n2801, Q => registers_22_9_port);
   registers_reg_22_8_inst : HS65_LH_DFPRQX9 port map( D => n2114, CP => clk, 
                           RN => n2801, Q => registers_22_8_port);
   registers_reg_22_7_inst : HS65_LH_DFPRQX9 port map( D => n2113, CP => clk, 
                           RN => n2808, Q => registers_22_7_port);
   registers_reg_22_6_inst : HS65_LH_DFPRQX9 port map( D => n2112, CP => clk, 
                           RN => n2825, Q => registers_22_6_port);
   registers_reg_22_5_inst : HS65_LH_DFPRQX9 port map( D => n2111, CP => clk, 
                           RN => n2825, Q => registers_22_5_port);
   registers_reg_22_4_inst : HS65_LH_DFPRQX9 port map( D => n2110, CP => clk, 
                           RN => n2825, Q => registers_22_4_port);
   registers_reg_22_3_inst : HS65_LH_DFPRQX9 port map( D => n2109, CP => clk, 
                           RN => n2825, Q => registers_22_3_port);
   registers_reg_22_2_inst : HS65_LH_DFPRQX9 port map( D => n2108, CP => clk, 
                           RN => n2825, Q => registers_22_2_port);
   registers_reg_22_1_inst : HS65_LH_DFPRQX9 port map( D => n2107, CP => clk, 
                           RN => n2825, Q => registers_22_1_port);
   registers_reg_22_0_inst : HS65_LH_DFPRQX9 port map( D => n2106, CP => clk, 
                           RN => n2825, Q => registers_22_0_port);
   registers_reg_21_31_inst : HS65_LH_DFPRQX9 port map( D => n2105, CP => clk, 
                           RN => n2825, Q => registers_21_31_port);
   registers_reg_21_30_inst : HS65_LH_DFPRQX9 port map( D => n2104, CP => clk, 
                           RN => n2826, Q => registers_21_30_port);
   registers_reg_21_29_inst : HS65_LH_DFPRQX9 port map( D => n2103, CP => clk, 
                           RN => n2825, Q => registers_21_29_port);
   registers_reg_21_28_inst : HS65_LH_DFPRQX9 port map( D => n2102, CP => clk, 
                           RN => n2826, Q => registers_21_28_port);
   registers_reg_21_27_inst : HS65_LH_DFPRQX9 port map( D => n2101, CP => clk, 
                           RN => n2825, Q => registers_21_27_port);
   registers_reg_21_26_inst : HS65_LH_DFPRQX9 port map( D => n2100, CP => clk, 
                           RN => n2826, Q => registers_21_26_port);
   registers_reg_21_25_inst : HS65_LH_DFPRQX9 port map( D => n2099, CP => clk, 
                           RN => n2825, Q => registers_21_25_port);
   registers_reg_21_24_inst : HS65_LH_DFPRQX9 port map( D => n2098, CP => clk, 
                           RN => n2826, Q => registers_21_24_port);
   registers_reg_21_23_inst : HS65_LH_DFPRQX9 port map( D => n2097, CP => clk, 
                           RN => n2825, Q => registers_21_23_port);
   registers_reg_21_22_inst : HS65_LH_DFPRQX9 port map( D => n2096, CP => clk, 
                           RN => n2824, Q => registers_21_22_port);
   registers_reg_21_21_inst : HS65_LH_DFPRQX9 port map( D => n2095, CP => clk, 
                           RN => n2824, Q => registers_21_21_port);
   registers_reg_21_20_inst : HS65_LH_DFPRQX9 port map( D => n2094, CP => clk, 
                           RN => n2824, Q => registers_21_20_port);
   registers_reg_21_19_inst : HS65_LH_DFPRQX9 port map( D => n2093, CP => clk, 
                           RN => n2824, Q => registers_21_19_port);
   registers_reg_21_18_inst : HS65_LH_DFPRQX9 port map( D => n2092, CP => clk, 
                           RN => n2824, Q => registers_21_18_port);
   registers_reg_21_17_inst : HS65_LH_DFPRQX9 port map( D => n2091, CP => clk, 
                           RN => n2824, Q => registers_21_17_port);
   registers_reg_21_16_inst : HS65_LH_DFPRQX9 port map( D => n2090, CP => clk, 
                           RN => n2824, Q => registers_21_16_port);
   registers_reg_21_15_inst : HS65_LH_DFPRQX9 port map( D => n2089, CP => clk, 
                           RN => n2824, Q => registers_21_15_port);
   registers_reg_21_14_inst : HS65_LH_DFPRQX9 port map( D => n2088, CP => clk, 
                           RN => n2824, Q => registers_21_14_port);
   registers_reg_21_13_inst : HS65_LH_DFPRQX9 port map( D => n2087, CP => clk, 
                           RN => n2824, Q => registers_21_13_port);
   registers_reg_21_12_inst : HS65_LH_DFPRQX9 port map( D => n2086, CP => clk, 
                           RN => n2824, Q => registers_21_12_port);
   registers_reg_21_11_inst : HS65_LH_DFPRQX9 port map( D => n2085, CP => clk, 
                           RN => n2824, Q => registers_21_11_port);
   registers_reg_21_10_inst : HS65_LH_DFPRQX9 port map( D => n2084, CP => clk, 
                           RN => n2823, Q => registers_21_10_port);
   registers_reg_21_9_inst : HS65_LH_DFPRQX9 port map( D => n2083, CP => clk, 
                           RN => n2823, Q => registers_21_9_port);
   registers_reg_21_8_inst : HS65_LH_DFPRQX9 port map( D => n2082, CP => clk, 
                           RN => n2823, Q => registers_21_8_port);
   registers_reg_21_7_inst : HS65_LH_DFPRQX9 port map( D => n2081, CP => clk, 
                           RN => n2823, Q => registers_21_7_port);
   registers_reg_21_6_inst : HS65_LH_DFPRQX9 port map( D => n2080, CP => clk, 
                           RN => n2823, Q => registers_21_6_port);
   registers_reg_21_5_inst : HS65_LH_DFPRQX9 port map( D => n2079, CP => clk, 
                           RN => n2823, Q => registers_21_5_port);
   registers_reg_21_4_inst : HS65_LH_DFPRQX9 port map( D => n2078, CP => clk, 
                           RN => n2823, Q => registers_21_4_port);
   registers_reg_21_3_inst : HS65_LH_DFPRQX9 port map( D => n2077, CP => clk, 
                           RN => n2823, Q => registers_21_3_port);
   registers_reg_21_2_inst : HS65_LH_DFPRQX9 port map( D => n2076, CP => clk, 
                           RN => n2823, Q => registers_21_2_port);
   registers_reg_21_1_inst : HS65_LH_DFPRQX9 port map( D => n2075, CP => clk, 
                           RN => n2823, Q => registers_21_1_port);
   registers_reg_21_0_inst : HS65_LH_DFPRQX9 port map( D => n2074, CP => clk, 
                           RN => n2823, Q => registers_21_0_port);
   registers_reg_20_31_inst : HS65_LH_DFPRQX9 port map( D => n2073, CP => clk, 
                           RN => n2823, Q => registers_20_31_port);
   registers_reg_20_30_inst : HS65_LH_DFPRQX9 port map( D => n2072, CP => clk, 
                           RN => n2816, Q => registers_20_30_port);
   registers_reg_20_29_inst : HS65_LH_DFPRQX9 port map( D => n2071, CP => clk, 
                           RN => n2816, Q => registers_20_29_port);
   registers_reg_20_28_inst : HS65_LH_DFPRQX9 port map( D => n2070, CP => clk, 
                           RN => n2816, Q => registers_20_28_port);
   registers_reg_20_27_inst : HS65_LH_DFPRQX9 port map( D => n2069, CP => clk, 
                           RN => n2816, Q => registers_20_27_port);
   registers_reg_20_26_inst : HS65_LH_DFPRQX9 port map( D => n2068, CP => clk, 
                           RN => n2816, Q => registers_20_26_port);
   registers_reg_20_25_inst : HS65_LH_DFPRQX9 port map( D => n2067, CP => clk, 
                           RN => n2816, Q => registers_20_25_port);
   registers_reg_20_24_inst : HS65_LH_DFPRQX9 port map( D => n2066, CP => clk, 
                           RN => n2816, Q => registers_20_24_port);
   registers_reg_20_23_inst : HS65_LH_DFPRQX9 port map( D => n2065, CP => clk, 
                           RN => n2816, Q => registers_20_23_port);
   registers_reg_20_22_inst : HS65_LH_DFPRQX9 port map( D => n2064, CP => clk, 
                           RN => n2817, Q => registers_20_22_port);
   registers_reg_20_21_inst : HS65_LH_DFPRQX9 port map( D => n2063, CP => clk, 
                           RN => n2821, Q => registers_20_21_port);
   registers_reg_20_20_inst : HS65_LH_DFPRQX9 port map( D => n2062, CP => clk, 
                           RN => n2817, Q => registers_20_20_port);
   registers_reg_20_19_inst : HS65_LH_DFPRQX9 port map( D => n2061, CP => clk, 
                           RN => n2817, Q => registers_20_19_port);
   registers_reg_20_18_inst : HS65_LH_DFPRQX9 port map( D => n2060, CP => clk, 
                           RN => n2817, Q => registers_20_18_port);
   registers_reg_20_17_inst : HS65_LH_DFPRQX9 port map( D => n2059, CP => clk, 
                           RN => n2817, Q => registers_20_17_port);
   registers_reg_20_16_inst : HS65_LH_DFPRQX9 port map( D => n2058, CP => clk, 
                           RN => n2817, Q => registers_20_16_port);
   registers_reg_20_15_inst : HS65_LH_DFPRQX9 port map( D => n2057, CP => clk, 
                           RN => n2817, Q => registers_20_15_port);
   registers_reg_20_14_inst : HS65_LH_DFPRQX9 port map( D => n2056, CP => clk, 
                           RN => n2817, Q => registers_20_14_port);
   registers_reg_20_13_inst : HS65_LH_DFPRQX9 port map( D => n2055, CP => clk, 
                           RN => n2817, Q => registers_20_13_port);
   registers_reg_20_12_inst : HS65_LH_DFPRQX9 port map( D => n2054, CP => clk, 
                           RN => n2817, Q => registers_20_12_port);
   registers_reg_20_11_inst : HS65_LH_DFPRQX9 port map( D => n2053, CP => clk, 
                           RN => n2817, Q => registers_20_11_port);
   registers_reg_20_10_inst : HS65_LH_DFPRQX9 port map( D => n2052, CP => clk, 
                           RN => n2818, Q => registers_20_10_port);
   registers_reg_20_9_inst : HS65_LH_DFPRQX9 port map( D => n2051, CP => clk, 
                           RN => n2818, Q => registers_20_9_port);
   registers_reg_20_8_inst : HS65_LH_DFPRQX9 port map( D => n2050, CP => clk, 
                           RN => n2818, Q => registers_20_8_port);
   registers_reg_20_7_inst : HS65_LH_DFPRQX9 port map( D => n2049, CP => clk, 
                           RN => n2818, Q => registers_20_7_port);
   registers_reg_20_6_inst : HS65_LH_DFPRQX9 port map( D => n2048, CP => clk, 
                           RN => n2818, Q => registers_20_6_port);
   registers_reg_20_5_inst : HS65_LH_DFPRQX9 port map( D => n2047, CP => clk, 
                           RN => n2818, Q => registers_20_5_port);
   registers_reg_20_4_inst : HS65_LH_DFPRQX9 port map( D => n2046, CP => clk, 
                           RN => n2818, Q => registers_20_4_port);
   registers_reg_20_3_inst : HS65_LH_DFPRQX9 port map( D => n2045, CP => clk, 
                           RN => n2818, Q => registers_20_3_port);
   registers_reg_20_2_inst : HS65_LH_DFPRQX9 port map( D => n2044, CP => clk, 
                           RN => n2818, Q => registers_20_2_port);
   registers_reg_20_1_inst : HS65_LH_DFPRQX9 port map( D => n2043, CP => clk, 
                           RN => n2818, Q => registers_20_1_port);
   registers_reg_20_0_inst : HS65_LH_DFPRQX9 port map( D => n2042, CP => clk, 
                           RN => n2818, Q => registers_20_0_port);
   registers_reg_19_31_inst : HS65_LH_DFPRQX9 port map( D => n2041, CP => clk, 
                           RN => n2819, Q => registers_19_31_port);
   registers_reg_19_30_inst : HS65_LH_DFPRQX9 port map( D => n2040, CP => clk, 
                           RN => n2819, Q => registers_19_30_port);
   registers_reg_19_29_inst : HS65_LH_DFPRQX9 port map( D => n2039, CP => clk, 
                           RN => n2819, Q => registers_19_29_port);
   registers_reg_19_28_inst : HS65_LH_DFPRQX9 port map( D => n2038, CP => clk, 
                           RN => n2819, Q => registers_19_28_port);
   registers_reg_19_27_inst : HS65_LH_DFPRQX9 port map( D => n2037, CP => clk, 
                           RN => n2819, Q => registers_19_27_port);
   registers_reg_19_26_inst : HS65_LH_DFPRQX9 port map( D => n2036, CP => clk, 
                           RN => n2819, Q => registers_19_26_port);
   registers_reg_19_25_inst : HS65_LH_DFPRQX9 port map( D => n2035, CP => clk, 
                           RN => n2819, Q => registers_19_25_port);
   registers_reg_19_24_inst : HS65_LH_DFPRQX9 port map( D => n2034, CP => clk, 
                           RN => n2819, Q => registers_19_24_port);
   registers_reg_19_23_inst : HS65_LH_DFPRQX9 port map( D => n2033, CP => clk, 
                           RN => n2819, Q => registers_19_23_port);
   registers_reg_19_22_inst : HS65_LH_DFPRQX9 port map( D => n2032, CP => clk, 
                           RN => n2819, Q => registers_19_22_port);
   registers_reg_19_21_inst : HS65_LH_DFPRQX9 port map( D => n2031, CP => clk, 
                           RN => n2819, Q => registers_19_21_port);
   registers_reg_19_20_inst : HS65_LH_DFPRQX9 port map( D => n2030, CP => clk, 
                           RN => n2819, Q => registers_19_20_port);
   registers_reg_19_19_inst : HS65_LH_DFPRQX9 port map( D => n2029, CP => clk, 
                           RN => n2820, Q => registers_19_19_port);
   registers_reg_19_18_inst : HS65_LH_DFPRQX9 port map( D => n2028, CP => clk, 
                           RN => n2820, Q => registers_19_18_port);
   registers_reg_19_17_inst : HS65_LH_DFPRQX9 port map( D => n2027, CP => clk, 
                           RN => n2820, Q => registers_19_17_port);
   registers_reg_19_16_inst : HS65_LH_DFPRQX9 port map( D => n2026, CP => clk, 
                           RN => n2820, Q => registers_19_16_port);
   registers_reg_19_15_inst : HS65_LH_DFPRQX9 port map( D => n2025, CP => clk, 
                           RN => n2820, Q => registers_19_15_port);
   registers_reg_19_14_inst : HS65_LH_DFPRQX9 port map( D => n2024, CP => clk, 
                           RN => n2820, Q => registers_19_14_port);
   registers_reg_19_13_inst : HS65_LH_DFPRQX9 port map( D => n2023, CP => clk, 
                           RN => n2820, Q => registers_19_13_port);
   registers_reg_19_12_inst : HS65_LH_DFPRQX9 port map( D => n2022, CP => clk, 
                           RN => n2820, Q => registers_19_12_port);
   registers_reg_19_11_inst : HS65_LH_DFPRQX9 port map( D => n2021, CP => clk, 
                           RN => n2820, Q => registers_19_11_port);
   registers_reg_19_10_inst : HS65_LH_DFPRQX9 port map( D => n2020, CP => clk, 
                           RN => n2820, Q => registers_19_10_port);
   registers_reg_19_9_inst : HS65_LH_DFPRQX9 port map( D => n2019, CP => clk, 
                           RN => n2820, Q => registers_19_9_port);
   registers_reg_19_8_inst : HS65_LH_DFPRQX9 port map( D => n2018, CP => clk, 
                           RN => n2820, Q => registers_19_8_port);
   registers_reg_19_7_inst : HS65_LH_DFPRQX9 port map( D => n2017, CP => clk, 
                           RN => n2821, Q => registers_19_7_port);
   registers_reg_19_6_inst : HS65_LH_DFPRQX9 port map( D => n2016, CP => clk, 
                           RN => n2821, Q => registers_19_6_port);
   registers_reg_19_5_inst : HS65_LH_DFPRQX9 port map( D => n2015, CP => clk, 
                           RN => n2821, Q => registers_19_5_port);
   registers_reg_19_4_inst : HS65_LH_DFPRQX9 port map( D => n2014, CP => clk, 
                           RN => n2821, Q => registers_19_4_port);
   registers_reg_19_3_inst : HS65_LH_DFPRQX9 port map( D => n2013, CP => clk, 
                           RN => n2821, Q => registers_19_3_port);
   registers_reg_19_2_inst : HS65_LH_DFPRQX9 port map( D => n2012, CP => clk, 
                           RN => n2821, Q => registers_19_2_port);
   registers_reg_19_1_inst : HS65_LH_DFPRQX9 port map( D => n2011, CP => clk, 
                           RN => n2821, Q => registers_19_1_port);
   registers_reg_19_0_inst : HS65_LH_DFPRQX9 port map( D => n2010, CP => clk, 
                           RN => n2821, Q => registers_19_0_port);
   registers_reg_18_31_inst : HS65_LH_DFPRQX9 port map( D => n2009, CP => clk, 
                           RN => n2821, Q => registers_18_31_port);
   registers_reg_18_30_inst : HS65_LH_DFPRQX9 port map( D => n2008, CP => clk, 
                           RN => n2821, Q => registers_18_30_port);
   registers_reg_18_29_inst : HS65_LH_DFPRQX9 port map( D => n2007, CP => clk, 
                           RN => n2821, Q => registers_18_29_port);
   registers_reg_18_28_inst : HS65_LH_DFPRQX9 port map( D => n2006, CP => clk, 
                           RN => n2822, Q => registers_18_28_port);
   registers_reg_18_27_inst : HS65_LH_DFPRQX9 port map( D => n2005, CP => clk, 
                           RN => n2822, Q => registers_18_27_port);
   registers_reg_18_26_inst : HS65_LH_DFPRQX9 port map( D => n2004, CP => clk, 
                           RN => n2822, Q => registers_18_26_port);
   registers_reg_18_25_inst : HS65_LH_DFPRQX9 port map( D => n2003, CP => clk, 
                           RN => n2822, Q => registers_18_25_port);
   registers_reg_18_24_inst : HS65_LH_DFPRQX9 port map( D => n2002, CP => clk, 
                           RN => n2822, Q => registers_18_24_port);
   registers_reg_18_23_inst : HS65_LH_DFPRQX9 port map( D => n2001, CP => clk, 
                           RN => n2822, Q => registers_18_23_port);
   registers_reg_18_22_inst : HS65_LH_DFPRQX9 port map( D => n2000, CP => clk, 
                           RN => n2822, Q => registers_18_22_port);
   registers_reg_18_21_inst : HS65_LH_DFPRQX9 port map( D => n1999, CP => clk, 
                           RN => n2822, Q => registers_18_21_port);
   registers_reg_18_20_inst : HS65_LH_DFPRQX9 port map( D => n1998, CP => clk, 
                           RN => n2822, Q => registers_18_20_port);
   registers_reg_18_19_inst : HS65_LH_DFPRQX9 port map( D => n1997, CP => clk, 
                           RN => n2822, Q => registers_18_19_port);
   registers_reg_18_18_inst : HS65_LH_DFPRQX9 port map( D => n1996, CP => clk, 
                           RN => n2822, Q => registers_18_18_port);
   registers_reg_18_17_inst : HS65_LH_DFPRQX9 port map( D => n1995, CP => clk, 
                           RN => n2822, Q => registers_18_17_port);
   registers_reg_18_16_inst : HS65_LH_DFPRQX9 port map( D => n1994, CP => clk, 
                           RN => n2818, Q => registers_18_16_port);
   registers_reg_18_15_inst : HS65_LH_DFPRQX9 port map( D => n1993, CP => clk, 
                           RN => n2783, Q => registers_18_15_port);
   registers_reg_18_14_inst : HS65_LH_DFPRQX9 port map( D => n1992, CP => clk, 
                           RN => n2778, Q => registers_18_14_port);
   registers_reg_18_13_inst : HS65_LH_DFPRQX9 port map( D => n1991, CP => clk, 
                           RN => n2774, Q => registers_18_13_port);
   registers_reg_18_12_inst : HS65_LH_DFPRQX9 port map( D => n1990, CP => clk, 
                           RN => n2774, Q => registers_18_12_port);
   registers_reg_18_11_inst : HS65_LH_DFPRQX9 port map( D => n1989, CP => clk, 
                           RN => n2774, Q => registers_18_11_port);
   registers_reg_18_10_inst : HS65_LH_DFPRQX9 port map( D => n1988, CP => clk, 
                           RN => n2774, Q => registers_18_10_port);
   registers_reg_18_9_inst : HS65_LH_DFPRQX9 port map( D => n1987, CP => clk, 
                           RN => n2774, Q => registers_18_9_port);
   registers_reg_18_8_inst : HS65_LH_DFPRQX9 port map( D => n1986, CP => clk, 
                           RN => n2774, Q => registers_18_8_port);
   registers_reg_18_7_inst : HS65_LH_DFPRQX9 port map( D => n1985, CP => clk, 
                           RN => n2774, Q => registers_18_7_port);
   registers_reg_18_6_inst : HS65_LH_DFPRQX9 port map( D => n1984, CP => clk, 
                           RN => n2774, Q => registers_18_6_port);
   registers_reg_18_5_inst : HS65_LH_DFPRQX9 port map( D => n1983, CP => clk, 
                           RN => n2774, Q => registers_18_5_port);
   registers_reg_18_4_inst : HS65_LH_DFPRQX9 port map( D => n1982, CP => clk, 
                           RN => n2774, Q => registers_18_4_port);
   registers_reg_18_3_inst : HS65_LH_DFPRQX9 port map( D => n1981, CP => clk, 
                           RN => n2774, Q => registers_18_3_port);
   registers_reg_18_2_inst : HS65_LH_DFPRQX9 port map( D => n1980, CP => clk, 
                           RN => n2775, Q => registers_18_2_port);
   registers_reg_18_1_inst : HS65_LH_DFPRQX9 port map( D => n1979, CP => clk, 
                           RN => n2775, Q => registers_18_1_port);
   registers_reg_18_0_inst : HS65_LH_DFPRQX9 port map( D => n1978, CP => clk, 
                           RN => n2775, Q => registers_18_0_port);
   registers_reg_17_31_inst : HS65_LH_DFPRQX9 port map( D => n1977, CP => clk, 
                           RN => n2775, Q => registers_17_31_port);
   registers_reg_17_30_inst : HS65_LH_DFPRQX9 port map( D => n1976, CP => clk, 
                           RN => n2775, Q => registers_17_30_port);
   registers_reg_17_29_inst : HS65_LH_DFPRQX9 port map( D => n1975, CP => clk, 
                           RN => n2775, Q => registers_17_29_port);
   registers_reg_17_28_inst : HS65_LH_DFPRQX9 port map( D => n1974, CP => clk, 
                           RN => n2775, Q => registers_17_28_port);
   registers_reg_17_27_inst : HS65_LH_DFPRQX9 port map( D => n1973, CP => clk, 
                           RN => n2775, Q => registers_17_27_port);
   registers_reg_17_26_inst : HS65_LH_DFPRQX9 port map( D => n1972, CP => clk, 
                           RN => n2775, Q => registers_17_26_port);
   registers_reg_17_25_inst : HS65_LH_DFPRQX9 port map( D => n1971, CP => clk, 
                           RN => n2775, Q => registers_17_25_port);
   registers_reg_17_24_inst : HS65_LH_DFPRQX9 port map( D => n1970, CP => clk, 
                           RN => n2775, Q => registers_17_24_port);
   registers_reg_17_23_inst : HS65_LH_DFPRQX9 port map( D => n1969, CP => clk, 
                           RN => n2775, Q => registers_17_23_port);
   registers_reg_17_22_inst : HS65_LH_DFPRQX9 port map( D => n1968, CP => clk, 
                           RN => n2776, Q => registers_17_22_port);
   registers_reg_17_21_inst : HS65_LH_DFPRQX9 port map( D => n1967, CP => clk, 
                           RN => n2776, Q => registers_17_21_port);
   registers_reg_17_20_inst : HS65_LH_DFPRQX9 port map( D => n1966, CP => clk, 
                           RN => n2776, Q => registers_17_20_port);
   registers_reg_17_19_inst : HS65_LH_DFPRQX9 port map( D => n1965, CP => clk, 
                           RN => n2776, Q => registers_17_19_port);
   registers_reg_17_18_inst : HS65_LH_DFPRQX9 port map( D => n1964, CP => clk, 
                           RN => n2776, Q => registers_17_18_port);
   registers_reg_17_17_inst : HS65_LH_DFPRQX9 port map( D => n1963, CP => clk, 
                           RN => n2776, Q => registers_17_17_port);
   registers_reg_17_16_inst : HS65_LH_DFPRQX9 port map( D => n1962, CP => clk, 
                           RN => n2776, Q => registers_17_16_port);
   registers_reg_17_15_inst : HS65_LH_DFPRQX9 port map( D => n1961, CP => clk, 
                           RN => n2776, Q => registers_17_15_port);
   registers_reg_17_14_inst : HS65_LH_DFPRQX9 port map( D => n1960, CP => clk, 
                           RN => n2776, Q => registers_17_14_port);
   registers_reg_17_13_inst : HS65_LH_DFPRQX9 port map( D => n1959, CP => clk, 
                           RN => n2776, Q => registers_17_13_port);
   registers_reg_17_12_inst : HS65_LH_DFPRQX9 port map( D => n1958, CP => clk, 
                           RN => n2776, Q => registers_17_12_port);
   registers_reg_17_11_inst : HS65_LH_DFPRQX9 port map( D => n1957, CP => clk, 
                           RN => n2776, Q => registers_17_11_port);
   registers_reg_17_10_inst : HS65_LH_DFPRQX9 port map( D => n1956, CP => clk, 
                           RN => n2777, Q => registers_17_10_port);
   registers_reg_17_9_inst : HS65_LH_DFPRQX9 port map( D => n1955, CP => clk, 
                           RN => n2777, Q => registers_17_9_port);
   registers_reg_17_8_inst : HS65_LH_DFPRQX9 port map( D => n1954, CP => clk, 
                           RN => n2777, Q => registers_17_8_port);
   registers_reg_17_7_inst : HS65_LH_DFPRQX9 port map( D => n1953, CP => clk, 
                           RN => n2777, Q => registers_17_7_port);
   registers_reg_17_6_inst : HS65_LH_DFPRQX9 port map( D => n1952, CP => clk, 
                           RN => n2777, Q => registers_17_6_port);
   registers_reg_17_5_inst : HS65_LH_DFPRQX9 port map( D => n1951, CP => clk, 
                           RN => n2777, Q => registers_17_5_port);
   registers_reg_17_4_inst : HS65_LH_DFPRQX9 port map( D => n1950, CP => clk, 
                           RN => n2777, Q => registers_17_4_port);
   registers_reg_17_3_inst : HS65_LH_DFPRQX9 port map( D => n1949, CP => clk, 
                           RN => n2777, Q => registers_17_3_port);
   registers_reg_17_2_inst : HS65_LH_DFPRQX9 port map( D => n1948, CP => clk, 
                           RN => n2777, Q => registers_17_2_port);
   registers_reg_17_1_inst : HS65_LH_DFPRQX9 port map( D => n1947, CP => clk, 
                           RN => n2777, Q => registers_17_1_port);
   registers_reg_17_0_inst : HS65_LH_DFPRQX9 port map( D => n1946, CP => clk, 
                           RN => n2777, Q => registers_17_0_port);
   registers_reg_16_31_inst : HS65_LH_DFPRQX9 port map( D => n1945, CP => clk, 
                           RN => n2777, Q => registers_16_31_port);
   registers_reg_16_30_inst : HS65_LH_DFPRQX9 port map( D => n1944, CP => clk, 
                           RN => n2778, Q => registers_16_30_port);
   registers_reg_16_29_inst : HS65_LH_DFPRQX9 port map( D => n1943, CP => clk, 
                           RN => n2778, Q => registers_16_29_port);
   registers_reg_16_28_inst : HS65_LH_DFPRQX9 port map( D => n1942, CP => clk, 
                           RN => n2778, Q => registers_16_28_port);
   registers_reg_16_27_inst : HS65_LH_DFPRQX9 port map( D => n1941, CP => clk, 
                           RN => n2778, Q => registers_16_27_port);
   registers_reg_16_26_inst : HS65_LH_DFPRQX9 port map( D => n1940, CP => clk, 
                           RN => n2778, Q => registers_16_26_port);
   registers_reg_16_25_inst : HS65_LH_DFPRQX9 port map( D => n1939, CP => clk, 
                           RN => n2778, Q => registers_16_25_port);
   registers_reg_16_24_inst : HS65_LH_DFPRQX9 port map( D => n1938, CP => clk, 
                           RN => n2778, Q => registers_16_24_port);
   registers_reg_16_23_inst : HS65_LH_DFPRQX9 port map( D => n1937, CP => clk, 
                           RN => n2778, Q => registers_16_23_port);
   registers_reg_16_22_inst : HS65_LH_DFPRQX9 port map( D => n1936, CP => clk, 
                           RN => n2778, Q => registers_16_22_port);
   registers_reg_16_21_inst : HS65_LH_DFPRQX9 port map( D => n1935, CP => clk, 
                           RN => n2778, Q => registers_16_21_port);
   registers_reg_16_20_inst : HS65_LH_DFPRQX9 port map( D => n1934, CP => clk, 
                           RN => n2778, Q => registers_16_20_port);
   registers_reg_16_19_inst : HS65_LH_DFPRQX9 port map( D => n1933, CP => clk, 
                           RN => n2779, Q => registers_16_19_port);
   registers_reg_16_18_inst : HS65_LH_DFPRQX9 port map( D => n1932, CP => clk, 
                           RN => n2779, Q => registers_16_18_port);
   registers_reg_16_17_inst : HS65_LH_DFPRQX9 port map( D => n1931, CP => clk, 
                           RN => n2779, Q => registers_16_17_port);
   registers_reg_16_16_inst : HS65_LH_DFPRQX9 port map( D => n1930, CP => clk, 
                           RN => n2779, Q => registers_16_16_port);
   registers_reg_16_15_inst : HS65_LH_DFPRQX9 port map( D => n1929, CP => clk, 
                           RN => n2779, Q => registers_16_15_port);
   registers_reg_16_14_inst : HS65_LH_DFPRQX9 port map( D => n1928, CP => clk, 
                           RN => n2779, Q => registers_16_14_port);
   registers_reg_16_13_inst : HS65_LH_DFPRQX9 port map( D => n1927, CP => clk, 
                           RN => n2779, Q => registers_16_13_port);
   registers_reg_16_12_inst : HS65_LH_DFPRQX9 port map( D => n1926, CP => clk, 
                           RN => n2779, Q => registers_16_12_port);
   registers_reg_16_11_inst : HS65_LH_DFPRQX9 port map( D => n1925, CP => clk, 
                           RN => n2779, Q => registers_16_11_port);
   registers_reg_16_10_inst : HS65_LH_DFPRQX9 port map( D => n1924, CP => clk, 
                           RN => n2779, Q => registers_16_10_port);
   registers_reg_16_9_inst : HS65_LH_DFPRQX9 port map( D => n1923, CP => clk, 
                           RN => n2779, Q => registers_16_9_port);
   registers_reg_16_8_inst : HS65_LH_DFPRQX9 port map( D => n1922, CP => clk, 
                           RN => n2779, Q => registers_16_8_port);
   registers_reg_16_7_inst : HS65_LH_DFPRQX9 port map( D => n1921, CP => clk, 
                           RN => n2780, Q => registers_16_7_port);
   registers_reg_16_6_inst : HS65_LH_DFPRQX9 port map( D => n1920, CP => clk, 
                           RN => n2780, Q => registers_16_6_port);
   registers_reg_16_5_inst : HS65_LH_DFPRQX9 port map( D => n1919, CP => clk, 
                           RN => n2780, Q => registers_16_5_port);
   registers_reg_16_4_inst : HS65_LH_DFPRQX9 port map( D => n1918, CP => clk, 
                           RN => n2780, Q => registers_16_4_port);
   registers_reg_16_3_inst : HS65_LH_DFPRQX9 port map( D => n1917, CP => clk, 
                           RN => n2780, Q => registers_16_3_port);
   registers_reg_16_2_inst : HS65_LH_DFPRQX9 port map( D => n1916, CP => clk, 
                           RN => n2780, Q => registers_16_2_port);
   registers_reg_16_1_inst : HS65_LH_DFPRQX9 port map( D => n1915, CP => clk, 
                           RN => n2780, Q => registers_16_1_port);
   registers_reg_16_0_inst : HS65_LH_DFPRQX9 port map( D => n1914, CP => clk, 
                           RN => n2780, Q => registers_16_0_port);
   registers_reg_13_31_inst : HS65_LH_DFPRQX9 port map( D => n1849, CP => clk, 
                           RN => n2780, Q => registers_13_31_port);
   registers_reg_13_30_inst : HS65_LH_DFPRQX9 port map( D => n1848, CP => clk, 
                           RN => n2780, Q => registers_13_30_port);
   registers_reg_13_29_inst : HS65_LH_DFPRQX9 port map( D => n1847, CP => clk, 
                           RN => n2780, Q => registers_13_29_port);
   registers_reg_13_28_inst : HS65_LH_DFPRQX9 port map( D => n1846, CP => clk, 
                           RN => n2780, Q => registers_13_28_port);
   registers_reg_13_27_inst : HS65_LH_DFPRQX9 port map( D => n1845, CP => clk, 
                           RN => n2781, Q => registers_13_27_port);
   registers_reg_13_26_inst : HS65_LH_DFPRQX9 port map( D => n1844, CP => clk, 
                           RN => n2781, Q => registers_13_26_port);
   registers_reg_13_25_inst : HS65_LH_DFPRQX9 port map( D => n1843, CP => clk, 
                           RN => n2781, Q => registers_13_25_port);
   registers_reg_13_24_inst : HS65_LH_DFPRQX9 port map( D => n1842, CP => clk, 
                           RN => n2781, Q => registers_13_24_port);
   registers_reg_13_23_inst : HS65_LH_DFPRQX9 port map( D => n1841, CP => clk, 
                           RN => n2781, Q => registers_13_23_port);
   registers_reg_13_22_inst : HS65_LH_DFPRQX9 port map( D => n1840, CP => clk, 
                           RN => n2781, Q => registers_13_22_port);
   registers_reg_13_21_inst : HS65_LH_DFPRQX9 port map( D => n1839, CP => clk, 
                           RN => n2781, Q => registers_13_21_port);
   registers_reg_13_20_inst : HS65_LH_DFPRQX9 port map( D => n1838, CP => clk, 
                           RN => n2781, Q => registers_13_20_port);
   registers_reg_13_19_inst : HS65_LH_DFPRQX9 port map( D => n1837, CP => clk, 
                           RN => n2781, Q => registers_13_19_port);
   registers_reg_13_18_inst : HS65_LH_DFPRQX9 port map( D => n1836, CP => clk, 
                           RN => n2781, Q => registers_13_18_port);
   registers_reg_13_17_inst : HS65_LH_DFPRQX9 port map( D => n1835, CP => clk, 
                           RN => n2781, Q => registers_13_17_port);
   registers_reg_13_16_inst : HS65_LH_DFPRQX9 port map( D => n1834, CP => clk, 
                           RN => n2781, Q => registers_13_16_port);
   registers_reg_13_15_inst : HS65_LH_DFPRQX9 port map( D => n1833, CP => clk, 
                           RN => n2782, Q => registers_13_15_port);
   registers_reg_13_14_inst : HS65_LH_DFPRQX9 port map( D => n1832, CP => clk, 
                           RN => n2782, Q => registers_13_14_port);
   registers_reg_13_13_inst : HS65_LH_DFPRQX9 port map( D => n1831, CP => clk, 
                           RN => n2782, Q => registers_13_13_port);
   registers_reg_13_12_inst : HS65_LH_DFPRQX9 port map( D => n1830, CP => clk, 
                           RN => n2782, Q => registers_13_12_port);
   registers_reg_13_11_inst : HS65_LH_DFPRQX9 port map( D => n1829, CP => clk, 
                           RN => n2782, Q => registers_13_11_port);
   registers_reg_13_10_inst : HS65_LH_DFPRQX9 port map( D => n1828, CP => clk, 
                           RN => n2782, Q => registers_13_10_port);
   registers_reg_13_9_inst : HS65_LH_DFPRQX9 port map( D => n1827, CP => clk, 
                           RN => n2782, Q => registers_13_9_port);
   registers_reg_13_8_inst : HS65_LH_DFPRQX9 port map( D => n1826, CP => clk, 
                           RN => n2782, Q => registers_13_8_port);
   registers_reg_13_7_inst : HS65_LH_DFPRQX9 port map( D => n1825, CP => clk, 
                           RN => n2782, Q => registers_13_7_port);
   registers_reg_13_6_inst : HS65_LH_DFPRQX9 port map( D => n1824, CP => clk, 
                           RN => n2782, Q => registers_13_6_port);
   registers_reg_13_5_inst : HS65_LH_DFPRQX9 port map( D => n1823, CP => clk, 
                           RN => n2782, Q => registers_13_5_port);
   registers_reg_13_4_inst : HS65_LH_DFPRQX9 port map( D => n1822, CP => clk, 
                           RN => n2782, Q => registers_13_4_port);
   registers_reg_13_3_inst : HS65_LH_DFPRQX9 port map( D => n1821, CP => clk, 
                           RN => n2769, Q => registers_13_3_port);
   registers_reg_13_2_inst : HS65_LH_DFPRQX9 port map( D => n1820, CP => clk, 
                           RN => n2765, Q => registers_13_2_port);
   registers_reg_13_1_inst : HS65_LH_DFPRQX9 port map( D => n1819, CP => clk, 
                           RN => n2765, Q => registers_13_1_port);
   registers_reg_13_0_inst : HS65_LH_DFPRQX9 port map( D => n1818, CP => clk, 
                           RN => n2765, Q => registers_13_0_port);
   registers_reg_12_31_inst : HS65_LH_DFPRQX9 port map( D => n1817, CP => clk, 
                           RN => n2765, Q => registers_12_31_port);
   registers_reg_12_30_inst : HS65_LH_DFPRQX9 port map( D => n1816, CP => clk, 
                           RN => n2765, Q => registers_12_30_port);
   registers_reg_12_29_inst : HS65_LH_DFPRQX9 port map( D => n1815, CP => clk, 
                           RN => n2765, Q => registers_12_29_port);
   registers_reg_12_28_inst : HS65_LH_DFPRQX9 port map( D => n1814, CP => clk, 
                           RN => n2765, Q => registers_12_28_port);
   registers_reg_12_27_inst : HS65_LH_DFPRQX9 port map( D => n1813, CP => clk, 
                           RN => n2765, Q => registers_12_27_port);
   registers_reg_12_26_inst : HS65_LH_DFPRQX9 port map( D => n1812, CP => clk, 
                           RN => n2765, Q => registers_12_26_port);
   registers_reg_12_25_inst : HS65_LH_DFPRQX9 port map( D => n1811, CP => clk, 
                           RN => n2765, Q => registers_12_25_port);
   registers_reg_12_24_inst : HS65_LH_DFPRQX9 port map( D => n1810, CP => clk, 
                           RN => n2765, Q => registers_12_24_port);
   registers_reg_12_23_inst : HS65_LH_DFPRQX9 port map( D => n1809, CP => clk, 
                           RN => n2766, Q => registers_12_23_port);
   registers_reg_12_22_inst : HS65_LH_DFPRQX9 port map( D => n1808, CP => clk, 
                           RN => n2766, Q => registers_12_22_port);
   registers_reg_12_21_inst : HS65_LH_DFPRQX9 port map( D => n1807, CP => clk, 
                           RN => n2766, Q => registers_12_21_port);
   registers_reg_12_20_inst : HS65_LH_DFPRQX9 port map( D => n1806, CP => clk, 
                           RN => n2766, Q => registers_12_20_port);
   registers_reg_12_19_inst : HS65_LH_DFPRQX9 port map( D => n1805, CP => clk, 
                           RN => n2766, Q => registers_12_19_port);
   registers_reg_12_18_inst : HS65_LH_DFPRQX9 port map( D => n1804, CP => clk, 
                           RN => n2766, Q => registers_12_18_port);
   registers_reg_12_17_inst : HS65_LH_DFPRQX9 port map( D => n1803, CP => clk, 
                           RN => n2766, Q => registers_12_17_port);
   registers_reg_12_16_inst : HS65_LH_DFPRQX9 port map( D => n1802, CP => clk, 
                           RN => n2766, Q => registers_12_16_port);
   registers_reg_12_15_inst : HS65_LH_DFPRQX9 port map( D => n1801, CP => clk, 
                           RN => n2766, Q => registers_12_15_port);
   registers_reg_12_14_inst : HS65_LH_DFPRQX9 port map( D => n1800, CP => clk, 
                           RN => n2766, Q => registers_12_14_port);
   registers_reg_12_13_inst : HS65_LH_DFPRQX9 port map( D => n1799, CP => clk, 
                           RN => n2766, Q => registers_12_13_port);
   registers_reg_12_12_inst : HS65_LH_DFPRQX9 port map( D => n1798, CP => clk, 
                           RN => n2766, Q => registers_12_12_port);
   registers_reg_12_11_inst : HS65_LH_DFPRQX9 port map( D => n1797, CP => clk, 
                           RN => n2767, Q => registers_12_11_port);
   registers_reg_12_10_inst : HS65_LH_DFPRQX9 port map( D => n1796, CP => clk, 
                           RN => n2767, Q => registers_12_10_port);
   registers_reg_12_9_inst : HS65_LH_DFPRQX9 port map( D => n1795, CP => clk, 
                           RN => n2767, Q => registers_12_9_port);
   registers_reg_12_8_inst : HS65_LH_DFPRQX9 port map( D => n1794, CP => clk, 
                           RN => n2767, Q => registers_12_8_port);
   registers_reg_12_7_inst : HS65_LH_DFPRQX9 port map( D => n1793, CP => clk, 
                           RN => n2767, Q => registers_12_7_port);
   registers_reg_12_6_inst : HS65_LH_DFPRQX9 port map( D => n1792, CP => clk, 
                           RN => n2767, Q => registers_12_6_port);
   registers_reg_12_5_inst : HS65_LH_DFPRQX9 port map( D => n1791, CP => clk, 
                           RN => n2767, Q => registers_12_5_port);
   registers_reg_12_4_inst : HS65_LH_DFPRQX9 port map( D => n1790, CP => clk, 
                           RN => n2767, Q => registers_12_4_port);
   registers_reg_12_3_inst : HS65_LH_DFPRQX9 port map( D => n1789, CP => clk, 
                           RN => n2767, Q => registers_12_3_port);
   registers_reg_12_2_inst : HS65_LH_DFPRQX9 port map( D => n1788, CP => clk, 
                           RN => n2767, Q => registers_12_2_port);
   registers_reg_12_1_inst : HS65_LH_DFPRQX9 port map( D => n1787, CP => clk, 
                           RN => n2767, Q => registers_12_1_port);
   registers_reg_12_0_inst : HS65_LH_DFPRQX9 port map( D => n1786, CP => clk, 
                           RN => n2767, Q => registers_12_0_port);
   registers_reg_11_31_inst : HS65_LH_DFPRQX9 port map( D => n1785, CP => clk, 
                           RN => n2768, Q => registers_11_31_port);
   registers_reg_11_30_inst : HS65_LH_DFPRQX9 port map( D => n1784, CP => clk, 
                           RN => n2768, Q => registers_11_30_port);
   registers_reg_11_29_inst : HS65_LH_DFPRQX9 port map( D => n1783, CP => clk, 
                           RN => n2768, Q => registers_11_29_port);
   registers_reg_11_28_inst : HS65_LH_DFPRQX9 port map( D => n1782, CP => clk, 
                           RN => n2768, Q => registers_11_28_port);
   registers_reg_11_27_inst : HS65_LH_DFPRQX9 port map( D => n1781, CP => clk, 
                           RN => n2768, Q => registers_11_27_port);
   registers_reg_11_26_inst : HS65_LH_DFPRQX9 port map( D => n1780, CP => clk, 
                           RN => n2768, Q => registers_11_26_port);
   registers_reg_11_25_inst : HS65_LH_DFPRQX9 port map( D => n1779, CP => clk, 
                           RN => n2768, Q => registers_11_25_port);
   registers_reg_11_24_inst : HS65_LH_DFPRQX9 port map( D => n1778, CP => clk, 
                           RN => n2768, Q => registers_11_24_port);
   registers_reg_11_23_inst : HS65_LH_DFPRQX9 port map( D => n1777, CP => clk, 
                           RN => n2768, Q => registers_11_23_port);
   registers_reg_11_22_inst : HS65_LH_DFPRQX9 port map( D => n1776, CP => clk, 
                           RN => n2768, Q => registers_11_22_port);
   registers_reg_11_21_inst : HS65_LH_DFPRQX9 port map( D => n1775, CP => clk, 
                           RN => n2768, Q => registers_11_21_port);
   registers_reg_11_20_inst : HS65_LH_DFPRQX9 port map( D => n1774, CP => clk, 
                           RN => n2768, Q => registers_11_20_port);
   registers_reg_11_19_inst : HS65_LH_DFPRQX9 port map( D => n1773, CP => clk, 
                           RN => n2769, Q => registers_11_19_port);
   registers_reg_11_18_inst : HS65_LH_DFPRQX9 port map( D => n1772, CP => clk, 
                           RN => n2769, Q => registers_11_18_port);
   registers_reg_11_17_inst : HS65_LH_DFPRQX9 port map( D => n1771, CP => clk, 
                           RN => n2769, Q => registers_11_17_port);
   registers_reg_11_16_inst : HS65_LH_DFPRQX9 port map( D => n1770, CP => clk, 
                           RN => n2769, Q => registers_11_16_port);
   registers_reg_11_15_inst : HS65_LH_DFPRQX9 port map( D => n1769, CP => clk, 
                           RN => n2769, Q => registers_11_15_port);
   registers_reg_11_14_inst : HS65_LH_DFPRQX9 port map( D => n1768, CP => clk, 
                           RN => n2769, Q => registers_11_14_port);
   registers_reg_11_13_inst : HS65_LH_DFPRQX9 port map( D => n1767, CP => clk, 
                           RN => n2769, Q => registers_11_13_port);
   registers_reg_11_12_inst : HS65_LH_DFPRQX9 port map( D => n1766, CP => clk, 
                           RN => n2769, Q => registers_11_12_port);
   registers_reg_11_11_inst : HS65_LH_DFPRQX9 port map( D => n1765, CP => clk, 
                           RN => n2769, Q => registers_11_11_port);
   registers_reg_11_10_inst : HS65_LH_DFPRQX9 port map( D => n1764, CP => clk, 
                           RN => n2769, Q => registers_11_10_port);
   registers_reg_11_9_inst : HS65_LH_DFPRQX9 port map( D => n1763, CP => clk, 
                           RN => n2769, Q => registers_11_9_port);
   registers_reg_11_8_inst : HS65_LH_DFPRQX9 port map( D => n1762, CP => clk, 
                           RN => n2770, Q => registers_11_8_port);
   registers_reg_11_7_inst : HS65_LH_DFPRQX9 port map( D => n1761, CP => clk, 
                           RN => n2770, Q => registers_11_7_port);
   registers_reg_11_6_inst : HS65_LH_DFPRQX9 port map( D => n1760, CP => clk, 
                           RN => n2770, Q => registers_11_6_port);
   registers_reg_11_5_inst : HS65_LH_DFPRQX9 port map( D => n1759, CP => clk, 
                           RN => n2770, Q => registers_11_5_port);
   registers_reg_11_4_inst : HS65_LH_DFPRQX9 port map( D => n1758, CP => clk, 
                           RN => n2770, Q => registers_11_4_port);
   registers_reg_11_3_inst : HS65_LH_DFPRQX9 port map( D => n1757, CP => clk, 
                           RN => n2770, Q => registers_11_3_port);
   registers_reg_11_2_inst : HS65_LH_DFPRQX9 port map( D => n1756, CP => clk, 
                           RN => n2770, Q => registers_11_2_port);
   registers_reg_11_1_inst : HS65_LH_DFPRQX9 port map( D => n1755, CP => clk, 
                           RN => n2770, Q => registers_11_1_port);
   registers_reg_11_0_inst : HS65_LH_DFPRQX9 port map( D => n1754, CP => clk, 
                           RN => n2770, Q => registers_11_0_port);
   registers_reg_10_31_inst : HS65_LH_DFPRQX9 port map( D => n1753, CP => clk, 
                           RN => n2770, Q => registers_10_31_port);
   registers_reg_10_30_inst : HS65_LH_DFPRQX9 port map( D => n1752, CP => clk, 
                           RN => n2770, Q => registers_10_30_port);
   registers_reg_10_29_inst : HS65_LH_DFPRQX9 port map( D => n1751, CP => clk, 
                           RN => n2770, Q => registers_10_29_port);
   registers_reg_10_28_inst : HS65_LH_DFPRQX9 port map( D => n1750, CP => clk, 
                           RN => n2771, Q => registers_10_28_port);
   registers_reg_10_27_inst : HS65_LH_DFPRQX9 port map( D => n1749, CP => clk, 
                           RN => n2771, Q => registers_10_27_port);
   registers_reg_10_26_inst : HS65_LH_DFPRQX9 port map( D => n1748, CP => clk, 
                           RN => n2771, Q => registers_10_26_port);
   registers_reg_10_25_inst : HS65_LH_DFPRQX9 port map( D => n1747, CP => clk, 
                           RN => n2771, Q => registers_10_25_port);
   registers_reg_10_24_inst : HS65_LH_DFPRQX9 port map( D => n1746, CP => clk, 
                           RN => n2771, Q => registers_10_24_port);
   registers_reg_10_23_inst : HS65_LH_DFPRQX9 port map( D => n1745, CP => clk, 
                           RN => n2771, Q => registers_10_23_port);
   registers_reg_10_22_inst : HS65_LH_DFPRQX9 port map( D => n1744, CP => clk, 
                           RN => n2771, Q => registers_10_22_port);
   registers_reg_10_21_inst : HS65_LH_DFPRQX9 port map( D => n1743, CP => clk, 
                           RN => n2771, Q => registers_10_21_port);
   registers_reg_10_20_inst : HS65_LH_DFPRQX9 port map( D => n1742, CP => clk, 
                           RN => n2771, Q => registers_10_20_port);
   registers_reg_10_19_inst : HS65_LH_DFPRQX9 port map( D => n1741, CP => clk, 
                           RN => n2771, Q => registers_10_19_port);
   registers_reg_10_18_inst : HS65_LH_DFPRQX9 port map( D => n1740, CP => clk, 
                           RN => n2771, Q => registers_10_18_port);
   registers_reg_10_17_inst : HS65_LH_DFPRQX9 port map( D => n1739, CP => clk, 
                           RN => n2771, Q => registers_10_17_port);
   registers_reg_10_16_inst : HS65_LH_DFPRQX9 port map( D => n1738, CP => clk, 
                           RN => n2772, Q => registers_10_16_port);
   registers_reg_10_15_inst : HS65_LH_DFPRQX9 port map( D => n1737, CP => clk, 
                           RN => n2772, Q => registers_10_15_port);
   registers_reg_10_14_inst : HS65_LH_DFPRQX9 port map( D => n1736, CP => clk, 
                           RN => n2772, Q => registers_10_14_port);
   registers_reg_10_13_inst : HS65_LH_DFPRQX9 port map( D => n1735, CP => clk, 
                           RN => n2772, Q => registers_10_13_port);
   registers_reg_10_12_inst : HS65_LH_DFPRQX9 port map( D => n1734, CP => clk, 
                           RN => n2772, Q => registers_10_12_port);
   registers_reg_10_11_inst : HS65_LH_DFPRQX9 port map( D => n1733, CP => clk, 
                           RN => n2772, Q => registers_10_11_port);
   registers_reg_10_10_inst : HS65_LH_DFPRQX9 port map( D => n1732, CP => clk, 
                           RN => n2772, Q => registers_10_10_port);
   registers_reg_10_9_inst : HS65_LH_DFPRQX9 port map( D => n1731, CP => clk, 
                           RN => n2772, Q => registers_10_9_port);
   registers_reg_10_8_inst : HS65_LH_DFPRQX9 port map( D => n1730, CP => clk, 
                           RN => n2772, Q => registers_10_8_port);
   registers_reg_10_7_inst : HS65_LH_DFPRQX9 port map( D => n1729, CP => clk, 
                           RN => n2772, Q => registers_10_7_port);
   registers_reg_10_6_inst : HS65_LH_DFPRQX9 port map( D => n1728, CP => clk, 
                           RN => n2772, Q => registers_10_6_port);
   registers_reg_10_5_inst : HS65_LH_DFPRQX9 port map( D => n1727, CP => clk, 
                           RN => n2772, Q => registers_10_5_port);
   registers_reg_10_4_inst : HS65_LH_DFPRQX9 port map( D => n1726, CP => clk, 
                           RN => n2773, Q => registers_10_4_port);
   registers_reg_10_3_inst : HS65_LH_DFPRQX9 port map( D => n1725, CP => clk, 
                           RN => n2773, Q => registers_10_3_port);
   registers_reg_10_2_inst : HS65_LH_DFPRQX9 port map( D => n1724, CP => clk, 
                           RN => n2773, Q => registers_10_2_port);
   registers_reg_10_1_inst : HS65_LH_DFPRQX9 port map( D => n1723, CP => clk, 
                           RN => n2773, Q => registers_10_1_port);
   registers_reg_10_0_inst : HS65_LH_DFPRQX9 port map( D => n1722, CP => clk, 
                           RN => n2773, Q => registers_10_0_port);
   registers_reg_7_31_inst : HS65_LH_DFPRQX9 port map( D => n1657, CP => clk, 
                           RN => n2773, Q => registers_7_31_port);
   registers_reg_7_30_inst : HS65_LH_DFPRQX9 port map( D => n1656, CP => clk, 
                           RN => n2773, Q => registers_7_30_port);
   registers_reg_7_29_inst : HS65_LH_DFPRQX9 port map( D => n1655, CP => clk, 
                           RN => n2773, Q => registers_7_29_port);
   registers_reg_7_28_inst : HS65_LH_DFPRQX9 port map( D => n1654, CP => clk, 
                           RN => n2773, Q => registers_7_28_port);
   registers_reg_7_27_inst : HS65_LH_DFPRQX9 port map( D => n1653, CP => clk, 
                           RN => n2773, Q => registers_7_27_port);
   registers_reg_7_26_inst : HS65_LH_DFPRQX9 port map( D => n1652, CP => clk, 
                           RN => n2773, Q => registers_7_26_port);
   registers_reg_7_25_inst : HS65_LH_DFPRQX9 port map( D => n1651, CP => clk, 
                           RN => n2773, Q => registers_7_25_port);
   registers_reg_7_24_inst : HS65_LH_DFPRQX9 port map( D => n1650, CP => clk, 
                           RN => n2774, Q => registers_7_24_port);
   registers_reg_7_23_inst : HS65_LH_DFPRQX9 port map( D => n1649, CP => clk, 
                           RN => n2796, Q => registers_7_23_port);
   registers_reg_7_22_inst : HS65_LH_DFPRQX9 port map( D => n1648, CP => clk, 
                           RN => n2792, Q => registers_7_22_port);
   registers_reg_7_21_inst : HS65_LH_DFPRQX9 port map( D => n1647, CP => clk, 
                           RN => n2792, Q => registers_7_21_port);
   registers_reg_7_20_inst : HS65_LH_DFPRQX9 port map( D => n1646, CP => clk, 
                           RN => n2792, Q => registers_7_20_port);
   registers_reg_7_19_inst : HS65_LH_DFPRQX9 port map( D => n1645, CP => clk, 
                           RN => n2792, Q => registers_7_19_port);
   registers_reg_7_18_inst : HS65_LH_DFPRQX9 port map( D => n1644, CP => clk, 
                           RN => n2792, Q => registers_7_18_port);
   registers_reg_7_17_inst : HS65_LH_DFPRQX9 port map( D => n1643, CP => clk, 
                           RN => n2792, Q => registers_7_17_port);
   registers_reg_7_16_inst : HS65_LH_DFPRQX9 port map( D => n1642, CP => clk, 
                           RN => n2792, Q => registers_7_16_port);
   registers_reg_7_15_inst : HS65_LH_DFPRQX9 port map( D => n1641, CP => clk, 
                           RN => n2792, Q => registers_7_15_port);
   registers_reg_7_14_inst : HS65_LH_DFPRQX9 port map( D => n1640, CP => clk, 
                           RN => n2792, Q => registers_7_14_port);
   registers_reg_7_13_inst : HS65_LH_DFPRQX9 port map( D => n1639, CP => clk, 
                           RN => n2792, Q => registers_7_13_port);
   registers_reg_7_12_inst : HS65_LH_DFPRQX9 port map( D => n1638, CP => clk, 
                           RN => n2792, Q => registers_7_12_port);
   registers_reg_7_11_inst : HS65_LH_DFPRQX9 port map( D => n1637, CP => clk, 
                           RN => n2793, Q => registers_7_11_port);
   registers_reg_7_10_inst : HS65_LH_DFPRQX9 port map( D => n1636, CP => clk, 
                           RN => n2793, Q => registers_7_10_port);
   registers_reg_7_9_inst : HS65_LH_DFPRQX9 port map( D => n1635, CP => clk, RN
                           => n2793, Q => registers_7_9_port);
   registers_reg_7_8_inst : HS65_LH_DFPRQX9 port map( D => n1634, CP => clk, RN
                           => n2793, Q => registers_7_8_port);
   registers_reg_7_7_inst : HS65_LH_DFPRQX9 port map( D => n1633, CP => clk, RN
                           => n2793, Q => registers_7_7_port);
   registers_reg_7_6_inst : HS65_LH_DFPRQX9 port map( D => n1632, CP => clk, RN
                           => n2793, Q => registers_7_6_port);
   registers_reg_7_5_inst : HS65_LH_DFPRQX9 port map( D => n1631, CP => clk, RN
                           => n2793, Q => registers_7_5_port);
   registers_reg_7_4_inst : HS65_LH_DFPRQX9 port map( D => n1630, CP => clk, RN
                           => n2793, Q => registers_7_4_port);
   registers_reg_7_3_inst : HS65_LH_DFPRQX9 port map( D => n1629, CP => clk, RN
                           => n2793, Q => registers_7_3_port);
   registers_reg_7_2_inst : HS65_LH_DFPRQX9 port map( D => n1628, CP => clk, RN
                           => n2793, Q => registers_7_2_port);
   registers_reg_7_1_inst : HS65_LH_DFPRQX9 port map( D => n1627, CP => clk, RN
                           => n2793, Q => registers_7_1_port);
   registers_reg_7_0_inst : HS65_LH_DFPRQX9 port map( D => n1626, CP => clk, RN
                           => n2793, Q => registers_7_0_port);
   registers_reg_6_31_inst : HS65_LH_DFPRQX9 port map( D => n1625, CP => clk, 
                           RN => n2794, Q => registers_6_31_port);
   registers_reg_6_30_inst : HS65_LH_DFPRQX9 port map( D => n1624, CP => clk, 
                           RN => n2794, Q => registers_6_30_port);
   registers_reg_6_29_inst : HS65_LH_DFPRQX9 port map( D => n1623, CP => clk, 
                           RN => n2794, Q => registers_6_29_port);
   registers_reg_6_28_inst : HS65_LH_DFPRQX9 port map( D => n1622, CP => clk, 
                           RN => n2794, Q => registers_6_28_port);
   registers_reg_6_27_inst : HS65_LH_DFPRQX9 port map( D => n1621, CP => clk, 
                           RN => n2794, Q => registers_6_27_port);
   registers_reg_6_26_inst : HS65_LH_DFPRQX9 port map( D => n1620, CP => clk, 
                           RN => n2794, Q => registers_6_26_port);
   registers_reg_6_25_inst : HS65_LH_DFPRQX9 port map( D => n1619, CP => clk, 
                           RN => n2794, Q => registers_6_25_port);
   registers_reg_6_24_inst : HS65_LH_DFPRQX9 port map( D => n1618, CP => clk, 
                           RN => n2794, Q => registers_6_24_port);
   registers_reg_6_23_inst : HS65_LH_DFPRQX9 port map( D => n1617, CP => clk, 
                           RN => n2794, Q => registers_6_23_port);
   registers_reg_6_22_inst : HS65_LH_DFPRQX9 port map( D => n1616, CP => clk, 
                           RN => n2794, Q => registers_6_22_port);
   registers_reg_6_21_inst : HS65_LH_DFPRQX9 port map( D => n1615, CP => clk, 
                           RN => n2794, Q => registers_6_21_port);
   registers_reg_6_20_inst : HS65_LH_DFPRQX9 port map( D => n1614, CP => clk, 
                           RN => n2794, Q => registers_6_20_port);
   registers_reg_6_19_inst : HS65_LH_DFPRQX9 port map( D => n1613, CP => clk, 
                           RN => n2795, Q => registers_6_19_port);
   registers_reg_6_18_inst : HS65_LH_DFPRQX9 port map( D => n1612, CP => clk, 
                           RN => n2795, Q => registers_6_18_port);
   registers_reg_6_17_inst : HS65_LH_DFPRQX9 port map( D => n1611, CP => clk, 
                           RN => n2795, Q => registers_6_17_port);
   registers_reg_6_16_inst : HS65_LH_DFPRQX9 port map( D => n1610, CP => clk, 
                           RN => n2795, Q => registers_6_16_port);
   registers_reg_6_15_inst : HS65_LH_DFPRQX9 port map( D => n1609, CP => clk, 
                           RN => n2795, Q => registers_6_15_port);
   registers_reg_6_14_inst : HS65_LH_DFPRQX9 port map( D => n1608, CP => clk, 
                           RN => n2795, Q => registers_6_14_port);
   registers_reg_6_13_inst : HS65_LH_DFPRQX9 port map( D => n1607, CP => clk, 
                           RN => n2795, Q => registers_6_13_port);
   registers_reg_6_12_inst : HS65_LH_DFPRQX9 port map( D => n1606, CP => clk, 
                           RN => n2795, Q => registers_6_12_port);
   registers_reg_6_11_inst : HS65_LH_DFPRQX9 port map( D => n1605, CP => clk, 
                           RN => n2795, Q => registers_6_11_port);
   registers_reg_6_10_inst : HS65_LH_DFPRQX9 port map( D => n1604, CP => clk, 
                           RN => n2795, Q => registers_6_10_port);
   registers_reg_6_9_inst : HS65_LH_DFPRQX9 port map( D => n1603, CP => clk, RN
                           => n2795, Q => registers_6_9_port);
   registers_reg_6_8_inst : HS65_LH_DFPRQX9 port map( D => n1602, CP => clk, RN
                           => n2795, Q => registers_6_8_port);
   registers_reg_6_7_inst : HS65_LH_DFPRQX9 port map( D => n1601, CP => clk, RN
                           => n2796, Q => registers_6_7_port);
   registers_reg_6_6_inst : HS65_LH_DFPRQX9 port map( D => n1600, CP => clk, RN
                           => n2796, Q => registers_6_6_port);
   registers_reg_6_5_inst : HS65_LH_DFPRQX9 port map( D => n1599, CP => clk, RN
                           => n2796, Q => registers_6_5_port);
   registers_reg_6_4_inst : HS65_LH_DFPRQX9 port map( D => n1598, CP => clk, RN
                           => n2796, Q => registers_6_4_port);
   registers_reg_6_3_inst : HS65_LH_DFPRQX9 port map( D => n1597, CP => clk, RN
                           => n2796, Q => registers_6_3_port);
   registers_reg_6_2_inst : HS65_LH_DFPRQX9 port map( D => n1596, CP => clk, RN
                           => n2796, Q => registers_6_2_port);
   registers_reg_6_1_inst : HS65_LH_DFPRQX9 port map( D => n1595, CP => clk, RN
                           => n2796, Q => registers_6_1_port);
   registers_reg_6_0_inst : HS65_LH_DFPRQX9 port map( D => n1594, CP => clk, RN
                           => n2796, Q => registers_6_0_port);
   registers_reg_5_31_inst : HS65_LH_DFPRQX9 port map( D => n1593, CP => clk, 
                           RN => n2796, Q => registers_5_31_port);
   registers_reg_5_30_inst : HS65_LH_DFPRQX9 port map( D => n1592, CP => clk, 
                           RN => n2796, Q => registers_5_30_port);
   registers_reg_5_29_inst : HS65_LH_DFPRQX9 port map( D => n1591, CP => clk, 
                           RN => n2796, Q => registers_5_29_port);
   registers_reg_5_28_inst : HS65_LH_DFPRQX9 port map( D => n1590, CP => clk, 
                           RN => n2797, Q => registers_5_28_port);
   registers_reg_5_27_inst : HS65_LH_DFPRQX9 port map( D => n1589, CP => clk, 
                           RN => n2797, Q => registers_5_27_port);
   registers_reg_5_26_inst : HS65_LH_DFPRQX9 port map( D => n1588, CP => clk, 
                           RN => n2797, Q => registers_5_26_port);
   registers_reg_5_25_inst : HS65_LH_DFPRQX9 port map( D => n1587, CP => clk, 
                           RN => n2797, Q => registers_5_25_port);
   registers_reg_5_24_inst : HS65_LH_DFPRQX9 port map( D => n1586, CP => clk, 
                           RN => n2797, Q => registers_5_24_port);
   registers_reg_5_23_inst : HS65_LH_DFPRQX9 port map( D => n1585, CP => clk, 
                           RN => n2797, Q => registers_5_23_port);
   registers_reg_5_22_inst : HS65_LH_DFPRQX9 port map( D => n1584, CP => clk, 
                           RN => n2797, Q => registers_5_22_port);
   registers_reg_5_21_inst : HS65_LH_DFPRQX9 port map( D => n1583, CP => clk, 
                           RN => n2797, Q => registers_5_21_port);
   registers_reg_5_20_inst : HS65_LH_DFPRQX9 port map( D => n1582, CP => clk, 
                           RN => n2797, Q => registers_5_20_port);
   registers_reg_5_19_inst : HS65_LH_DFPRQX9 port map( D => n1581, CP => clk, 
                           RN => n2797, Q => registers_5_19_port);
   registers_reg_5_18_inst : HS65_LH_DFPRQX9 port map( D => n1580, CP => clk, 
                           RN => n2797, Q => registers_5_18_port);
   registers_reg_5_17_inst : HS65_LH_DFPRQX9 port map( D => n1579, CP => clk, 
                           RN => n2797, Q => registers_5_17_port);
   registers_reg_5_16_inst : HS65_LH_DFPRQX9 port map( D => n1578, CP => clk, 
                           RN => n2798, Q => registers_5_16_port);
   registers_reg_5_15_inst : HS65_LH_DFPRQX9 port map( D => n1577, CP => clk, 
                           RN => n2798, Q => registers_5_15_port);
   registers_reg_5_14_inst : HS65_LH_DFPRQX9 port map( D => n1576, CP => clk, 
                           RN => n2798, Q => registers_5_14_port);
   registers_reg_5_13_inst : HS65_LH_DFPRQX9 port map( D => n1575, CP => clk, 
                           RN => n2798, Q => registers_5_13_port);
   registers_reg_5_12_inst : HS65_LH_DFPRQX9 port map( D => n1574, CP => clk, 
                           RN => n2798, Q => registers_5_12_port);
   registers_reg_5_11_inst : HS65_LH_DFPRQX9 port map( D => n1573, CP => clk, 
                           RN => n2798, Q => registers_5_11_port);
   registers_reg_5_10_inst : HS65_LH_DFPRQX9 port map( D => n1572, CP => clk, 
                           RN => n2798, Q => registers_5_10_port);
   registers_reg_5_9_inst : HS65_LH_DFPRQX9 port map( D => n1571, CP => clk, RN
                           => n2798, Q => registers_5_9_port);
   registers_reg_5_8_inst : HS65_LH_DFPRQX9 port map( D => n1570, CP => clk, RN
                           => n2798, Q => registers_5_8_port);
   registers_reg_5_7_inst : HS65_LH_DFPRQX9 port map( D => n1569, CP => clk, RN
                           => n2798, Q => registers_5_7_port);
   registers_reg_5_6_inst : HS65_LH_DFPRQX9 port map( D => n1568, CP => clk, RN
                           => n2798, Q => registers_5_6_port);
   registers_reg_5_5_inst : HS65_LH_DFPRQX9 port map( D => n1567, CP => clk, RN
                           => n2798, Q => registers_5_5_port);
   registers_reg_5_4_inst : HS65_LH_DFPRQX9 port map( D => n1566, CP => clk, RN
                           => n2799, Q => registers_5_4_port);
   registers_reg_5_3_inst : HS65_LH_DFPRQX9 port map( D => n1565, CP => clk, RN
                           => n2799, Q => registers_5_3_port);
   registers_reg_5_2_inst : HS65_LH_DFPRQX9 port map( D => n1564, CP => clk, RN
                           => n2799, Q => registers_5_2_port);
   registers_reg_5_1_inst : HS65_LH_DFPRQX9 port map( D => n1563, CP => clk, RN
                           => n2799, Q => registers_5_1_port);
   registers_reg_5_0_inst : HS65_LH_DFPRQX9 port map( D => n1562, CP => clk, RN
                           => n2799, Q => registers_5_0_port);
   registers_reg_4_31_inst : HS65_LH_DFPRQX9 port map( D => n1561, CP => clk, 
                           RN => n2799, Q => registers_4_31_port);
   registers_reg_4_30_inst : HS65_LH_DFPRQX9 port map( D => n1560, CP => clk, 
                           RN => n2799, Q => registers_4_30_port);
   registers_reg_4_29_inst : HS65_LH_DFPRQX9 port map( D => n1559, CP => clk, 
                           RN => n2799, Q => registers_4_29_port);
   registers_reg_4_28_inst : HS65_LH_DFPRQX9 port map( D => n1558, CP => clk, 
                           RN => n2801, Q => registers_4_28_port);
   registers_reg_4_27_inst : HS65_LH_DFPRQX9 port map( D => n1557, CP => clk, 
                           RN => n2799, Q => registers_4_27_port);
   registers_reg_4_26_inst : HS65_LH_DFPRQX9 port map( D => n1556, CP => clk, 
                           RN => n2799, Q => registers_4_26_port);
   registers_reg_4_25_inst : HS65_LH_DFPRQX9 port map( D => n1555, CP => clk, 
                           RN => n2799, Q => registers_4_25_port);
   registers_reg_4_24_inst : HS65_LH_DFPRQX9 port map( D => n1554, CP => clk, 
                           RN => n2800, Q => registers_4_24_port);
   registers_reg_4_23_inst : HS65_LH_DFPRQX9 port map( D => n1553, CP => clk, 
                           RN => n2800, Q => registers_4_23_port);
   registers_reg_4_22_inst : HS65_LH_DFPRQX9 port map( D => n1552, CP => clk, 
                           RN => n2800, Q => registers_4_22_port);
   registers_reg_4_21_inst : HS65_LH_DFPRQX9 port map( D => n1551, CP => clk, 
                           RN => n2800, Q => registers_4_21_port);
   registers_reg_4_20_inst : HS65_LH_DFPRQX9 port map( D => n1550, CP => clk, 
                           RN => n2800, Q => registers_4_20_port);
   registers_reg_4_19_inst : HS65_LH_DFPRQX9 port map( D => n1549, CP => clk, 
                           RN => n2800, Q => registers_4_19_port);
   registers_reg_4_18_inst : HS65_LH_DFPRQX9 port map( D => n1548, CP => clk, 
                           RN => n2800, Q => registers_4_18_port);
   registers_reg_4_17_inst : HS65_LH_DFPRQX9 port map( D => n1547, CP => clk, 
                           RN => n2800, Q => registers_4_17_port);
   registers_reg_4_16_inst : HS65_LH_DFPRQX9 port map( D => n1546, CP => clk, 
                           RN => n2800, Q => registers_4_16_port);
   registers_reg_4_15_inst : HS65_LH_DFPRQX9 port map( D => n1545, CP => clk, 
                           RN => n2800, Q => registers_4_15_port);
   registers_reg_4_14_inst : HS65_LH_DFPRQX9 port map( D => n1544, CP => clk, 
                           RN => n2800, Q => registers_4_14_port);
   registers_reg_4_13_inst : HS65_LH_DFPRQX9 port map( D => n1543, CP => clk, 
                           RN => n2800, Q => registers_4_13_port);
   registers_reg_4_12_inst : HS65_LH_DFPRQX9 port map( D => n1542, CP => clk, 
                           RN => n2787, Q => registers_4_12_port);
   registers_reg_4_11_inst : HS65_LH_DFPRQX9 port map( D => n1541, CP => clk, 
                           RN => n2783, Q => registers_4_11_port);
   registers_reg_4_10_inst : HS65_LH_DFPRQX9 port map( D => n1540, CP => clk, 
                           RN => n2783, Q => registers_4_10_port);
   registers_reg_4_9_inst : HS65_LH_DFPRQX9 port map( D => n1539, CP => clk, RN
                           => n2783, Q => registers_4_9_port);
   registers_reg_4_8_inst : HS65_LH_DFPRQX9 port map( D => n1538, CP => clk, RN
                           => n2783, Q => registers_4_8_port);
   registers_reg_4_7_inst : HS65_LH_DFPRQX9 port map( D => n1537, CP => clk, RN
                           => n2783, Q => registers_4_7_port);
   registers_reg_4_6_inst : HS65_LH_DFPRQX9 port map( D => n1536, CP => clk, RN
                           => n2783, Q => registers_4_6_port);
   registers_reg_4_5_inst : HS65_LH_DFPRQX9 port map( D => n1535, CP => clk, RN
                           => n2783, Q => registers_4_5_port);
   registers_reg_4_4_inst : HS65_LH_DFPRQX9 port map( D => n1534, CP => clk, RN
                           => n2783, Q => registers_4_4_port);
   registers_reg_4_3_inst : HS65_LH_DFPRQX9 port map( D => n1533, CP => clk, RN
                           => n2783, Q => registers_4_3_port);
   registers_reg_4_2_inst : HS65_LH_DFPRQX9 port map( D => n1532, CP => clk, RN
                           => n2783, Q => registers_4_2_port);
   registers_reg_4_1_inst : HS65_LH_DFPRQX9 port map( D => n1531, CP => clk, RN
                           => n2783, Q => registers_4_1_port);
   registers_reg_4_0_inst : HS65_LH_DFPRQX9 port map( D => n1530, CP => clk, RN
                           => n2784, Q => registers_4_0_port);
   registers_reg_3_31_inst : HS65_LH_DFPRQX9 port map( D => n1529, CP => clk, 
                           RN => n2784, Q => registers_3_31_port);
   registers_reg_3_30_inst : HS65_LH_DFPRQX9 port map( D => n1528, CP => clk, 
                           RN => n2784, Q => registers_3_30_port);
   registers_reg_3_29_inst : HS65_LH_DFPRQX9 port map( D => n1527, CP => clk, 
                           RN => n2784, Q => registers_3_29_port);
   registers_reg_3_28_inst : HS65_LH_DFPRQX9 port map( D => n1526, CP => clk, 
                           RN => n2784, Q => registers_3_28_port);
   registers_reg_3_27_inst : HS65_LH_DFPRQX9 port map( D => n1525, CP => clk, 
                           RN => n2784, Q => registers_3_27_port);
   registers_reg_3_26_inst : HS65_LH_DFPRQX9 port map( D => n1524, CP => clk, 
                           RN => n2784, Q => registers_3_26_port);
   registers_reg_3_25_inst : HS65_LH_DFPRQX9 port map( D => n1523, CP => clk, 
                           RN => n2784, Q => registers_3_25_port);
   registers_reg_3_24_inst : HS65_LH_DFPRQX9 port map( D => n1522, CP => clk, 
                           RN => n2784, Q => registers_3_24_port);
   registers_reg_3_23_inst : HS65_LH_DFPRQX9 port map( D => n1521, CP => clk, 
                           RN => n2784, Q => registers_3_23_port);
   registers_reg_3_22_inst : HS65_LH_DFPRQX9 port map( D => n1520, CP => clk, 
                           RN => n2784, Q => registers_3_22_port);
   registers_reg_3_21_inst : HS65_LH_DFPRQX9 port map( D => n1519, CP => clk, 
                           RN => n2784, Q => registers_3_21_port);
   registers_reg_3_20_inst : HS65_LH_DFPRQX9 port map( D => n1518, CP => clk, 
                           RN => n2785, Q => registers_3_20_port);
   registers_reg_3_19_inst : HS65_LH_DFPRQX9 port map( D => n1517, CP => clk, 
                           RN => n2785, Q => registers_3_19_port);
   registers_reg_3_18_inst : HS65_LH_DFPRQX9 port map( D => n1516, CP => clk, 
                           RN => n2785, Q => registers_3_18_port);
   registers_reg_3_17_inst : HS65_LH_DFPRQX9 port map( D => n1515, CP => clk, 
                           RN => n2785, Q => registers_3_17_port);
   registers_reg_3_16_inst : HS65_LH_DFPRQX9 port map( D => n1514, CP => clk, 
                           RN => n2785, Q => registers_3_16_port);
   registers_reg_3_15_inst : HS65_LH_DFPRQX9 port map( D => n1513, CP => clk, 
                           RN => n2785, Q => registers_3_15_port);
   registers_reg_3_14_inst : HS65_LH_DFPRQX9 port map( D => n1512, CP => clk, 
                           RN => n2785, Q => registers_3_14_port);
   registers_reg_3_13_inst : HS65_LH_DFPRQX9 port map( D => n1511, CP => clk, 
                           RN => n2785, Q => registers_3_13_port);
   registers_reg_3_12_inst : HS65_LH_DFPRQX9 port map( D => n1510, CP => clk, 
                           RN => n2785, Q => registers_3_12_port);
   registers_reg_3_11_inst : HS65_LH_DFPRQX9 port map( D => n1509, CP => clk, 
                           RN => n2785, Q => registers_3_11_port);
   registers_reg_3_10_inst : HS65_LH_DFPRQX9 port map( D => n1508, CP => clk, 
                           RN => n2785, Q => registers_3_10_port);
   registers_reg_3_9_inst : HS65_LH_DFPRQX9 port map( D => n1507, CP => clk, RN
                           => n2785, Q => registers_3_9_port);
   registers_reg_3_8_inst : HS65_LH_DFPRQX9 port map( D => n1506, CP => clk, RN
                           => n2786, Q => registers_3_8_port);
   registers_reg_3_7_inst : HS65_LH_DFPRQX9 port map( D => n1505, CP => clk, RN
                           => n2786, Q => registers_3_7_port);
   registers_reg_3_6_inst : HS65_LH_DFPRQX9 port map( D => n1504, CP => clk, RN
                           => n2786, Q => registers_3_6_port);
   registers_reg_3_5_inst : HS65_LH_DFPRQX9 port map( D => n1503, CP => clk, RN
                           => n2786, Q => registers_3_5_port);
   registers_reg_3_4_inst : HS65_LH_DFPRQX9 port map( D => n1502, CP => clk, RN
                           => n2786, Q => registers_3_4_port);
   registers_reg_3_3_inst : HS65_LH_DFPRQX9 port map( D => n1501, CP => clk, RN
                           => n2786, Q => registers_3_3_port);
   registers_reg_3_2_inst : HS65_LH_DFPRQX9 port map( D => n1500, CP => clk, RN
                           => n2786, Q => registers_3_2_port);
   registers_reg_3_1_inst : HS65_LH_DFPRQX9 port map( D => n1499, CP => clk, RN
                           => n2786, Q => registers_3_1_port);
   registers_reg_3_0_inst : HS65_LH_DFPRQX9 port map( D => n1498, CP => clk, RN
                           => n2786, Q => registers_3_0_port);
   registers_reg_2_31_inst : HS65_LH_DFPRQX9 port map( D => n1497, CP => clk, 
                           RN => n2786, Q => registers_2_31_port);
   registers_reg_2_30_inst : HS65_LH_DFPRQX9 port map( D => n1496, CP => clk, 
                           RN => n2786, Q => registers_2_30_port);
   registers_reg_2_29_inst : HS65_LH_DFPRQX9 port map( D => n1495, CP => clk, 
                           RN => n2786, Q => registers_2_29_port);
   registers_reg_2_28_inst : HS65_LH_DFPRQX9 port map( D => n1494, CP => clk, 
                           RN => n2787, Q => registers_2_28_port);
   registers_reg_2_27_inst : HS65_LH_DFPRQX9 port map( D => n1493, CP => clk, 
                           RN => n2787, Q => registers_2_27_port);
   registers_reg_2_26_inst : HS65_LH_DFPRQX9 port map( D => n1492, CP => clk, 
                           RN => n2787, Q => registers_2_26_port);
   registers_reg_2_25_inst : HS65_LH_DFPRQX9 port map( D => n1491, CP => clk, 
                           RN => n2787, Q => registers_2_25_port);
   registers_reg_2_24_inst : HS65_LH_DFPRQX9 port map( D => n1490, CP => clk, 
                           RN => n2787, Q => registers_2_24_port);
   registers_reg_2_23_inst : HS65_LH_DFPRQX9 port map( D => n1489, CP => clk, 
                           RN => n2787, Q => registers_2_23_port);
   registers_reg_2_22_inst : HS65_LH_DFPRQX9 port map( D => n1488, CP => clk, 
                           RN => n2787, Q => registers_2_22_port);
   registers_reg_2_21_inst : HS65_LH_DFPRQX9 port map( D => n1487, CP => clk, 
                           RN => n2787, Q => registers_2_21_port);
   registers_reg_2_20_inst : HS65_LH_DFPRQX9 port map( D => n1486, CP => clk, 
                           RN => n2787, Q => registers_2_20_port);
   registers_reg_2_19_inst : HS65_LH_DFPRQX9 port map( D => n1485, CP => clk, 
                           RN => n2787, Q => registers_2_19_port);
   registers_reg_2_18_inst : HS65_LH_DFPRQX9 port map( D => n1484, CP => clk, 
                           RN => n2787, Q => registers_2_18_port);
   registers_reg_2_17_inst : HS65_LH_DFPRQX9 port map( D => n1483, CP => clk, 
                           RN => n2788, Q => registers_2_17_port);
   registers_reg_2_16_inst : HS65_LH_DFPRQX9 port map( D => n1482, CP => clk, 
                           RN => n2788, Q => registers_2_16_port);
   registers_reg_2_15_inst : HS65_LH_DFPRQX9 port map( D => n1481, CP => clk, 
                           RN => n2788, Q => registers_2_15_port);
   registers_reg_2_14_inst : HS65_LH_DFPRQX9 port map( D => n1480, CP => clk, 
                           RN => n2788, Q => registers_2_14_port);
   registers_reg_2_13_inst : HS65_LH_DFPRQX9 port map( D => n1479, CP => clk, 
                           RN => n2788, Q => registers_2_13_port);
   registers_reg_2_12_inst : HS65_LH_DFPRQX9 port map( D => n1478, CP => clk, 
                           RN => n2788, Q => registers_2_12_port);
   registers_reg_2_11_inst : HS65_LH_DFPRQX9 port map( D => n1477, CP => clk, 
                           RN => n2788, Q => registers_2_11_port);
   registers_reg_2_10_inst : HS65_LH_DFPRQX9 port map( D => n1476, CP => clk, 
                           RN => n2788, Q => registers_2_10_port);
   registers_reg_2_9_inst : HS65_LH_DFPRQX9 port map( D => n1475, CP => clk, RN
                           => n2788, Q => registers_2_9_port);
   registers_reg_2_8_inst : HS65_LH_DFPRQX9 port map( D => n1474, CP => clk, RN
                           => n2788, Q => registers_2_8_port);
   registers_reg_2_7_inst : HS65_LH_DFPRQX9 port map( D => n1473, CP => clk, RN
                           => n2788, Q => registers_2_7_port);
   registers_reg_2_6_inst : HS65_LH_DFPRQX9 port map( D => n1472, CP => clk, RN
                           => n2788, Q => registers_2_6_port);
   registers_reg_2_5_inst : HS65_LH_DFPRQX9 port map( D => n1471, CP => clk, RN
                           => n2789, Q => registers_2_5_port);
   registers_reg_2_4_inst : HS65_LH_DFPRQX9 port map( D => n1470, CP => clk, RN
                           => n2789, Q => registers_2_4_port);
   registers_reg_2_3_inst : HS65_LH_DFPRQX9 port map( D => n1469, CP => clk, RN
                           => n2789, Q => registers_2_3_port);
   registers_reg_2_2_inst : HS65_LH_DFPRQX9 port map( D => n1468, CP => clk, RN
                           => n2789, Q => registers_2_2_port);
   registers_reg_2_1_inst : HS65_LH_DFPRQX9 port map( D => n1467, CP => clk, RN
                           => n2789, Q => registers_2_1_port);
   registers_reg_2_0_inst : HS65_LH_DFPRQX9 port map( D => n1466, CP => clk, RN
                           => n2789, Q => registers_2_0_port);
   registers_reg_1_31_inst : HS65_LH_DFPRQX9 port map( D => n1465, CP => clk, 
                           RN => n2789, Q => registers_1_31_port);
   registers_reg_1_30_inst : HS65_LH_DFPRQX9 port map( D => n1464, CP => clk, 
                           RN => n2789, Q => registers_1_30_port);
   registers_reg_1_29_inst : HS65_LH_DFPRQX9 port map( D => n1463, CP => clk, 
                           RN => n2789, Q => registers_1_29_port);
   registers_reg_1_28_inst : HS65_LH_DFPRQX9 port map( D => n1462, CP => clk, 
                           RN => n2789, Q => registers_1_28_port);
   registers_reg_1_27_inst : HS65_LH_DFPRQX9 port map( D => n1461, CP => clk, 
                           RN => n2789, Q => registers_1_27_port);
   registers_reg_1_26_inst : HS65_LH_DFPRQX9 port map( D => n1460, CP => clk, 
                           RN => n2789, Q => registers_1_26_port);
   registers_reg_1_25_inst : HS65_LH_DFPRQX9 port map( D => n1459, CP => clk, 
                           RN => n2790, Q => registers_1_25_port);
   registers_reg_1_24_inst : HS65_LH_DFPRQX9 port map( D => n1458, CP => clk, 
                           RN => n2790, Q => registers_1_24_port);
   registers_reg_1_23_inst : HS65_LH_DFPRQX9 port map( D => n1457, CP => clk, 
                           RN => n2790, Q => registers_1_23_port);
   registers_reg_1_22_inst : HS65_LH_DFPRQX9 port map( D => n1456, CP => clk, 
                           RN => n2790, Q => registers_1_22_port);
   registers_reg_1_21_inst : HS65_LH_DFPRQX9 port map( D => n1455, CP => clk, 
                           RN => n2790, Q => registers_1_21_port);
   registers_reg_1_20_inst : HS65_LH_DFPRQX9 port map( D => n1454, CP => clk, 
                           RN => n2790, Q => registers_1_20_port);
   registers_reg_1_19_inst : HS65_LH_DFPRQX9 port map( D => n1453, CP => clk, 
                           RN => n2790, Q => registers_1_19_port);
   registers_reg_1_18_inst : HS65_LH_DFPRQX9 port map( D => n1452, CP => clk, 
                           RN => n2790, Q => registers_1_18_port);
   registers_reg_1_17_inst : HS65_LH_DFPRQX9 port map( D => n1451, CP => clk, 
                           RN => n2790, Q => registers_1_17_port);
   registers_reg_1_16_inst : HS65_LH_DFPRQX9 port map( D => n1450, CP => clk, 
                           RN => n2790, Q => registers_1_16_port);
   registers_reg_1_15_inst : HS65_LH_DFPRQX9 port map( D => n1449, CP => clk, 
                           RN => n2790, Q => registers_1_15_port);
   registers_reg_1_14_inst : HS65_LH_DFPRQX9 port map( D => n1448, CP => clk, 
                           RN => n2790, Q => registers_1_14_port);
   registers_reg_1_13_inst : HS65_LH_DFPRQX9 port map( D => n1447, CP => clk, 
                           RN => n2791, Q => registers_1_13_port);
   registers_reg_1_12_inst : HS65_LH_DFPRQX9 port map( D => n1446, CP => clk, 
                           RN => n2791, Q => registers_1_12_port);
   registers_reg_1_11_inst : HS65_LH_DFPRQX9 port map( D => n1445, CP => clk, 
                           RN => n2791, Q => registers_1_11_port);
   registers_reg_1_10_inst : HS65_LH_DFPRQX9 port map( D => n1444, CP => clk, 
                           RN => n2791, Q => registers_1_10_port);
   registers_reg_1_9_inst : HS65_LH_DFPRQX9 port map( D => n1443, CP => clk, RN
                           => n2791, Q => registers_1_9_port);
   registers_reg_1_8_inst : HS65_LH_DFPRQX9 port map( D => n1442, CP => clk, RN
                           => n2791, Q => registers_1_8_port);
   registers_reg_1_7_inst : HS65_LH_DFPRQX9 port map( D => n1441, CP => clk, RN
                           => n2791, Q => registers_1_7_port);
   registers_reg_1_6_inst : HS65_LH_DFPRQX9 port map( D => n1440, CP => clk, RN
                           => n2791, Q => registers_1_6_port);
   registers_reg_1_5_inst : HS65_LH_DFPRQX9 port map( D => n1439, CP => clk, RN
                           => n2791, Q => registers_1_5_port);
   registers_reg_1_4_inst : HS65_LH_DFPRQX9 port map( D => n1438, CP => clk, RN
                           => n2791, Q => registers_1_4_port);
   registers_reg_1_3_inst : HS65_LH_DFPRQX9 port map( D => n1437, CP => clk, RN
                           => n2791, Q => registers_1_3_port);
   registers_reg_1_2_inst : HS65_LH_DFPRQX9 port map( D => n1436, CP => clk, RN
                           => n2791, Q => registers_1_2_port);
   registers_reg_1_1_inst : HS65_LH_DFPRQX9 port map( D => n1435, CP => clk, RN
                           => n2792, Q => registers_1_1_port);
   registers_reg_1_0_inst : HS65_LH_DFPRQX9 port map( D => n1434, CP => clk, RN
                           => n2799, Q => registers_1_0_port);
   registers_reg_29_31_inst : HS65_LH_DFPRQNX9 port map( D => n2361, CP => clk,
                           RN => n2833, QN => n1);
   registers_reg_29_30_inst : HS65_LH_DFPRQNX9 port map( D => n2360, CP => clk,
                           RN => n2833, QN => n2);
   registers_reg_29_29_inst : HS65_LH_DFPRQNX9 port map( D => n2359, CP => clk,
                           RN => n2833, QN => n3);
   registers_reg_29_28_inst : HS65_LH_DFPRQNX9 port map( D => n2358, CP => clk,
                           RN => n2832, QN => n4);
   registers_reg_29_27_inst : HS65_LH_DFPRQNX9 port map( D => n2357, CP => clk,
                           RN => n2832, QN => n5);
   registers_reg_29_26_inst : HS65_LH_DFPRQNX9 port map( D => n2356, CP => clk,
                           RN => n2832, QN => n6);
   registers_reg_29_25_inst : HS65_LH_DFPRQNX9 port map( D => n2355, CP => clk,
                           RN => n2832, QN => n7);
   registers_reg_29_24_inst : HS65_LH_DFPRQNX9 port map( D => n2354, CP => clk,
                           RN => n2832, QN => n8);
   registers_reg_29_23_inst : HS65_LH_DFPRQNX9 port map( D => n2353, CP => clk,
                           RN => n2832, QN => n9);
   registers_reg_29_22_inst : HS65_LH_DFPRQNX9 port map( D => n2352, CP => clk,
                           RN => n2832, QN => n10);
   registers_reg_29_21_inst : HS65_LH_DFPRQNX9 port map( D => n2351, CP => clk,
                           RN => n2832, QN => n11);
   registers_reg_29_20_inst : HS65_LH_DFPRQNX9 port map( D => n2350, CP => clk,
                           RN => n2832, QN => n12);
   registers_reg_29_19_inst : HS65_LH_DFPRQNX9 port map( D => n2349, CP => clk,
                           RN => n2832, QN => n13);
   registers_reg_29_18_inst : HS65_LH_DFPRQNX9 port map( D => n2348, CP => clk,
                           RN => n2832, QN => n14);
   registers_reg_29_17_inst : HS65_LH_DFPRQNX9 port map( D => n2347, CP => clk,
                           RN => n2832, QN => n15);
   registers_reg_29_16_inst : HS65_LH_DFPRQNX9 port map( D => n2346, CP => clk,
                           RN => n2832, QN => n16);
   registers_reg_29_15_inst : HS65_LH_DFPRQNX9 port map( D => n2345, CP => clk,
                           RN => n2832, QN => n17);
   registers_reg_29_14_inst : HS65_LH_DFPRQNX9 port map( D => n2344, CP => clk,
                           RN => n2831, QN => n18);
   registers_reg_29_13_inst : HS65_LH_DFPRQNX9 port map( D => n2343, CP => clk,
                           RN => n2831, QN => n19);
   registers_reg_29_12_inst : HS65_LH_DFPRQNX9 port map( D => n2342, CP => clk,
                           RN => n2831, QN => n20);
   registers_reg_29_11_inst : HS65_LH_DFPRQNX9 port map( D => n2341, CP => clk,
                           RN => n2831, QN => n21);
   registers_reg_29_10_inst : HS65_LH_DFPRQNX9 port map( D => n2340, CP => clk,
                           RN => n2831, QN => n22);
   registers_reg_29_9_inst : HS65_LH_DFPRQNX9 port map( D => n2339, CP => clk, 
                           RN => n2831, QN => n23);
   registers_reg_29_8_inst : HS65_LH_DFPRQNX9 port map( D => n2338, CP => clk, 
                           RN => n2831, QN => n24);
   registers_reg_29_7_inst : HS65_LH_DFPRQNX9 port map( D => n2337, CP => clk, 
                           RN => n2831, QN => n25);
   registers_reg_29_6_inst : HS65_LH_DFPRQNX9 port map( D => n2336, CP => clk, 
                           RN => n2831, QN => n26);
   registers_reg_29_5_inst : HS65_LH_DFPRQNX9 port map( D => n2335, CP => clk, 
                           RN => n2831, QN => n27);
   registers_reg_29_4_inst : HS65_LH_DFPRQNX9 port map( D => n2334, CP => clk, 
                           RN => n2831, QN => n28);
   registers_reg_29_3_inst : HS65_LH_DFPRQNX9 port map( D => n2333, CP => clk, 
                           RN => n2831, QN => n29);
   registers_reg_29_2_inst : HS65_LH_DFPRQNX9 port map( D => n2332, CP => clk, 
                           RN => n2831, QN => n30);
   registers_reg_29_1_inst : HS65_LH_DFPRQNX9 port map( D => n2331, CP => clk, 
                           RN => n2831, QN => n31);
   registers_reg_29_0_inst : HS65_LH_DFPRQNX9 port map( D => n2330, CP => clk, 
                           RN => n2830, QN => n32);
   registers_reg_27_31_inst : HS65_LH_DFPRQNX9 port map( D => n2297, CP => clk,
                           RN => n2826, QN => n65);
   registers_reg_27_30_inst : HS65_LH_DFPRQNX9 port map( D => n2296, CP => clk,
                           RN => n2826, QN => n66);
   registers_reg_27_29_inst : HS65_LH_DFPRQNX9 port map( D => n2295, CP => clk,
                           RN => n2827, QN => n67);
   registers_reg_27_28_inst : HS65_LH_DFPRQNX9 port map( D => n2294, CP => clk,
                           RN => n2827, QN => n68);
   registers_reg_27_27_inst : HS65_LH_DFPRQNX9 port map( D => n2293, CP => clk,
                           RN => n2827, QN => n69);
   registers_reg_27_26_inst : HS65_LH_DFPRQNX9 port map( D => n2292, CP => clk,
                           RN => n2827, QN => n70);
   registers_reg_27_25_inst : HS65_LH_DFPRQNX9 port map( D => n2291, CP => clk,
                           RN => n2827, QN => n71);
   registers_reg_27_24_inst : HS65_LH_DFPRQNX9 port map( D => n2290, CP => clk,
                           RN => n2827, QN => n72);
   registers_reg_27_23_inst : HS65_LH_DFPRQNX9 port map( D => n2289, CP => clk,
                           RN => n2827, QN => n73);
   registers_reg_27_22_inst : HS65_LH_DFPRQNX9 port map( D => n2288, CP => clk,
                           RN => n2827, QN => n74);
   registers_reg_27_21_inst : HS65_LH_DFPRQNX9 port map( D => n2287, CP => clk,
                           RN => n2827, QN => n75);
   registers_reg_27_20_inst : HS65_LH_DFPRQNX9 port map( D => n2286, CP => clk,
                           RN => n2827, QN => n76);
   registers_reg_27_19_inst : HS65_LH_DFPRQNX9 port map( D => n2285, CP => clk,
                           RN => n2827, QN => n77);
   registers_reg_27_18_inst : HS65_LH_DFPRQNX9 port map( D => n2284, CP => clk,
                           RN => n2827, QN => n78);
   registers_reg_27_17_inst : HS65_LH_DFPRQNX9 port map( D => n2283, CP => clk,
                           RN => n2827, QN => n79);
   registers_reg_27_16_inst : HS65_LH_DFPRQNX9 port map( D => n2282, CP => clk,
                           RN => n2828, QN => n80);
   registers_reg_27_15_inst : HS65_LH_DFPRQNX9 port map( D => n2281, CP => clk,
                           RN => n2828, QN => n81);
   registers_reg_27_14_inst : HS65_LH_DFPRQNX9 port map( D => n2280, CP => clk,
                           RN => n2828, QN => n82);
   registers_reg_27_13_inst : HS65_LH_DFPRQNX9 port map( D => n2279, CP => clk,
                           RN => n2828, QN => n83);
   registers_reg_27_12_inst : HS65_LH_DFPRQNX9 port map( D => n2278, CP => clk,
                           RN => n2828, QN => n84);
   registers_reg_27_11_inst : HS65_LH_DFPRQNX9 port map( D => n2277, CP => clk,
                           RN => n2828, QN => n85);
   registers_reg_27_10_inst : HS65_LH_DFPRQNX9 port map( D => n2276, CP => clk,
                           RN => n2828, QN => n86);
   registers_reg_27_9_inst : HS65_LH_DFPRQNX9 port map( D => n2275, CP => clk, 
                           RN => n2828, QN => n87);
   registers_reg_27_8_inst : HS65_LH_DFPRQNX9 port map( D => n2274, CP => clk, 
                           RN => n2828, QN => n88);
   registers_reg_27_7_inst : HS65_LH_DFPRQNX9 port map( D => n2273, CP => clk, 
                           RN => n2828, QN => n89);
   registers_reg_27_6_inst : HS65_LH_DFPRQNX9 port map( D => n2272, CP => clk, 
                           RN => n2828, QN => n90);
   registers_reg_27_5_inst : HS65_LH_DFPRQNX9 port map( D => n2271, CP => clk, 
                           RN => n2828, QN => n91);
   registers_reg_27_4_inst : HS65_LH_DFPRQNX9 port map( D => n2270, CP => clk, 
                           RN => n2828, QN => n92);
   registers_reg_27_3_inst : HS65_LH_DFPRQNX9 port map( D => n2269, CP => clk, 
                           RN => n2828, QN => n93);
   registers_reg_27_2_inst : HS65_LH_DFPRQNX9 port map( D => n2268, CP => clk, 
                           RN => n2829, QN => n94);
   registers_reg_27_1_inst : HS65_LH_DFPRQNX9 port map( D => n2267, CP => clk, 
                           RN => n2829, QN => n95);
   registers_reg_27_0_inst : HS65_LH_DFPRQNX9 port map( D => n2266, CP => clk, 
                           RN => n2829, QN => n96);
   registers_reg_15_31_inst : HS65_LH_DFPRQNX9 port map( D => n1913, CP => clk,
                           RN => n2842, QN => n129);
   registers_reg_15_30_inst : HS65_LH_DFPRQNX9 port map( D => n1912, CP => clk,
                           RN => n2842, QN => n130);
   registers_reg_15_29_inst : HS65_LH_DFPRQNX9 port map( D => n1911, CP => clk,
                           RN => n2842, QN => n131);
   registers_reg_15_28_inst : HS65_LH_DFPRQNX9 port map( D => n1910, CP => clk,
                           RN => n2842, QN => n132);
   registers_reg_15_27_inst : HS65_LH_DFPRQNX9 port map( D => n1909, CP => clk,
                           RN => n2841, QN => n133);
   registers_reg_15_26_inst : HS65_LH_DFPRQNX9 port map( D => n1908, CP => clk,
                           RN => n2841, QN => n134);
   registers_reg_15_25_inst : HS65_LH_DFPRQNX9 port map( D => n1907, CP => clk,
                           RN => n2841, QN => n135);
   registers_reg_15_24_inst : HS65_LH_DFPRQNX9 port map( D => n1906, CP => clk,
                           RN => n2841, QN => n136);
   registers_reg_15_23_inst : HS65_LH_DFPRQNX9 port map( D => n1905, CP => clk,
                           RN => n2841, QN => n137);
   registers_reg_15_22_inst : HS65_LH_DFPRQNX9 port map( D => n1904, CP => clk,
                           RN => n2841, QN => n138);
   registers_reg_15_21_inst : HS65_LH_DFPRQNX9 port map( D => n1903, CP => clk,
                           RN => n2841, QN => n139);
   registers_reg_15_20_inst : HS65_LH_DFPRQNX9 port map( D => n1902, CP => clk,
                           RN => n2841, QN => n140);
   registers_reg_15_19_inst : HS65_LH_DFPRQNX9 port map( D => n1901, CP => clk,
                           RN => n2841, QN => n141);
   registers_reg_15_18_inst : HS65_LH_DFPRQNX9 port map( D => n1900, CP => clk,
                           RN => n2841, QN => n142);
   registers_reg_15_17_inst : HS65_LH_DFPRQNX9 port map( D => n1899, CP => clk,
                           RN => n2841, QN => n143);
   registers_reg_15_16_inst : HS65_LH_DFPRQNX9 port map( D => n1898, CP => clk,
                           RN => n2841, QN => n144);
   registers_reg_15_15_inst : HS65_LH_DFPRQNX9 port map( D => n1897, CP => clk,
                           RN => n2841, QN => n145);
   registers_reg_15_14_inst : HS65_LH_DFPRQNX9 port map( D => n1896, CP => clk,
                           RN => n2836, QN => n146);
   registers_reg_15_13_inst : HS65_LH_DFPRQNX9 port map( D => n1895, CP => clk,
                           RN => n2836, QN => n147);
   registers_reg_15_12_inst : HS65_LH_DFPRQNX9 port map( D => n1894, CP => clk,
                           RN => n2836, QN => n148);
   registers_reg_15_11_inst : HS65_LH_DFPRQNX9 port map( D => n1893, CP => clk,
                           RN => n2836, QN => n149);
   registers_reg_15_10_inst : HS65_LH_DFPRQNX9 port map( D => n1892, CP => clk,
                           RN => n2836, QN => n150);
   registers_reg_15_9_inst : HS65_LH_DFPRQNX9 port map( D => n1891, CP => clk, 
                           RN => n2836, QN => n151);
   registers_reg_15_8_inst : HS65_LH_DFPRQNX9 port map( D => n1890, CP => clk, 
                           RN => n2836, QN => n152);
   registers_reg_15_7_inst : HS65_LH_DFPRQNX9 port map( D => n1889, CP => clk, 
                           RN => n2835, QN => n153);
   registers_reg_15_6_inst : HS65_LH_DFPRQNX9 port map( D => n1888, CP => clk, 
                           RN => n2835, QN => n154);
   registers_reg_15_5_inst : HS65_LH_DFPRQNX9 port map( D => n1887, CP => clk, 
                           RN => n2835, QN => n155);
   registers_reg_15_4_inst : HS65_LH_DFPRQNX9 port map( D => n1886, CP => clk, 
                           RN => n2835, QN => n156);
   registers_reg_15_3_inst : HS65_LH_DFPRQNX9 port map( D => n1885, CP => clk, 
                           RN => n2835, QN => n157);
   registers_reg_15_2_inst : HS65_LH_DFPRQNX9 port map( D => n1884, CP => clk, 
                           RN => n2835, QN => n158);
   registers_reg_15_1_inst : HS65_LH_DFPRQNX9 port map( D => n1883, CP => clk, 
                           RN => n2835, QN => n159);
   registers_reg_15_0_inst : HS65_LH_DFPRQNX9 port map( D => n1882, CP => clk, 
                           RN => n2835, QN => n160);
   registers_reg_9_31_inst : HS65_LH_DFPRQNX9 port map( D => n1721, CP => clk, 
                           RN => n2836, QN => n193);
   registers_reg_9_30_inst : HS65_LH_DFPRQNX9 port map( D => n1720, CP => clk, 
                           RN => n2836, QN => n194);
   registers_reg_9_29_inst : HS65_LH_DFPRQNX9 port map( D => n1719, CP => clk, 
                           RN => n2836, QN => n195);
   registers_reg_9_28_inst : HS65_LH_DFPRQNX9 port map( D => n1718, CP => clk, 
                           RN => n2836, QN => n196);
   registers_reg_9_27_inst : HS65_LH_DFPRQNX9 port map( D => n1717, CP => clk, 
                           RN => n2836, QN => n197);
   registers_reg_9_26_inst : HS65_LH_DFPRQNX9 port map( D => n1716, CP => clk, 
                           RN => n2836, QN => n198);
   registers_reg_9_25_inst : HS65_LH_DFPRQNX9 port map( D => n1715, CP => clk, 
                           RN => n2833, QN => n199);
   registers_reg_9_24_inst : HS65_LH_DFPRQNX9 port map( D => n1714, CP => clk, 
                           RN => n2836, QN => n200);
   registers_reg_9_23_inst : HS65_LH_DFPRQNX9 port map( D => n1713, CP => clk, 
                           RN => n2837, QN => n201);
   registers_reg_9_22_inst : HS65_LH_DFPRQNX9 port map( D => n1712, CP => clk, 
                           RN => n2837, QN => n202);
   registers_reg_9_21_inst : HS65_LH_DFPRQNX9 port map( D => n1711, CP => clk, 
                           RN => n2837, QN => n203);
   registers_reg_9_20_inst : HS65_LH_DFPRQNX9 port map( D => n1710, CP => clk, 
                           RN => n2837, QN => n204);
   registers_reg_9_19_inst : HS65_LH_DFPRQNX9 port map( D => n1709, CP => clk, 
                           RN => n2837, QN => n205);
   registers_reg_9_18_inst : HS65_LH_DFPRQNX9 port map( D => n1708, CP => clk, 
                           RN => n2837, QN => n206);
   registers_reg_9_17_inst : HS65_LH_DFPRQNX9 port map( D => n1707, CP => clk, 
                           RN => n2837, QN => n207);
   registers_reg_9_16_inst : HS65_LH_DFPRQNX9 port map( D => n1706, CP => clk, 
                           RN => n2837, QN => n208);
   registers_reg_9_15_inst : HS65_LH_DFPRQNX9 port map( D => n1705, CP => clk, 
                           RN => n2837, QN => n209);
   registers_reg_9_14_inst : HS65_LH_DFPRQNX9 port map( D => n1704, CP => clk, 
                           RN => n2837, QN => n210);
   registers_reg_9_13_inst : HS65_LH_DFPRQNX9 port map( D => n1703, CP => clk, 
                           RN => n2837, QN => n211);
   registers_reg_9_12_inst : HS65_LH_DFPRQNX9 port map( D => n1702, CP => clk, 
                           RN => n2837, QN => n212);
   registers_reg_9_11_inst : HS65_LH_DFPRQNX9 port map( D => n1701, CP => clk, 
                           RN => n2837, QN => n213);
   registers_reg_9_10_inst : HS65_LH_DFPRQNX9 port map( D => n1700, CP => clk, 
                           RN => n2837, QN => n214);
   registers_reg_9_9_inst : HS65_LH_DFPRQNX9 port map( D => n1699, CP => clk, 
                           RN => n2838, QN => n215);
   registers_reg_9_8_inst : HS65_LH_DFPRQNX9 port map( D => n1698, CP => clk, 
                           RN => n2838, QN => n216);
   registers_reg_9_7_inst : HS65_LH_DFPRQNX9 port map( D => n1697, CP => clk, 
                           RN => n2838, QN => n217);
   registers_reg_9_6_inst : HS65_LH_DFPRQNX9 port map( D => n1696, CP => clk, 
                           RN => n2838, QN => n218);
   registers_reg_9_5_inst : HS65_LH_DFPRQNX9 port map( D => n1695, CP => clk, 
                           RN => n2838, QN => n219);
   registers_reg_9_4_inst : HS65_LH_DFPRQNX9 port map( D => n1694, CP => clk, 
                           RN => n2838, QN => n220);
   registers_reg_9_3_inst : HS65_LH_DFPRQNX9 port map( D => n1693, CP => clk, 
                           RN => n2838, QN => n221);
   registers_reg_9_2_inst : HS65_LH_DFPRQNX9 port map( D => n1692, CP => clk, 
                           RN => n2838, QN => n222);
   registers_reg_9_1_inst : HS65_LH_DFPRQNX9 port map( D => n1691, CP => clk, 
                           RN => n2838, QN => n223);
   registers_reg_9_0_inst : HS65_LH_DFPRQNX9 port map( D => n1690, CP => clk, 
                           RN => n2838, QN => n224);
   registers_reg_28_31_inst : HS65_LH_DFPRQNX9 port map( D => n2329, CP => clk,
                           RN => n2830, QN => n33);
   registers_reg_28_30_inst : HS65_LH_DFPRQNX9 port map( D => n2328, CP => clk,
                           RN => n2830, QN => n34);
   registers_reg_28_29_inst : HS65_LH_DFPRQNX9 port map( D => n2327, CP => clk,
                           RN => n2830, QN => n35);
   registers_reg_28_28_inst : HS65_LH_DFPRQNX9 port map( D => n2326, CP => clk,
                           RN => n2830, QN => n36);
   registers_reg_28_27_inst : HS65_LH_DFPRQNX9 port map( D => n2325, CP => clk,
                           RN => n2830, QN => n37);
   registers_reg_28_26_inst : HS65_LH_DFPRQNX9 port map( D => n2324, CP => clk,
                           RN => n2830, QN => n38);
   registers_reg_28_25_inst : HS65_LH_DFPRQNX9 port map( D => n2323, CP => clk,
                           RN => n2830, QN => n39);
   registers_reg_28_24_inst : HS65_LH_DFPRQNX9 port map( D => n2322, CP => clk,
                           RN => n2830, QN => n40);
   registers_reg_28_23_inst : HS65_LH_DFPRQNX9 port map( D => n2321, CP => clk,
                           RN => n2830, QN => n41);
   registers_reg_28_22_inst : HS65_LH_DFPRQNX9 port map( D => n2320, CP => clk,
                           RN => n2830, QN => n42);
   registers_reg_28_21_inst : HS65_LH_DFPRQNX9 port map( D => n2319, CP => clk,
                           RN => n2830, QN => n43);
   registers_reg_28_20_inst : HS65_LH_DFPRQNX9 port map( D => n2318, CP => clk,
                           RN => n2830, QN => n44);
   registers_reg_28_19_inst : HS65_LH_DFPRQNX9 port map( D => n2317, CP => clk,
                           RN => n2830, QN => n45);
   registers_reg_28_18_inst : HS65_LH_DFPRQNX9 port map( D => n2316, CP => clk,
                           RN => n2829, QN => n46);
   registers_reg_28_17_inst : HS65_LH_DFPRQNX9 port map( D => n2315, CP => clk,
                           RN => n2829, QN => n47);
   registers_reg_28_16_inst : HS65_LH_DFPRQNX9 port map( D => n2314, CP => clk,
                           RN => n2829, QN => n48);
   registers_reg_28_15_inst : HS65_LH_DFPRQNX9 port map( D => n2313, CP => clk,
                           RN => n2829, QN => n49);
   registers_reg_28_14_inst : HS65_LH_DFPRQNX9 port map( D => n2312, CP => clk,
                           RN => n2829, QN => n50);
   registers_reg_28_13_inst : HS65_LH_DFPRQNX9 port map( D => n2311, CP => clk,
                           RN => n2829, QN => n51);
   registers_reg_28_12_inst : HS65_LH_DFPRQNX9 port map( D => n2310, CP => clk,
                           RN => n2829, QN => n52);
   registers_reg_28_11_inst : HS65_LH_DFPRQNX9 port map( D => n2309, CP => clk,
                           RN => n2829, QN => n53);
   registers_reg_28_10_inst : HS65_LH_DFPRQNX9 port map( D => n2308, CP => clk,
                           RN => n2829, QN => n54);
   registers_reg_28_9_inst : HS65_LH_DFPRQNX9 port map( D => n2307, CP => clk, 
                           RN => n2829, QN => n55);
   registers_reg_28_8_inst : HS65_LH_DFPRQNX9 port map( D => n2306, CP => clk, 
                           RN => n2829, QN => n56);
   registers_reg_28_7_inst : HS65_LH_DFPRQNX9 port map( D => n2305, CP => clk, 
                           RN => n2827, QN => n57);
   registers_reg_28_6_inst : HS65_LH_DFPRQNX9 port map( D => n2304, CP => clk, 
                           RN => n2826, QN => n58);
   registers_reg_28_5_inst : HS65_LH_DFPRQNX9 port map( D => n2303, CP => clk, 
                           RN => n2826, QN => n59);
   registers_reg_28_4_inst : HS65_LH_DFPRQNX9 port map( D => n2302, CP => clk, 
                           RN => n2826, QN => n60);
   registers_reg_28_3_inst : HS65_LH_DFPRQNX9 port map( D => n2301, CP => clk, 
                           RN => n2826, QN => n61);
   registers_reg_28_2_inst : HS65_LH_DFPRQNX9 port map( D => n2300, CP => clk, 
                           RN => n2826, QN => n62);
   registers_reg_28_1_inst : HS65_LH_DFPRQNX9 port map( D => n2299, CP => clk, 
                           RN => n2826, QN => n63);
   registers_reg_28_0_inst : HS65_LH_DFPRQNX9 port map( D => n2298, CP => clk, 
                           RN => n2826, QN => n64);
   registers_reg_26_31_inst : HS65_LH_DFPRQNX9 port map( D => n2265, CP => clk,
                           RN => n2844, QN => n97);
   registers_reg_26_30_inst : HS65_LH_DFPRQNX9 port map( D => n2264, CP => clk,
                           RN => n2844, QN => n98);
   registers_reg_26_29_inst : HS65_LH_DFPRQNX9 port map( D => n2263, CP => clk,
                           RN => n2844, QN => n99);
   registers_reg_26_28_inst : HS65_LH_DFPRQNX9 port map( D => n2262, CP => clk,
                           RN => n2844, QN => n100);
   registers_reg_26_27_inst : HS65_LH_DFPRQNX9 port map( D => n2261, CP => clk,
                           RN => n2844, QN => n101);
   registers_reg_26_26_inst : HS65_LH_DFPRQNX9 port map( D => n2260, CP => clk,
                           RN => n2844, QN => n102);
   registers_reg_26_25_inst : HS65_LH_DFPRQNX9 port map( D => n2259, CP => clk,
                           RN => n2844, QN => n103);
   registers_reg_26_24_inst : HS65_LH_DFPRQNX9 port map( D => n2258, CP => clk,
                           RN => n2844, QN => n104);
   registers_reg_26_23_inst : HS65_LH_DFPRQNX9 port map( D => n2257, CP => clk,
                           RN => n2843, QN => n105);
   registers_reg_26_22_inst : HS65_LH_DFPRQNX9 port map( D => n2256, CP => clk,
                           RN => n2843, QN => n106);
   registers_reg_26_21_inst : HS65_LH_DFPRQNX9 port map( D => n2255, CP => clk,
                           RN => n2843, QN => n107);
   registers_reg_26_20_inst : HS65_LH_DFPRQNX9 port map( D => n2254, CP => clk,
                           RN => n2843, QN => n108);
   registers_reg_26_19_inst : HS65_LH_DFPRQNX9 port map( D => n2253, CP => clk,
                           RN => n2843, QN => n109);
   registers_reg_26_18_inst : HS65_LH_DFPRQNX9 port map( D => n2252, CP => clk,
                           RN => n2843, QN => n110);
   registers_reg_26_17_inst : HS65_LH_DFPRQNX9 port map( D => n2251, CP => clk,
                           RN => n2843, QN => n111);
   registers_reg_26_16_inst : HS65_LH_DFPRQNX9 port map( D => n2250, CP => clk,
                           RN => n2843, QN => n112);
   registers_reg_26_15_inst : HS65_LH_DFPRQNX9 port map( D => n2249, CP => clk,
                           RN => n2843, QN => n113);
   registers_reg_26_14_inst : HS65_LH_DFPRQNX9 port map( D => n2248, CP => clk,
                           RN => n2843, QN => n114);
   registers_reg_26_13_inst : HS65_LH_DFPRQNX9 port map( D => n2247, CP => clk,
                           RN => n2843, QN => n115);
   registers_reg_26_12_inst : HS65_LH_DFPRQNX9 port map( D => n2246, CP => clk,
                           RN => n2843, QN => n116);
   registers_reg_26_11_inst : HS65_LH_DFPRQNX9 port map( D => n2245, CP => clk,
                           RN => n2843, QN => n117);
   registers_reg_26_10_inst : HS65_LH_DFPRQNX9 port map( D => n2244, CP => clk,
                           RN => n2843, QN => n118);
   registers_reg_26_9_inst : HS65_LH_DFPRQNX9 port map( D => n2243, CP => clk, 
                           RN => n2842, QN => n119);
   registers_reg_26_8_inst : HS65_LH_DFPRQNX9 port map( D => n2242, CP => clk, 
                           RN => n2842, QN => n120);
   registers_reg_26_7_inst : HS65_LH_DFPRQNX9 port map( D => n2241, CP => clk, 
                           RN => n2842, QN => n121);
   registers_reg_26_6_inst : HS65_LH_DFPRQNX9 port map( D => n2240, CP => clk, 
                           RN => n2842, QN => n122);
   registers_reg_26_5_inst : HS65_LH_DFPRQNX9 port map( D => n2239, CP => clk, 
                           RN => n2842, QN => n123);
   registers_reg_26_4_inst : HS65_LH_DFPRQNX9 port map( D => n2238, CP => clk, 
                           RN => n2842, QN => n124);
   registers_reg_26_3_inst : HS65_LH_DFPRQNX9 port map( D => n2237, CP => clk, 
                           RN => n2842, QN => n125);
   registers_reg_26_2_inst : HS65_LH_DFPRQNX9 port map( D => n2236, CP => clk, 
                           RN => n2842, QN => n126);
   registers_reg_26_1_inst : HS65_LH_DFPRQNX9 port map( D => n2235, CP => clk, 
                           RN => n2842, QN => n127);
   registers_reg_26_0_inst : HS65_LH_DFPRQNX9 port map( D => n2234, CP => clk, 
                           RN => n2842, QN => n128);
   registers_reg_14_31_inst : HS65_LH_DFPRQNX9 port map( D => n1881, CP => clk,
                           RN => n2835, QN => n161);
   registers_reg_14_30_inst : HS65_LH_DFPRQNX9 port map( D => n1880, CP => clk,
                           RN => n2835, QN => n162);
   registers_reg_14_29_inst : HS65_LH_DFPRQNX9 port map( D => n1879, CP => clk,
                           RN => n2835, QN => n163);
   registers_reg_14_28_inst : HS65_LH_DFPRQNX9 port map( D => n1878, CP => clk,
                           RN => n2835, QN => n164);
   registers_reg_14_27_inst : HS65_LH_DFPRQNX9 port map( D => n1877, CP => clk,
                           RN => n2835, QN => n165);
   registers_reg_14_26_inst : HS65_LH_DFPRQNX9 port map( D => n1876, CP => clk,
                           RN => n2835, QN => n166);
   registers_reg_14_25_inst : HS65_LH_DFPRQNX9 port map( D => n1875, CP => clk,
                           RN => n2834, QN => n167);
   registers_reg_14_24_inst : HS65_LH_DFPRQNX9 port map( D => n1874, CP => clk,
                           RN => n2834, QN => n168);
   registers_reg_14_23_inst : HS65_LH_DFPRQNX9 port map( D => n1873, CP => clk,
                           RN => n2834, QN => n169);
   registers_reg_14_22_inst : HS65_LH_DFPRQNX9 port map( D => n1872, CP => clk,
                           RN => n2834, QN => n170);
   registers_reg_14_21_inst : HS65_LH_DFPRQNX9 port map( D => n1871, CP => clk,
                           RN => n2834, QN => n171);
   registers_reg_14_20_inst : HS65_LH_DFPRQNX9 port map( D => n1870, CP => clk,
                           RN => n2834, QN => n172);
   registers_reg_14_19_inst : HS65_LH_DFPRQNX9 port map( D => n1869, CP => clk,
                           RN => n2834, QN => n173);
   registers_reg_14_18_inst : HS65_LH_DFPRQNX9 port map( D => n1868, CP => clk,
                           RN => n2834, QN => n174);
   registers_reg_14_17_inst : HS65_LH_DFPRQNX9 port map( D => n1867, CP => clk,
                           RN => n2834, QN => n175);
   registers_reg_14_16_inst : HS65_LH_DFPRQNX9 port map( D => n1866, CP => clk,
                           RN => n2834, QN => n176);
   registers_reg_14_15_inst : HS65_LH_DFPRQNX9 port map( D => n1865, CP => clk,
                           RN => n2834, QN => n177);
   registers_reg_14_14_inst : HS65_LH_DFPRQNX9 port map( D => n1864, CP => clk,
                           RN => n2834, QN => n178);
   registers_reg_14_13_inst : HS65_LH_DFPRQNX9 port map( D => n1863, CP => clk,
                           RN => n2834, QN => n179);
   registers_reg_14_12_inst : HS65_LH_DFPRQNX9 port map( D => n1862, CP => clk,
                           RN => n2834, QN => n180);
   registers_reg_14_11_inst : HS65_LH_DFPRQNX9 port map( D => n1861, CP => clk,
                           RN => n2833, QN => n181);
   registers_reg_14_10_inst : HS65_LH_DFPRQNX9 port map( D => n1860, CP => clk,
                           RN => n2833, QN => n182);
   registers_reg_14_9_inst : HS65_LH_DFPRQNX9 port map( D => n1859, CP => clk, 
                           RN => n2833, QN => n183);
   registers_reg_14_8_inst : HS65_LH_DFPRQNX9 port map( D => n1858, CP => clk, 
                           RN => n2833, QN => n184);
   registers_reg_14_7_inst : HS65_LH_DFPRQNX9 port map( D => n1857, CP => clk, 
                           RN => n2833, QN => n185);
   registers_reg_14_6_inst : HS65_LH_DFPRQNX9 port map( D => n1856, CP => clk, 
                           RN => n2833, QN => n186);
   registers_reg_14_5_inst : HS65_LH_DFPRQNX9 port map( D => n1855, CP => clk, 
                           RN => n2833, QN => n187);
   registers_reg_14_4_inst : HS65_LH_DFPRQNX9 port map( D => n1854, CP => clk, 
                           RN => n2833, QN => n188);
   registers_reg_14_3_inst : HS65_LH_DFPRQNX9 port map( D => n1853, CP => clk, 
                           RN => n2833, QN => n189);
   registers_reg_14_2_inst : HS65_LH_DFPRQNX9 port map( D => n1852, CP => clk, 
                           RN => n2833, QN => n190);
   registers_reg_14_1_inst : HS65_LH_DFPRQNX9 port map( D => n1851, CP => clk, 
                           RN => n2838, QN => n191);
   registers_reg_14_0_inst : HS65_LH_DFPRQNX9 port map( D => n1850, CP => clk, 
                           RN => n2826, QN => n192);
   registers_reg_8_31_inst : HS65_LH_DFPRQNX9 port map( D => n1689, CP => clk, 
                           RN => n2838, QN => n225);
   registers_reg_8_30_inst : HS65_LH_DFPRQNX9 port map( D => n1688, CP => clk, 
                           RN => n2838, QN => n226);
   registers_reg_8_29_inst : HS65_LH_DFPRQNX9 port map( D => n1687, CP => clk, 
                           RN => n2838, QN => n227);
   registers_reg_8_28_inst : HS65_LH_DFPRQNX9 port map( D => n1686, CP => clk, 
                           RN => n2839, QN => n228);
   registers_reg_8_27_inst : HS65_LH_DFPRQNX9 port map( D => n1685, CP => clk, 
                           RN => n2839, QN => n229);
   registers_reg_8_26_inst : HS65_LH_DFPRQNX9 port map( D => n1684, CP => clk, 
                           RN => n2839, QN => n230);
   registers_reg_8_25_inst : HS65_LH_DFPRQNX9 port map( D => n1683, CP => clk, 
                           RN => n2839, QN => n231);
   registers_reg_8_24_inst : HS65_LH_DFPRQNX9 port map( D => n1682, CP => clk, 
                           RN => n2839, QN => n232);
   registers_reg_8_23_inst : HS65_LH_DFPRQNX9 port map( D => n1681, CP => clk, 
                           RN => n2839, QN => n233);
   registers_reg_8_22_inst : HS65_LH_DFPRQNX9 port map( D => n1680, CP => clk, 
                           RN => n2839, QN => n234);
   registers_reg_8_21_inst : HS65_LH_DFPRQNX9 port map( D => n1679, CP => clk, 
                           RN => n2839, QN => n235);
   registers_reg_8_20_inst : HS65_LH_DFPRQNX9 port map( D => n1678, CP => clk, 
                           RN => n2839, QN => n236);
   registers_reg_8_19_inst : HS65_LH_DFPRQNX9 port map( D => n1677, CP => clk, 
                           RN => n2839, QN => n237);
   registers_reg_8_18_inst : HS65_LH_DFPRQNX9 port map( D => n1676, CP => clk, 
                           RN => n2839, QN => n238);
   registers_reg_8_17_inst : HS65_LH_DFPRQNX9 port map( D => n1675, CP => clk, 
                           RN => n2839, QN => n239);
   registers_reg_8_16_inst : HS65_LH_DFPRQNX9 port map( D => n1674, CP => clk, 
                           RN => n2839, QN => n240);
   registers_reg_8_15_inst : HS65_LH_DFPRQNX9 port map( D => n1673, CP => clk, 
                           RN => n2839, QN => n241);
   registers_reg_8_14_inst : HS65_LH_DFPRQNX9 port map( D => n1672, CP => clk, 
                           RN => n2840, QN => n242);
   registers_reg_8_13_inst : HS65_LH_DFPRQNX9 port map( D => n1671, CP => clk, 
                           RN => n2840, QN => n243);
   registers_reg_8_12_inst : HS65_LH_DFPRQNX9 port map( D => n1670, CP => clk, 
                           RN => n2840, QN => n244);
   registers_reg_8_11_inst : HS65_LH_DFPRQNX9 port map( D => n1669, CP => clk, 
                           RN => n2840, QN => n245);
   registers_reg_8_10_inst : HS65_LH_DFPRQNX9 port map( D => n1668, CP => clk, 
                           RN => n2840, QN => n246);
   registers_reg_8_9_inst : HS65_LH_DFPRQNX9 port map( D => n1667, CP => clk, 
                           RN => n2840, QN => n247);
   registers_reg_8_8_inst : HS65_LH_DFPRQNX9 port map( D => n1666, CP => clk, 
                           RN => n2840, QN => n248);
   registers_reg_8_7_inst : HS65_LH_DFPRQNX9 port map( D => n1665, CP => clk, 
                           RN => n2840, QN => n249);
   registers_reg_8_6_inst : HS65_LH_DFPRQNX9 port map( D => n1664, CP => clk, 
                           RN => n2840, QN => n250);
   registers_reg_8_5_inst : HS65_LH_DFPRQNX9 port map( D => n1663, CP => clk, 
                           RN => n2840, QN => n251);
   registers_reg_8_4_inst : HS65_LH_DFPRQNX9 port map( D => n1662, CP => clk, 
                           RN => n2840, QN => n252);
   registers_reg_8_3_inst : HS65_LH_DFPRQNX9 port map( D => n1661, CP => clk, 
                           RN => n2840, QN => n253);
   registers_reg_8_2_inst : HS65_LH_DFPRQNX9 port map( D => n1660, CP => clk, 
                           RN => n2840, QN => n254);
   registers_reg_8_1_inst : HS65_LH_DFPRQNX9 port map( D => n1659, CP => clk, 
                           RN => n2840, QN => n255);
   registers_reg_8_0_inst : HS65_LH_DFPRQNX9 port map( D => n1658, CP => clk, 
                           RN => n2841, QN => n256);
   U3 : HS65_LH_AND2X4 port map( A => n1393, B => n1394, Z => n257);
   U4 : HS65_LH_AND2X4 port map( A => n1396, B => n1394, Z => n258);
   U5 : HS65_LH_AND2X4 port map( A => n1398, B => n1394, Z => n259);
   U6 : HS65_LH_AND2X4 port map( A => n1406, B => n1394, Z => n260);
   U7 : HS65_LH_AND2X4 port map( A => n1402, B => n1394, Z => n261);
   U8 : HS65_LH_AND2X4 port map( A => n1404, B => n1394, Z => n262);
   U9 : HS65_LH_AND2X4 port map( A => n1400, B => n1394, Z => n263);
   U10 : HS65_LH_AND2X4 port map( A => n1408, B => n1398, Z => n264);
   U11 : HS65_LH_AND2X4 port map( A => n1408, B => n1402, Z => n265);
   U12 : HS65_LH_AND2X4 port map( A => n1408, B => n1396, Z => n266);
   U13 : HS65_LH_AND2X4 port map( A => n1408, B => n1400, Z => n267);
   U14 : HS65_LH_AND2X4 port map( A => n1417, B => n1402, Z => n268);
   U15 : HS65_LH_AND2X4 port map( A => n1417, B => n1400, Z => n269);
   U16 : HS65_LH_AND2X4 port map( A => n1426, B => n1404, Z => n270);
   U17 : HS65_LH_AND2X4 port map( A => n1417, B => n1404, Z => n271);
   U18 : HS65_LH_AND2X4 port map( A => n1426, B => n1406, Z => n272);
   U19 : HS65_LH_AND2X4 port map( A => n1417, B => n1406, Z => n273);
   U20 : HS65_LH_AND2X4 port map( A => n1426, B => n1393, Z => n274);
   U21 : HS65_LH_AND2X4 port map( A => n1417, B => n1398, Z => n275);
   U22 : HS65_LH_AND2X4 port map( A => n1417, B => n1393, Z => n276);
   U23 : HS65_LH_AND2X4 port map( A => n1417, B => n1396, Z => n277);
   U24 : HS65_LH_AND2X4 port map( A => n861, B => n841, Z => n380);
   U25 : HS65_LH_AND2X4 port map( A => n849, B => n841, Z => n358);
   U26 : HS65_LH_AND2X4 port map( A => n1389, B => n1369, Z => n908);
   U27 : HS65_LH_AND2X4 port map( A => n1377, B => n1369, Z => n886);
   U28 : HS65_LH_AND2X4 port map( A => n857, B => n841, Z => n365);
   U29 : HS65_LH_AND2X4 port map( A => n1385, B => n1369, Z => n893);
   U30 : HS65_LH_AND2X4 port map( A => n861, B => n843, Z => n378);
   U31 : HS65_LH_AND2X4 port map( A => n860, B => n843, Z => n379);
   U32 : HS65_LH_AND2X4 port map( A => n861, B => n846, Z => n376);
   U33 : HS65_LH_AND2X4 port map( A => n860, B => n846, Z => n377);
   U34 : HS65_LH_AND2X4 port map( A => n849, B => n843, Z => n356);
   U35 : HS65_LH_AND2X4 port map( A => n848, B => n843, Z => n357);
   U36 : HS65_LH_AND2X4 port map( A => n1389, B => n1371, Z => n906);
   U37 : HS65_LH_AND2X4 port map( A => n1388, B => n1371, Z => n907);
   U38 : HS65_LH_AND2X4 port map( A => n1389, B => n1374, Z => n904);
   U39 : HS65_LH_AND2X4 port map( A => n1388, B => n1374, Z => n905);
   U40 : HS65_LH_AND2X4 port map( A => n1377, B => n1371, Z => n884);
   U41 : HS65_LH_AND2X4 port map( A => n1376, B => n1371, Z => n885);
   U42 : HS65_LH_AND2X4 port map( A => n1368, B => n1374, Z => n875);
   U43 : HS65_LH_AND2X4 port map( A => n860, B => n841, Z => n381);
   U44 : HS65_LH_AND2X4 port map( A => n1388, B => n1369, Z => n909);
   U45 : HS65_LH_AND2X4 port map( A => n1376, B => n1369, Z => n887);
   U46 : HS65_LH_AND2X4 port map( A => n861, B => n845, Z => n374);
   U47 : HS65_LH_AND2X4 port map( A => n860, B => n845, Z => n375);
   U48 : HS65_LH_AND2X4 port map( A => n1389, B => n1373, Z => n902);
   U49 : HS65_LH_AND2X4 port map( A => n1388, B => n1373, Z => n903);
   U50 : HS65_LH_AND2X4 port map( A => n1373, B => n1384, Z => n897);
   U51 : HS65_LH_IVX9 port map( A => regfile_i(9), Z => n2710);
   U52 : HS65_LH_IVX9 port map( A => regfile_i(10), Z => n2712);
   U53 : HS65_LH_IVX9 port map( A => regfile_i(11), Z => n2714);
   U54 : HS65_LH_IVX9 port map( A => regfile_i(13), Z => n2718);
   U55 : HS65_LH_IVX9 port map( A => regfile_i(14), Z => n2720);
   U56 : HS65_LH_IVX9 port map( A => regfile_i(15), Z => n2722);
   U57 : HS65_LH_IVX9 port map( A => regfile_i(16), Z => n2724);
   U58 : HS65_LH_IVX9 port map( A => regfile_i(17), Z => n2726);
   U59 : HS65_LH_IVX9 port map( A => regfile_i(18), Z => n2728);
   U60 : HS65_LH_IVX9 port map( A => regfile_i(19), Z => n2730);
   U61 : HS65_LH_IVX9 port map( A => regfile_i(20), Z => n2732);
   U62 : HS65_LH_IVX9 port map( A => regfile_i(21), Z => n2734);
   U63 : HS65_LH_IVX9 port map( A => regfile_i(22), Z => n2736);
   U64 : HS65_LH_IVX9 port map( A => regfile_i(23), Z => n2738);
   U65 : HS65_LH_IVX9 port map( A => regfile_i(24), Z => n2740);
   U66 : HS65_LH_IVX9 port map( A => regfile_i(25), Z => n2742);
   U67 : HS65_LH_IVX9 port map( A => regfile_i(26), Z => n2744);
   U68 : HS65_LH_IVX9 port map( A => regfile_i(27), Z => n2746);
   U69 : HS65_LH_IVX9 port map( A => regfile_i(28), Z => n2748);
   U70 : HS65_LH_IVX9 port map( A => regfile_i(29), Z => n2750);
   U71 : HS65_LH_IVX9 port map( A => regfile_i(30), Z => n2752);
   U72 : HS65_LH_IVX9 port map( A => regfile_i(31), Z => n2754);
   U73 : HS65_LH_IVX9 port map( A => regfile_i(32), Z => n2756);
   U74 : HS65_LH_IVX9 port map( A => regfile_i(33), Z => n2758);
   U75 : HS65_LH_IVX9 port map( A => regfile_i(34), Z => n2760);
   U76 : HS65_LH_AND2X4 port map( A => n849, B => n846, Z => n354);
   U77 : HS65_LH_AND2X4 port map( A => n848, B => n846, Z => n355);
   U78 : HS65_LH_AND2X4 port map( A => n1377, B => n1374, Z => n882);
   U79 : HS65_LH_AND2X4 port map( A => n1376, B => n1374, Z => n883);
   U80 : HS65_LH_AND2X4 port map( A => n840, B => n846, Z => n347);
   U81 : HS65_LH_AND2X4 port map( A => n842, B => n846, Z => n348);
   U82 : HS65_LH_AND2X4 port map( A => n840, B => n843, Z => n342);
   U83 : HS65_LH_AND2X4 port map( A => n842, B => n843, Z => n343);
   U84 : HS65_LH_AND2X4 port map( A => n1370, B => n1374, Z => n876);
   U85 : HS65_LH_AND2X4 port map( A => n1368, B => n1371, Z => n870);
   U86 : HS65_LH_AND2X4 port map( A => n1370, B => n1371, Z => n871);
   U87 : HS65_LH_AND2X4 port map( A => n848, B => n841, Z => n359);
   U88 : HS65_LH_AND2X4 port map( A => n848, B => n845, Z => n353);
   U89 : HS65_LH_AND2X4 port map( A => n1376, B => n1373, Z => n881);
   U90 : HS65_LH_AND2X4 port map( A => n841, B => n856, Z => n364);
   U91 : HS65_LH_AND2X4 port map( A => n1369, B => n1384, Z => n892);
   U92 : HS65_LH_AND2X4 port map( A => n845, B => n856, Z => n369);
   U93 : HS65_LH_AND2X4 port map( A => n845, B => n857, Z => n370);
   U94 : HS65_LH_AND2X4 port map( A => n1373, B => n1385, Z => n898);
   U95 : HS65_LH_IVX9 port map( A => regfile_i(4), Z => n2700);
   U96 : HS65_LH_IVX9 port map( A => regfile_i(5), Z => n2702);
   U97 : HS65_LH_IVX9 port map( A => regfile_i(6), Z => n2704);
   U98 : HS65_LH_IVX9 port map( A => regfile_i(7), Z => n2706);
   U99 : HS65_LH_IVX9 port map( A => regfile_i(8), Z => n2708);
   U100 : HS65_LH_IVX9 port map( A => regfile_i(12), Z => n2716);
   U101 : HS65_LH_IVX9 port map( A => regfile_i(3), Z => n2698);
   U102 : HS65_LH_IVX9 port map( A => regfile_i(2), Z => n2893);
   U103 : HS65_LH_NOR3AX2 port map( A => regfile_i(37), B => regfile_i(35), C 
                           => regfile_i(36), Z => n1400);
   U104 : HS65_LH_NOR3AX2 port map( A => regfile_i(37), B => n2897, C => 
                           regfile_i(36), Z => n1402);
   U105 : HS65_LH_NOR3AX2 port map( A => regfile_i(37), B => n2896, C => 
                           regfile_i(35), Z => n1404);
   U106 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => regfile_i(39), C =>
                           n2895, Z => n1408);
   U107 : HS65_LH_NOR3AX2 port map( A => regfile_i(37), B => n2896, C => n2897,
                           Z => n1406);
   U108 : HS65_LH_NOR3AX2 port map( A => regfile_i(0), B => regfile_i(38), C =>
                           regfile_i(39), Z => n1394);
   U109 : HS65_LH_BFX9 port map( A => n2854, Z => n2826);
   U110 : HS65_LH_BFX9 port map( A => n2847, Z => n2840);
   U111 : HS65_LH_BFX9 port map( A => n2847, Z => n2839);
   U112 : HS65_LH_BFX9 port map( A => n2848, Z => n2837);
   U113 : HS65_LH_BFX9 port map( A => n2848, Z => n2838);
   U114 : HS65_LH_BFX9 port map( A => n2850, Z => n2834);
   U115 : HS65_LH_BFX9 port map( A => n2849, Z => n2835);
   U116 : HS65_LH_BFX9 port map( A => n2849, Z => n2836);
   U117 : HS65_LH_BFX9 port map( A => n2846, Z => n2841);
   U118 : HS65_LH_BFX9 port map( A => n2846, Z => n2842);
   U119 : HS65_LH_BFX9 port map( A => n2845, Z => n2843);
   U120 : HS65_LH_BFX9 port map( A => n2853, Z => n2828);
   U121 : HS65_LH_BFX9 port map( A => n2853, Z => n2827);
   U122 : HS65_LH_BFX9 port map( A => n2852, Z => n2829);
   U123 : HS65_LH_BFX9 port map( A => n2852, Z => n2830);
   U124 : HS65_LH_BFX9 port map( A => n2851, Z => n2831);
   U125 : HS65_LH_BFX9 port map( A => n2851, Z => n2832);
   U126 : HS65_LH_BFX9 port map( A => n2850, Z => n2833);
   U127 : HS65_LH_BFX9 port map( A => n2871, Z => n2791);
   U128 : HS65_LH_BFX9 port map( A => n2872, Z => n2790);
   U129 : HS65_LH_BFX9 port map( A => n2872, Z => n2789);
   U130 : HS65_LH_BFX9 port map( A => n2873, Z => n2788);
   U131 : HS65_LH_BFX9 port map( A => n2874, Z => n2786);
   U132 : HS65_LH_BFX9 port map( A => n2874, Z => n2785);
   U133 : HS65_LH_BFX9 port map( A => n2875, Z => n2784);
   U134 : HS65_LH_BFX9 port map( A => n2873, Z => n2787);
   U135 : HS65_LH_BFX9 port map( A => n2867, Z => n2800);
   U136 : HS65_LH_BFX9 port map( A => n2867, Z => n2799);
   U137 : HS65_LH_BFX9 port map( A => n2868, Z => n2798);
   U138 : HS65_LH_BFX9 port map( A => n2868, Z => n2797);
   U139 : HS65_LH_BFX9 port map( A => n2869, Z => n2795);
   U140 : HS65_LH_BFX9 port map( A => n2870, Z => n2794);
   U141 : HS65_LH_BFX9 port map( A => n2870, Z => n2793);
   U142 : HS65_LH_BFX9 port map( A => n2871, Z => n2792);
   U143 : HS65_LH_BFX9 port map( A => n2869, Z => n2796);
   U144 : HS65_LH_BFX9 port map( A => n2880, Z => n2773);
   U145 : HS65_LH_BFX9 port map( A => n2881, Z => n2772);
   U146 : HS65_LH_BFX9 port map( A => n2881, Z => n2771);
   U147 : HS65_LH_BFX9 port map( A => n2882, Z => n2770);
   U148 : HS65_LH_BFX9 port map( A => n2883, Z => n2768);
   U149 : HS65_LH_BFX9 port map( A => n2883, Z => n2767);
   U150 : HS65_LH_BFX9 port map( A => n2884, Z => n2766);
   U151 : HS65_LH_BFX9 port map( A => n2882, Z => n2769);
   U152 : HS65_LH_BFX9 port map( A => n2876, Z => n2782);
   U153 : HS65_LH_BFX9 port map( A => n2876, Z => n2781);
   U154 : HS65_LH_BFX9 port map( A => n2877, Z => n2780);
   U155 : HS65_LH_BFX9 port map( A => n2877, Z => n2779);
   U156 : HS65_LH_BFX9 port map( A => n2878, Z => n2777);
   U157 : HS65_LH_BFX9 port map( A => n2879, Z => n2776);
   U158 : HS65_LH_BFX9 port map( A => n2879, Z => n2775);
   U159 : HS65_LH_BFX9 port map( A => n2880, Z => n2774);
   U160 : HS65_LH_BFX9 port map( A => n2878, Z => n2778);
   U161 : HS65_LH_BFX9 port map( A => n2875, Z => n2783);
   U162 : HS65_LH_BFX9 port map( A => n2856, Z => n2822);
   U163 : HS65_LH_BFX9 port map( A => n2857, Z => n2820);
   U164 : HS65_LH_BFX9 port map( A => n2857, Z => n2819);
   U165 : HS65_LH_BFX9 port map( A => n2858, Z => n2818);
   U166 : HS65_LH_BFX9 port map( A => n2856, Z => n2821);
   U167 : HS65_LH_BFX9 port map( A => n2855, Z => n2823);
   U168 : HS65_LH_BFX9 port map( A => n2855, Z => n2824);
   U169 : HS65_LH_BFX9 port map( A => n2854, Z => n2825);
   U170 : HS65_LH_BFX9 port map( A => n2866, Z => n2801);
   U171 : HS65_LH_BFX9 port map( A => n2866, Z => n2802);
   U172 : HS65_LH_BFX9 port map( A => n2865, Z => n2803);
   U173 : HS65_LH_BFX9 port map( A => n2865, Z => n2804);
   U174 : HS65_LH_BFX9 port map( A => n2864, Z => n2805);
   U175 : HS65_LH_BFX9 port map( A => n2864, Z => n2806);
   U176 : HS65_LH_BFX9 port map( A => n2863, Z => n2807);
   U177 : HS65_LH_BFX9 port map( A => n2863, Z => n2808);
   U178 : HS65_LH_BFX9 port map( A => n2862, Z => n2809);
   U179 : HS65_LH_BFX9 port map( A => n2862, Z => n2810);
   U180 : HS65_LH_BFX9 port map( A => n2861, Z => n2811);
   U181 : HS65_LH_BFX9 port map( A => n2861, Z => n2812);
   U182 : HS65_LH_BFX9 port map( A => n2860, Z => n2813);
   U183 : HS65_LH_BFX9 port map( A => n2860, Z => n2814);
   U184 : HS65_LH_BFX9 port map( A => n2859, Z => n2815);
   U185 : HS65_LH_BFX9 port map( A => n2859, Z => n2816);
   U186 : HS65_LH_BFX9 port map( A => n2858, Z => n2817);
   U187 : HS65_LH_BFX9 port map( A => n2884, Z => n2765);
   U188 : HS65_LH_BFX9 port map( A => n2845, Z => n2844);
   U189 : HS65_LH_BFX9 port map( A => n2887, Z => n2872);
   U190 : HS65_LH_BFX9 port map( A => n2887, Z => n2874);
   U191 : HS65_LH_BFX9 port map( A => n2887, Z => n2873);
   U192 : HS65_LH_BFX9 port map( A => n2888, Z => n2867);
   U193 : HS65_LH_BFX9 port map( A => n2888, Z => n2868);
   U194 : HS65_LH_BFX9 port map( A => n2887, Z => n2870);
   U195 : HS65_LH_BFX9 port map( A => n2887, Z => n2871);
   U196 : HS65_LH_BFX9 port map( A => n2888, Z => n2869);
   U197 : HS65_LH_BFX9 port map( A => n2885, Z => n2881);
   U198 : HS65_LH_BFX9 port map( A => n2885, Z => n2883);
   U199 : HS65_LH_BFX9 port map( A => n2885, Z => n2882);
   U200 : HS65_LH_BFX9 port map( A => n2886, Z => n2876);
   U201 : HS65_LH_BFX9 port map( A => n2886, Z => n2877);
   U202 : HS65_LH_BFX9 port map( A => n2886, Z => n2879);
   U203 : HS65_LH_BFX9 port map( A => n2885, Z => n2880);
   U204 : HS65_LH_BFX9 port map( A => n2886, Z => n2878);
   U205 : HS65_LH_BFX9 port map( A => n2886, Z => n2875);
   U206 : HS65_LH_BFX9 port map( A => n2890, Z => n2857);
   U207 : HS65_LH_BFX9 port map( A => n2890, Z => n2856);
   U208 : HS65_LH_BFX9 port map( A => n2890, Z => n2855);
   U209 : HS65_LH_BFX9 port map( A => n2888, Z => n2866);
   U210 : HS65_LH_BFX9 port map( A => n2888, Z => n2865);
   U211 : HS65_LH_BFX9 port map( A => n2889, Z => n2864);
   U212 : HS65_LH_BFX9 port map( A => n2889, Z => n2863);
   U213 : HS65_LH_BFX9 port map( A => n2889, Z => n2862);
   U214 : HS65_LH_BFX9 port map( A => n2889, Z => n2861);
   U215 : HS65_LH_BFX9 port map( A => n2889, Z => n2860);
   U216 : HS65_LH_BFX9 port map( A => n2890, Z => n2859);
   U217 : HS65_LH_BFX9 port map( A => n2890, Z => n2858);
   U218 : HS65_LH_BFX9 port map( A => n2885, Z => n2884);
   U219 : HS65_LH_BFX9 port map( A => n2892, Z => n2847);
   U220 : HS65_LH_BFX9 port map( A => n2892, Z => n2848);
   U221 : HS65_LH_BFX9 port map( A => n2892, Z => n2849);
   U222 : HS65_LH_BFX9 port map( A => n2892, Z => n2846);
   U223 : HS65_LH_BFX9 port map( A => n2892, Z => n2845);
   U224 : HS65_LH_BFX9 port map( A => n2891, Z => n2854);
   U225 : HS65_LH_BFX9 port map( A => n2891, Z => n2853);
   U226 : HS65_LH_BFX9 port map( A => n2891, Z => n2852);
   U227 : HS65_LH_BFX9 port map( A => n2891, Z => n2851);
   U228 : HS65_LH_BFX9 port map( A => n2891, Z => n2850);
   U229 : HS65_LH_BFX9 port map( A => n2761, Z => n2887);
   U230 : HS65_LH_BFX9 port map( A => n2761, Z => n2886);
   U231 : HS65_LH_BFX9 port map( A => n2762, Z => n2888);
   U232 : HS65_LH_BFX9 port map( A => n2762, Z => n2889);
   U233 : HS65_LH_BFX9 port map( A => n2762, Z => n2890);
   U234 : HS65_LH_BFX9 port map( A => n2761, Z => n2885);
   U235 : HS65_LH_BFX9 port map( A => n2763, Z => n2892);
   U236 : HS65_LH_BFX9 port map( A => n2763, Z => n2891);
   U237 : HS65_LH_BFX9 port map( A => n908, Z => n2514);
   U238 : HS65_LH_BFX9 port map( A => n886, Z => n2562);
   U239 : HS65_LH_BFX9 port map( A => n908, Z => n2515);
   U240 : HS65_LH_BFX9 port map( A => n886, Z => n2563);
   U241 : HS65_LH_BFX9 port map( A => n380, Z => n2607);
   U242 : HS65_LH_BFX9 port map( A => n358, Z => n2655);
   U243 : HS65_LH_BFX9 port map( A => n380, Z => n2608);
   U244 : HS65_LH_BFX9 port map( A => n358, Z => n2656);
   U245 : HS65_LH_BFX9 port map( A => n380, Z => n2609);
   U246 : HS65_LH_BFX9 port map( A => n358, Z => n2657);
   U247 : HS65_LH_BFX9 port map( A => n908, Z => n2516);
   U248 : HS65_LH_BFX9 port map( A => n886, Z => n2564);
   U249 : HS65_LH_BFX9 port map( A => n893, Z => n2553);
   U250 : HS65_LH_BFX9 port map( A => n893, Z => n2554);
   U251 : HS65_LH_BFX9 port map( A => n345, Z => n2688);
   U252 : HS65_LH_BFX9 port map( A => n345, Z => n2689);
   U253 : HS65_LH_BFX9 port map( A => n365, Z => n2646);
   U254 : HS65_LH_BFX9 port map( A => n365, Z => n2647);
   U255 : HS65_LH_BFX9 port map( A => n873, Z => n2595);
   U256 : HS65_LH_BFX9 port map( A => n873, Z => n2596);
   U257 : HS65_LH_BFX9 port map( A => n345, Z => n2690);
   U258 : HS65_LH_BFX9 port map( A => n873, Z => n2597);
   U259 : HS65_LH_BFX9 port map( A => n893, Z => n2555);
   U260 : HS65_LH_BFX9 port map( A => n365, Z => n2648);
   U261 : HS65_LH_IVX9 port map( A => n2473, Z => n2472);
   U262 : HS65_LH_IVX9 port map( A => n2473, Z => n2471);
   U263 : HS65_LH_IVX9 port map( A => n2468, Z => n2467);
   U264 : HS65_LH_IVX9 port map( A => n2468, Z => n2466);
   U265 : HS65_LH_IVX9 port map( A => n2443, Z => n2442);
   U266 : HS65_LH_IVX9 port map( A => n2443, Z => n2441);
   U267 : HS65_LH_IVX9 port map( A => n2438, Z => n2437);
   U268 : HS65_LH_IVX9 port map( A => n2438, Z => n2436);
   U269 : HS65_LH_IVX9 port map( A => n300, Z => n299);
   U270 : HS65_LH_IVX9 port map( A => n300, Z => n298);
   U271 : HS65_LH_BFX9 port map( A => n259, Z => n2499);
   U272 : HS65_LH_BFX9 port map( A => n263, Z => n2494);
   U273 : HS65_LH_BFX9 port map( A => n261, Z => n2489);
   U274 : HS65_LH_BFX9 port map( A => n262, Z => n2484);
   U275 : HS65_LH_BFX9 port map( A => n260, Z => n2479);
   U276 : HS65_LH_BFX9 port map( A => n266, Z => n2464);
   U277 : HS65_LH_BFX9 port map( A => n264, Z => n2459);
   U278 : HS65_LH_BFX9 port map( A => n267, Z => n2454);
   U279 : HS65_LH_BFX9 port map( A => n265, Z => n2449);
   U280 : HS65_LH_BFX9 port map( A => n269, Z => n1412);
   U281 : HS65_LH_BFX9 port map( A => n268, Z => n1401);
   U282 : HS65_LH_BFX9 port map( A => n271, Z => n880);
   U283 : HS65_LH_BFX9 port map( A => n270, Z => n296);
   U284 : HS65_LH_IVX9 port map( A => n2463, Z => n2462);
   U285 : HS65_LH_IVX9 port map( A => n2463, Z => n2461);
   U286 : HS65_LH_IVX9 port map( A => n2458, Z => n2457);
   U287 : HS65_LH_IVX9 port map( A => n2458, Z => n2456);
   U288 : HS65_LH_IVX9 port map( A => n2453, Z => n2452);
   U289 : HS65_LH_IVX9 port map( A => n2453, Z => n2451);
   U290 : HS65_LH_IVX9 port map( A => n2448, Z => n2447);
   U291 : HS65_LH_IVX9 port map( A => n2448, Z => n2446);
   U292 : HS65_LH_IVX9 port map( A => n2508, Z => n2507);
   U293 : HS65_LH_IVX9 port map( A => n2508, Z => n2506);
   U294 : HS65_LH_IVX9 port map( A => n2503, Z => n2502);
   U295 : HS65_LH_IVX9 port map( A => n2503, Z => n2501);
   U296 : HS65_LH_IVX9 port map( A => n2498, Z => n2497);
   U297 : HS65_LH_IVX9 port map( A => n2498, Z => n2496);
   U298 : HS65_LH_IVX9 port map( A => n2493, Z => n2492);
   U299 : HS65_LH_IVX9 port map( A => n2493, Z => n2491);
   U300 : HS65_LH_IVX9 port map( A => n2488, Z => n2487);
   U301 : HS65_LH_IVX9 port map( A => n2488, Z => n2486);
   U302 : HS65_LH_IVX9 port map( A => n2483, Z => n2482);
   U303 : HS65_LH_IVX9 port map( A => n2483, Z => n2481);
   U304 : HS65_LH_IVX9 port map( A => n2478, Z => n2477);
   U305 : HS65_LH_IVX9 port map( A => n2478, Z => n2476);
   U306 : HS65_LH_IVX9 port map( A => n2428, Z => n2427);
   U307 : HS65_LH_IVX9 port map( A => n2428, Z => n2426);
   U308 : HS65_LH_IVX9 port map( A => n1427, Z => n1424);
   U309 : HS65_LH_IVX9 port map( A => n1427, Z => n1423);
   U310 : HS65_LH_IVX9 port map( A => n1420, Z => n1419);
   U311 : HS65_LH_IVX9 port map( A => n1420, Z => n1418);
   U312 : HS65_LH_IVX9 port map( A => n1411, Z => n1410);
   U313 : HS65_LH_IVX9 port map( A => n1411, Z => n1405);
   U314 : HS65_LH_IVX9 port map( A => n1399, Z => n1397);
   U315 : HS65_LH_IVX9 port map( A => n1399, Z => n1395);
   U316 : HS65_LH_IVX9 port map( A => n352, Z => n334);
   U317 : HS65_LH_IVX9 port map( A => n352, Z => n333);
   U318 : HS65_LH_IVX9 port map( A => n320, Z => n319);
   U319 : HS65_LH_IVX9 port map( A => n320, Z => n318);
   U320 : HS65_LH_IVX9 port map( A => n295, Z => n294);
   U321 : HS65_LH_IVX9 port map( A => n295, Z => n293);
   U322 : HS65_LH_IVX9 port map( A => n330, Z => n329);
   U323 : HS65_LH_IVX9 port map( A => n330, Z => n328);
   U324 : HS65_LH_IVX9 port map( A => n290, Z => n289);
   U325 : HS65_LH_IVX9 port map( A => n290, Z => n288);
   U326 : HS65_LH_BFX9 port map( A => n259, Z => n2500);
   U327 : HS65_LH_BFX9 port map( A => n263, Z => n2495);
   U328 : HS65_LH_BFX9 port map( A => n261, Z => n2490);
   U329 : HS65_LH_BFX9 port map( A => n262, Z => n2485);
   U330 : HS65_LH_BFX9 port map( A => n266, Z => n2465);
   U331 : HS65_LH_BFX9 port map( A => n264, Z => n2460);
   U332 : HS65_LH_BFX9 port map( A => n267, Z => n2455);
   U333 : HS65_LH_BFX9 port map( A => n265, Z => n2450);
   U334 : HS65_LH_IVX9 port map( A => n305, Z => n304);
   U335 : HS65_LH_IVX9 port map( A => n305, Z => n303);
   U336 : HS65_LH_IVX9 port map( A => n315, Z => n314);
   U337 : HS65_LH_IVX9 port map( A => n315, Z => n313);
   U338 : HS65_LH_IVX9 port map( A => n310, Z => n309);
   U339 : HS65_LH_IVX9 port map( A => n310, Z => n308);
   U340 : HS65_LH_BFX9 port map( A => n257, Z => n2509);
   U341 : HS65_LH_BFX9 port map( A => n258, Z => n2504);
   U342 : HS65_LH_BFX9 port map( A => n276, Z => n2429);
   U343 : HS65_LH_BFX9 port map( A => n277, Z => n1432);
   U344 : HS65_LH_BFX9 port map( A => n275, Z => n1421);
   U345 : HS65_LH_BFX9 port map( A => n274, Z => n321);
   U346 : HS65_LH_BFX9 port map( A => n273, Z => n331);
   U347 : HS65_LH_BFX9 port map( A => n272, Z => n291);
   U348 : HS65_LH_BFX9 port map( A => n2435, Z => n2433);
   U349 : HS65_LH_BFX9 port map( A => n327, Z => n325);
   U350 : HS65_LH_IVX9 port map( A => n2432, Z => n2431);
   U351 : HS65_LH_IVX9 port map( A => n324, Z => n323);
   U352 : HS65_LH_BFX9 port map( A => n257, Z => n2510);
   U353 : HS65_LH_BFX9 port map( A => n258, Z => n2505);
   U354 : HS65_LH_BFX9 port map( A => n260, Z => n2480);
   U355 : HS65_LH_BFX9 port map( A => n269, Z => n1413);
   U356 : HS65_LH_BFX9 port map( A => n268, Z => n1403);
   U357 : HS65_LH_BFX9 port map( A => n271, Z => n1392);
   U358 : HS65_LH_BFX9 port map( A => n270, Z => n297);
   U359 : HS65_LH_BFX9 port map( A => n2428, Z => n2430);
   U360 : HS65_LH_BFX9 port map( A => n1427, Z => n1433);
   U361 : HS65_LH_BFX9 port map( A => n1420, Z => n1422);
   U362 : HS65_LH_BFX9 port map( A => n320, Z => n322);
   U363 : HS65_LH_BFX9 port map( A => n273, Z => n332);
   U364 : HS65_LH_BFX9 port map( A => n272, Z => n292);
   U365 : HS65_LH_BFX9 port map( A => n2432, Z => n2434);
   U366 : HS65_LH_BFX9 port map( A => n324, Z => n326);
   U367 : HS65_LH_BFX9 port map( A => n2764, Z => n2762);
   U368 : HS65_LH_BFX9 port map( A => n2764, Z => n2761);
   U369 : HS65_LH_BFX9 port map( A => n2764, Z => n2763);
   U370 : HS65_LH_BFX9 port map( A => n897, Z => n2544);
   U371 : HS65_LH_BFX9 port map( A => n892, Z => n2556);
   U372 : HS65_LH_BFX9 port map( A => n897, Z => n2545);
   U373 : HS65_LH_BFX9 port map( A => n892, Z => n2557);
   U374 : HS65_LH_BFX9 port map( A => n875, Z => n2589);
   U375 : HS65_LH_BFX9 port map( A => n870, Z => n2601);
   U376 : HS65_LH_BFX9 port map( A => n875, Z => n2590);
   U377 : HS65_LH_BFX9 port map( A => n870, Z => n2602);
   U378 : HS65_LH_BFX9 port map( A => n369, Z => n2637);
   U379 : HS65_LH_BFX9 port map( A => n369, Z => n2638);
   U380 : HS65_LH_BFX9 port map( A => n347, Z => n2682);
   U381 : HS65_LH_BFX9 port map( A => n347, Z => n2683);
   U382 : HS65_LH_BFX9 port map( A => n372, Z => n2631);
   U383 : HS65_LH_BFX9 port map( A => n372, Z => n2632);
   U384 : HS65_LH_BFX9 port map( A => n904, Z => n2526);
   U385 : HS65_LH_BFX9 port map( A => n904, Z => n2527);
   U386 : HS65_LH_BFX9 port map( A => n906, Z => n2520);
   U387 : HS65_LH_BFX9 port map( A => n902, Z => n2532);
   U388 : HS65_LH_BFX9 port map( A => n884, Z => n2568);
   U389 : HS65_LH_BFX9 port map( A => n906, Z => n2521);
   U390 : HS65_LH_BFX9 port map( A => n902, Z => n2533);
   U391 : HS65_LH_BFX9 port map( A => n884, Z => n2569);
   U392 : HS65_LH_BFX9 port map( A => n907, Z => n2517);
   U393 : HS65_LH_BFX9 port map( A => n903, Z => n2529);
   U394 : HS65_LH_BFX9 port map( A => n885, Z => n2565);
   U395 : HS65_LH_BFX9 port map( A => n907, Z => n2518);
   U396 : HS65_LH_BFX9 port map( A => n903, Z => n2530);
   U397 : HS65_LH_BFX9 port map( A => n885, Z => n2566);
   U398 : HS65_LH_BFX9 port map( A => n909, Z => n2511);
   U399 : HS65_LH_BFX9 port map( A => n905, Z => n2523);
   U400 : HS65_LH_BFX9 port map( A => n887, Z => n2559);
   U401 : HS65_LH_BFX9 port map( A => n909, Z => n2512);
   U402 : HS65_LH_BFX9 port map( A => n905, Z => n2524);
   U403 : HS65_LH_BFX9 port map( A => n887, Z => n2560);
   U404 : HS65_LH_BFX9 port map( A => n381, Z => n2604);
   U405 : HS65_LH_BFX9 port map( A => n377, Z => n2616);
   U406 : HS65_LH_BFX9 port map( A => n359, Z => n2652);
   U407 : HS65_LH_BFX9 port map( A => n381, Z => n2605);
   U408 : HS65_LH_BFX9 port map( A => n377, Z => n2617);
   U409 : HS65_LH_BFX9 port map( A => n359, Z => n2653);
   U410 : HS65_LH_BFX9 port map( A => n379, Z => n2610);
   U411 : HS65_LH_BFX9 port map( A => n375, Z => n2622);
   U412 : HS65_LH_BFX9 port map( A => n357, Z => n2658);
   U413 : HS65_LH_BFX9 port map( A => n379, Z => n2611);
   U414 : HS65_LH_BFX9 port map( A => n375, Z => n2623);
   U415 : HS65_LH_BFX9 port map( A => n357, Z => n2659);
   U416 : HS65_LH_BFX9 port map( A => n378, Z => n2613);
   U417 : HS65_LH_BFX9 port map( A => n374, Z => n2625);
   U418 : HS65_LH_BFX9 port map( A => n356, Z => n2661);
   U419 : HS65_LH_BFX9 port map( A => n378, Z => n2614);
   U420 : HS65_LH_BFX9 port map( A => n374, Z => n2626);
   U421 : HS65_LH_BFX9 port map( A => n356, Z => n2662);
   U422 : HS65_LH_BFX9 port map( A => n376, Z => n2619);
   U423 : HS65_LH_BFX9 port map( A => n376, Z => n2620);
   U424 : HS65_LH_BFX9 port map( A => n897, Z => n2546);
   U425 : HS65_LH_BFX9 port map( A => n875, Z => n2591);
   U426 : HS65_LH_BFX9 port map( A => n907, Z => n2519);
   U427 : HS65_LH_BFX9 port map( A => n903, Z => n2531);
   U428 : HS65_LH_BFX9 port map( A => n885, Z => n2567);
   U429 : HS65_LH_BFX9 port map( A => n909, Z => n2513);
   U430 : HS65_LH_BFX9 port map( A => n905, Z => n2525);
   U431 : HS65_LH_BFX9 port map( A => n887, Z => n2561);
   U432 : HS65_LH_BFX9 port map( A => n381, Z => n2606);
   U433 : HS65_LH_BFX9 port map( A => n377, Z => n2618);
   U434 : HS65_LH_BFX9 port map( A => n359, Z => n2654);
   U435 : HS65_LH_BFX9 port map( A => n379, Z => n2612);
   U436 : HS65_LH_BFX9 port map( A => n375, Z => n2624);
   U437 : HS65_LH_BFX9 port map( A => n357, Z => n2660);
   U438 : HS65_LH_BFX9 port map( A => n378, Z => n2615);
   U439 : HS65_LH_BFX9 port map( A => n374, Z => n2627);
   U440 : HS65_LH_BFX9 port map( A => n356, Z => n2663);
   U441 : HS65_LH_BFX9 port map( A => n376, Z => n2621);
   U442 : HS65_LH_BFX9 port map( A => n904, Z => n2528);
   U443 : HS65_LH_BFX9 port map( A => n906, Z => n2522);
   U444 : HS65_LH_BFX9 port map( A => n902, Z => n2534);
   U445 : HS65_LH_BFX9 port map( A => n884, Z => n2570);
   U446 : HS65_LH_NAND2X7 port map( A => n842, B => n841, Z => n345);
   U447 : HS65_LH_NAND2X7 port map( A => n1370, B => n1369, Z => n873);
   U448 : HS65_LH_BFX9 port map( A => n882, Z => n2574);
   U449 : HS65_LH_BFX9 port map( A => n883, Z => n2571);
   U450 : HS65_LH_BFX9 port map( A => n881, Z => n2577);
   U451 : HS65_LH_BFX9 port map( A => n882, Z => n2575);
   U452 : HS65_LH_BFX9 port map( A => n883, Z => n2572);
   U453 : HS65_LH_BFX9 port map( A => n881, Z => n2578);
   U454 : HS65_LH_BFX9 port map( A => n373, Z => n2628);
   U455 : HS65_LH_BFX9 port map( A => n368, Z => n2640);
   U456 : HS65_LH_BFX9 port map( A => n373, Z => n2629);
   U457 : HS65_LH_BFX9 port map( A => n368, Z => n2641);
   U458 : HS65_LH_BFX9 port map( A => n346, Z => n2685);
   U459 : HS65_LH_BFX9 port map( A => n346, Z => n2686);
   U460 : HS65_LH_BFX9 port map( A => n354, Z => n2667);
   U461 : HS65_LH_BFX9 port map( A => n355, Z => n2664);
   U462 : HS65_LH_BFX9 port map( A => n353, Z => n2670);
   U463 : HS65_LH_BFX9 port map( A => n354, Z => n2668);
   U464 : HS65_LH_BFX9 port map( A => n355, Z => n2665);
   U465 : HS65_LH_BFX9 port map( A => n353, Z => n2671);
   U466 : HS65_LH_BFX9 port map( A => n351, Z => n2673);
   U467 : HS65_LH_BFX9 port map( A => n351, Z => n2674);
   U468 : HS65_LH_BFX9 port map( A => n898, Z => n2541);
   U469 : HS65_LH_BFX9 port map( A => n898, Z => n2542);
   U470 : HS65_LH_BFX9 port map( A => n876, Z => n2586);
   U471 : HS65_LH_BFX9 port map( A => n871, Z => n2598);
   U472 : HS65_LH_BFX9 port map( A => n876, Z => n2587);
   U473 : HS65_LH_BFX9 port map( A => n871, Z => n2599);
   U474 : HS65_LH_BFX9 port map( A => n364, Z => n2649);
   U475 : HS65_LH_BFX9 port map( A => n364, Z => n2650);
   U476 : HS65_LH_BFX9 port map( A => n342, Z => n2694);
   U477 : HS65_LH_BFX9 port map( A => n342, Z => n2695);
   U478 : HS65_LH_BFX9 port map( A => n901, Z => n2535);
   U479 : HS65_LH_BFX9 port map( A => n896, Z => n2547);
   U480 : HS65_LH_BFX9 port map( A => n901, Z => n2536);
   U481 : HS65_LH_BFX9 port map( A => n896, Z => n2548);
   U482 : HS65_LH_BFX9 port map( A => n367, Z => n2643);
   U483 : HS65_LH_BFX9 port map( A => n367, Z => n2644);
   U484 : HS65_LH_BFX9 port map( A => n874, Z => n2592);
   U485 : HS65_LH_BFX9 port map( A => n874, Z => n2593);
   U486 : HS65_LH_BFX9 port map( A => n370, Z => n2634);
   U487 : HS65_LH_BFX9 port map( A => n370, Z => n2635);
   U488 : HS65_LH_BFX9 port map( A => n348, Z => n2679);
   U489 : HS65_LH_BFX9 port map( A => n343, Z => n2691);
   U490 : HS65_LH_BFX9 port map( A => n348, Z => n2680);
   U491 : HS65_LH_BFX9 port map( A => n343, Z => n2692);
   U492 : HS65_LH_BFX9 port map( A => n879, Z => n2580);
   U493 : HS65_LH_BFX9 port map( A => n879, Z => n2581);
   U494 : HS65_LH_BFX9 port map( A => n350, Z => n2676);
   U495 : HS65_LH_BFX9 port map( A => n350, Z => n2677);
   U496 : HS65_LH_BFX9 port map( A => n900, Z => n2538);
   U497 : HS65_LH_BFX9 port map( A => n895, Z => n2550);
   U498 : HS65_LH_BFX9 port map( A => n900, Z => n2539);
   U499 : HS65_LH_BFX9 port map( A => n895, Z => n2551);
   U500 : HS65_LH_BFX9 port map( A => n878, Z => n2583);
   U501 : HS65_LH_BFX9 port map( A => n878, Z => n2584);
   U502 : HS65_LH_BFX9 port map( A => n354, Z => n2669);
   U503 : HS65_LH_BFX9 port map( A => n355, Z => n2666);
   U504 : HS65_LH_BFX9 port map( A => n353, Z => n2672);
   U505 : HS65_LH_BFX9 port map( A => n369, Z => n2639);
   U506 : HS65_LH_BFX9 port map( A => n364, Z => n2651);
   U507 : HS65_LH_BFX9 port map( A => n347, Z => n2684);
   U508 : HS65_LH_BFX9 port map( A => n342, Z => n2696);
   U509 : HS65_LH_BFX9 port map( A => n372, Z => n2633);
   U510 : HS65_LH_BFX9 port map( A => n367, Z => n2645);
   U511 : HS65_LH_BFX9 port map( A => n350, Z => n2678);
   U512 : HS65_LH_BFX9 port map( A => n878, Z => n2585);
   U513 : HS65_LH_IVX9 port map( A => n2710, Z => n2709);
   U514 : HS65_LH_IVX9 port map( A => n2712, Z => n2711);
   U515 : HS65_LH_IVX9 port map( A => n2714, Z => n2713);
   U516 : HS65_LH_IVX9 port map( A => n2716, Z => n2715);
   U517 : HS65_LH_IVX9 port map( A => n2718, Z => n2717);
   U518 : HS65_LH_IVX9 port map( A => n2720, Z => n2719);
   U519 : HS65_LH_IVX9 port map( A => n2722, Z => n2721);
   U520 : HS65_LH_IVX9 port map( A => n2724, Z => n2723);
   U521 : HS65_LH_IVX9 port map( A => n2726, Z => n2725);
   U522 : HS65_LH_IVX9 port map( A => n2728, Z => n2727);
   U523 : HS65_LH_IVX9 port map( A => n2730, Z => n2729);
   U524 : HS65_LH_IVX9 port map( A => n2732, Z => n2731);
   U525 : HS65_LH_IVX9 port map( A => n2734, Z => n2733);
   U526 : HS65_LH_IVX9 port map( A => n2736, Z => n2735);
   U527 : HS65_LH_IVX9 port map( A => n2738, Z => n2737);
   U528 : HS65_LH_IVX9 port map( A => n2740, Z => n2739);
   U529 : HS65_LH_IVX9 port map( A => n2742, Z => n2741);
   U530 : HS65_LH_IVX9 port map( A => n2744, Z => n2743);
   U531 : HS65_LH_IVX9 port map( A => n2746, Z => n2745);
   U532 : HS65_LH_IVX9 port map( A => n2748, Z => n2747);
   U533 : HS65_LH_IVX9 port map( A => n2750, Z => n2749);
   U534 : HS65_LH_IVX9 port map( A => n2752, Z => n2751);
   U535 : HS65_LH_IVX9 port map( A => n2754, Z => n2753);
   U536 : HS65_LH_IVX9 port map( A => n2756, Z => n2755);
   U537 : HS65_LH_IVX9 port map( A => n2758, Z => n2757);
   U538 : HS65_LH_IVX9 port map( A => n2760, Z => n2759);
   U539 : HS65_LH_BFX9 port map( A => n900, Z => n2540);
   U540 : HS65_LH_BFX9 port map( A => n895, Z => n2552);
   U541 : HS65_LH_BFX9 port map( A => n882, Z => n2576);
   U542 : HS65_LH_BFX9 port map( A => n883, Z => n2573);
   U543 : HS65_LH_BFX9 port map( A => n881, Z => n2579);
   U544 : HS65_LH_IVX9 port map( A => n2698, Z => n2697);
   U545 : HS65_LH_IVX9 port map( A => n2700, Z => n2699);
   U546 : HS65_LH_IVX9 port map( A => n2702, Z => n2701);
   U547 : HS65_LH_IVX9 port map( A => n2704, Z => n2703);
   U548 : HS65_LH_IVX9 port map( A => n2706, Z => n2705);
   U549 : HS65_LH_IVX9 port map( A => n2708, Z => n2707);
   U550 : HS65_LH_BFX9 port map( A => n892, Z => n2558);
   U551 : HS65_LH_BFX9 port map( A => n870, Z => n2603);
   U552 : HS65_LH_BFX9 port map( A => n346, Z => n2687);
   U553 : HS65_LH_BFX9 port map( A => n351, Z => n2675);
   U554 : HS65_LH_BFX9 port map( A => n373, Z => n2630);
   U555 : HS65_LH_BFX9 port map( A => n368, Z => n2642);
   U556 : HS65_LH_BFX9 port map( A => n874, Z => n2594);
   U557 : HS65_LH_BFX9 port map( A => n879, Z => n2582);
   U558 : HS65_LH_BFX9 port map( A => n901, Z => n2537);
   U559 : HS65_LH_BFX9 port map( A => n896, Z => n2549);
   U560 : HS65_LH_BFX9 port map( A => n898, Z => n2543);
   U561 : HS65_LH_BFX9 port map( A => n876, Z => n2588);
   U562 : HS65_LH_BFX9 port map( A => n871, Z => n2600);
   U563 : HS65_LH_BFX9 port map( A => n370, Z => n2636);
   U564 : HS65_LH_BFX9 port map( A => n348, Z => n2681);
   U565 : HS65_LH_BFX9 port map( A => n343, Z => n2693);
   U566 : HS65_LH_BFX9 port map( A => n257, Z => n2508);
   U567 : HS65_LH_BFX9 port map( A => n258, Z => n2503);
   U568 : HS65_LH_BFX9 port map( A => n261, Z => n2488);
   U569 : HS65_LH_BFX9 port map( A => n262, Z => n2483);
   U570 : HS65_LH_BFX9 port map( A => n1407, Z => n2473);
   U571 : HS65_LH_BFX9 port map( A => n1409, Z => n2468);
   U572 : HS65_LH_BFX9 port map( A => n1414, Z => n2443);
   U573 : HS65_LH_BFX9 port map( A => n1415, Z => n2438);
   U574 : HS65_LH_BFX9 port map( A => n1431, Z => n300);
   U575 : HS65_LH_BFX9 port map( A => n259, Z => n2498);
   U576 : HS65_LH_BFX9 port map( A => n263, Z => n2493);
   U577 : HS65_LH_BFX9 port map( A => n260, Z => n2478);
   U578 : HS65_LH_BFX9 port map( A => n266, Z => n2463);
   U579 : HS65_LH_BFX9 port map( A => n264, Z => n2458);
   U580 : HS65_LH_BFX9 port map( A => n267, Z => n2453);
   U581 : HS65_LH_BFX9 port map( A => n265, Z => n2448);
   U582 : HS65_LH_BFX9 port map( A => n269, Z => n1411);
   U583 : HS65_LH_BFX9 port map( A => n268, Z => n1399);
   U584 : HS65_LH_BFX9 port map( A => n271, Z => n352);
   U585 : HS65_LH_BFX9 port map( A => n270, Z => n295);
   U586 : HS65_LH_BFX9 port map( A => n276, Z => n2428);
   U587 : HS65_LH_BFX9 port map( A => n277, Z => n1427);
   U588 : HS65_LH_BFX9 port map( A => n275, Z => n1420);
   U589 : HS65_LH_BFX9 port map( A => n274, Z => n320);
   U590 : HS65_LH_BFX9 port map( A => n273, Z => n330);
   U591 : HS65_LH_BFX9 port map( A => n272, Z => n290);
   U592 : HS65_LH_BFX9 port map( A => n1428, Z => n315);
   U593 : HS65_LH_BFX9 port map( A => n1429, Z => n310);
   U594 : HS65_LH_BFX9 port map( A => n1430, Z => n305);
   U595 : HS65_LH_BFX9 port map( A => n1407, Z => n2474);
   U596 : HS65_LH_BFX9 port map( A => n1409, Z => n2469);
   U597 : HS65_LH_BFX9 port map( A => n1414, Z => n2444);
   U598 : HS65_LH_BFX9 port map( A => n1415, Z => n2439);
   U599 : HS65_LH_BFX9 port map( A => n1428, Z => n316);
   U600 : HS65_LH_BFX9 port map( A => n1429, Z => n311);
   U601 : HS65_LH_BFX9 port map( A => n1430, Z => n306);
   U602 : HS65_LH_BFX9 port map( A => n1431, Z => n301);
   U603 : HS65_LH_BFX9 port map( A => n2435, Z => n2432);
   U604 : HS65_LH_IVX9 port map( A => n1416, Z => n2435);
   U605 : HS65_LH_BFX9 port map( A => n327, Z => n324);
   U606 : HS65_LH_IVX9 port map( A => n1425, Z => n327);
   U607 : HS65_LH_BFX9 port map( A => n1407, Z => n2475);
   U608 : HS65_LH_BFX9 port map( A => n1409, Z => n2470);
   U609 : HS65_LH_BFX9 port map( A => n1414, Z => n2445);
   U610 : HS65_LH_BFX9 port map( A => n1415, Z => n2440);
   U611 : HS65_LH_BFX9 port map( A => n1428, Z => n317);
   U612 : HS65_LH_BFX9 port map( A => n1429, Z => n312);
   U613 : HS65_LH_BFX9 port map( A => n1430, Z => n307);
   U614 : HS65_LH_BFX9 port map( A => n1431, Z => n302);
   U615 : HS65_LH_BFX9 port map( A => rst_n, Z => n2764);
   U616 : HS65_LH_NAND2X7 port map( A => n846, B => n857, Z => n372);
   U617 : HS65_LH_NOR2X6 port map( A => n2900, B => n2899, Z => n841);
   U618 : HS65_LH_NOR2X6 port map( A => n2905, B => n2904, Z => n1369);
   U619 : HS65_LH_AND2X4 port map( A => n859, B => n2898, Z => n857);
   U620 : HS65_LH_AND2X4 port map( A => n862, B => n2898, Z => n861);
   U621 : HS65_LH_AND2X4 port map( A => n1390, B => n2903, Z => n1389);
   U622 : HS65_LH_NOR2X6 port map( A => n2902, B => n2901, Z => n859);
   U623 : HS65_LH_NOR2X6 port map( A => n2907, B => n2906, Z => n1387);
   U624 : HS65_LH_AND2X4 port map( A => n850, B => n2898, Z => n849);
   U625 : HS65_LH_AND2X4 port map( A => n1378, B => n2903, Z => n1377);
   U626 : HS65_LH_BFX9 port map( A => n2893, Z => n280);
   U627 : HS65_LH_BFX9 port map( A => n2894, Z => n285);
   U628 : HS65_LH_BFX9 port map( A => n2893, Z => n278);
   U629 : HS65_LH_BFX9 port map( A => n2893, Z => n279);
   U630 : HS65_LH_BFX9 port map( A => n2894, Z => n283);
   U631 : HS65_LH_BFX9 port map( A => n2894, Z => n284);
   U632 : HS65_LH_NAND2X7 port map( A => n840, B => n841, Z => n346);
   U633 : HS65_LH_NAND2X7 port map( A => n1368, B => n1369, Z => n874);
   U634 : HS65_LH_NAND2X7 port map( A => n842, B => n845, Z => n350);
   U635 : HS65_LH_NAND2X7 port map( A => n840, B => n845, Z => n351);
   U636 : HS65_LH_NAND2X7 port map( A => n1370, B => n1373, Z => n878);
   U637 : HS65_LH_NAND2X7 port map( A => n1368, B => n1373, Z => n879);
   U638 : HS65_LH_NAND2X7 port map( A => n843, B => n857, Z => n367);
   U639 : HS65_LH_NAND2X7 port map( A => n843, B => n856, Z => n368);
   U640 : HS65_LH_NAND2X7 port map( A => n1371, B => n1385, Z => n895);
   U641 : HS65_LH_NAND2X7 port map( A => n1371, B => n1384, Z => n896);
   U642 : HS65_LH_NAND2X7 port map( A => n846, B => n856, Z => n373);
   U643 : HS65_LH_NAND2X7 port map( A => n1374, B => n1385, Z => n900);
   U644 : HS65_LH_NAND2X7 port map( A => n1374, B => n1384, Z => n901);
   U645 : HS65_LH_AND2X4 port map( A => n847, B => n2898, Z => n842);
   U646 : HS65_LH_AND2X4 port map( A => n1375, B => n2903, Z => n1370);
   U647 : HS65_LH_AND2X4 port map( A => n1387, B => n2903, Z => n1385);
   U648 : HS65_LH_BFX9 port map( A => n2893, Z => n281);
   U649 : HS65_LH_BFX9 port map( A => n2894, Z => n287);
   U650 : HS65_LH_BFX9 port map( A => n2894, Z => n286);
   U651 : HS65_LH_BFX9 port map( A => n2893, Z => n282);
   U652 : HS65_LH_NAND2X7 port map( A => n1408, B => n1391, Z => n1407);
   U653 : HS65_LH_NAND2X7 port map( A => n1408, B => n1393, Z => n1409);
   U654 : HS65_LH_NAND2X7 port map( A => n1408, B => n1404, Z => n1414);
   U655 : HS65_LH_NAND2X7 port map( A => n1408, B => n1406, Z => n1415);
   U656 : HS65_LH_NAND2X7 port map( A => n1426, B => n1402, Z => n1431);
   U657 : HS65_LH_NAND2X7 port map( A => n1417, B => n1391, Z => n1416);
   U658 : HS65_LH_NAND2X7 port map( A => n1426, B => n1391, Z => n1425);
   U659 : HS65_LH_NAND2X7 port map( A => n1426, B => n1400, Z => n1430);
   U660 : HS65_LH_NAND2X7 port map( A => n1426, B => n1396, Z => n1428);
   U661 : HS65_LH_NAND2X7 port map( A => n1426, B => n1398, Z => n1429);
   U662 : HS65_LH_IVX9 port map( A => regfile_i(1), Z => n2894);
   U663 : HS65_LH_NOR2X6 port map( A => n2900, B => regfile_i(41), Z => n843);
   U664 : HS65_LH_NOR2X6 port map( A => n2905, B => regfile_i(46), Z => n1371);
   U665 : HS65_LH_NOR2X6 port map( A => n2899, B => regfile_i(42), Z => n846);
   U666 : HS65_LH_NOR2X6 port map( A => n2904, B => regfile_i(47), Z => n1374);
   U667 : HS65_LH_NOR2X6 port map( A => regfile_i(41), B => regfile_i(42), Z =>
                           n845);
   U668 : HS65_LH_NOR2X6 port map( A => regfile_i(46), B => regfile_i(47), Z =>
                           n1373);
   U669 : HS65_LH_AOI212X4 port map( A => registers_11_0_port, B => n2682, C =>
                           registers_10_0_port, D => n2679, E => n844, Z => 
                           n837);
   U670 : HS65_LH_OAI22X6 port map( A => n2676, B => n256, C => n2673, D => 
                           n224, Z => n844);
   U671 : HS65_LH_AOI212X4 port map( A => registers_11_1_port, B => n2682, C =>
                           registers_10_1_port, D => n2679, E => n675, Z => 
                           n672);
   U672 : HS65_LH_OAI22X6 port map( A => n2676, B => n255, C => n2673, D => 
                           n223, Z => n675);
   U673 : HS65_LH_AOI212X4 port map( A => registers_11_2_port, B => n2683, C =>
                           registers_10_2_port, D => n2680, E => n510, Z => 
                           n507);
   U674 : HS65_LH_OAI22X6 port map( A => n2677, B => n254, C => n2674, D => 
                           n222, Z => n510);
   U675 : HS65_LH_AOI212X4 port map( A => registers_11_11_port, B => n2682, C 
                           => registers_10_11_port, D => n2679, E => n810, Z =>
                           n807);
   U676 : HS65_LH_OAI22X6 port map( A => n2676, B => n245, C => n2673, D => 
                           n213, Z => n810);
   U677 : HS65_LH_AOI212X4 port map( A => registers_11_12_port, B => n2682, C 
                           => registers_10_12_port, D => n2679, E => n795, Z =>
                           n792);
   U678 : HS65_LH_OAI22X6 port map( A => n2676, B => n244, C => n2673, D => 
                           n212, Z => n795);
   U679 : HS65_LH_AOI212X4 port map( A => registers_11_13_port, B => n2682, C 
                           => registers_10_13_port, D => n2679, E => n780, Z =>
                           n777);
   U680 : HS65_LH_OAI22X6 port map( A => n2676, B => n243, C => n2673, D => 
                           n211, Z => n780);
   U681 : HS65_LH_AOI212X4 port map( A => registers_11_14_port, B => n2682, C 
                           => registers_10_14_port, D => n2679, E => n765, Z =>
                           n762);
   U682 : HS65_LH_OAI22X6 port map( A => n2676, B => n242, C => n2673, D => 
                           n210, Z => n765);
   U683 : HS65_LH_AOI212X4 port map( A => registers_11_15_port, B => n2682, C 
                           => registers_10_15_port, D => n2679, E => n750, Z =>
                           n747);
   U684 : HS65_LH_OAI22X6 port map( A => n2676, B => n241, C => n2673, D => 
                           n209, Z => n750);
   U685 : HS65_LH_AOI212X4 port map( A => registers_11_16_port, B => n2682, C 
                           => registers_10_16_port, D => n2679, E => n735, Z =>
                           n732);
   U686 : HS65_LH_OAI22X6 port map( A => n2676, B => n240, C => n2673, D => 
                           n208, Z => n735);
   U687 : HS65_LH_AOI212X4 port map( A => registers_11_17_port, B => n2682, C 
                           => registers_10_17_port, D => n2679, E => n720, Z =>
                           n717);
   U688 : HS65_LH_OAI22X6 port map( A => n2676, B => n239, C => n2673, D => 
                           n207, Z => n720);
   U689 : HS65_LH_AOI212X4 port map( A => registers_11_18_port, B => n2682, C 
                           => registers_10_18_port, D => n2679, E => n705, Z =>
                           n702);
   U690 : HS65_LH_OAI22X6 port map( A => n2676, B => n238, C => n2673, D => 
                           n206, Z => n705);
   U691 : HS65_LH_AOI212X4 port map( A => registers_11_19_port, B => n2682, C 
                           => registers_10_19_port, D => n2679, E => n690, Z =>
                           n687);
   U692 : HS65_LH_OAI22X6 port map( A => n2676, B => n237, C => n2673, D => 
                           n205, Z => n690);
   U693 : HS65_LH_AOI212X4 port map( A => registers_11_20_port, B => n2683, C 
                           => registers_10_20_port, D => n2679, E => n660, Z =>
                           n657);
   U694 : HS65_LH_OAI22X6 port map( A => n2677, B => n236, C => n2673, D => 
                           n204, Z => n660);
   U695 : HS65_LH_AOI212X4 port map( A => registers_11_21_port, B => n2683, C 
                           => registers_10_21_port, D => n2680, E => n645, Z =>
                           n642);
   U696 : HS65_LH_OAI22X6 port map( A => n2677, B => n235, C => n2674, D => 
                           n203, Z => n645);
   U697 : HS65_LH_AOI212X4 port map( A => registers_11_22_port, B => n2683, C 
                           => registers_10_22_port, D => n2680, E => n630, Z =>
                           n627);
   U698 : HS65_LH_OAI22X6 port map( A => n2677, B => n234, C => n2674, D => 
                           n202, Z => n630);
   U699 : HS65_LH_AOI212X4 port map( A => registers_11_23_port, B => n2683, C 
                           => registers_10_23_port, D => n2680, E => n615, Z =>
                           n612);
   U700 : HS65_LH_OAI22X6 port map( A => n2677, B => n233, C => n2674, D => 
                           n201, Z => n615);
   U701 : HS65_LH_AOI212X4 port map( A => registers_11_24_port, B => n2683, C 
                           => registers_10_24_port, D => n2680, E => n600, Z =>
                           n597);
   U702 : HS65_LH_OAI22X6 port map( A => n2677, B => n232, C => n2674, D => 
                           n200, Z => n600);
   U703 : HS65_LH_AOI212X4 port map( A => registers_11_25_port, B => n2683, C 
                           => registers_10_25_port, D => n2680, E => n585, Z =>
                           n582);
   U704 : HS65_LH_OAI22X6 port map( A => n2677, B => n231, C => n2674, D => 
                           n199, Z => n585);
   U705 : HS65_LH_AOI212X4 port map( A => registers_11_26_port, B => n2683, C 
                           => registers_10_26_port, D => n2680, E => n570, Z =>
                           n567);
   U706 : HS65_LH_OAI22X6 port map( A => n2677, B => n230, C => n2674, D => 
                           n198, Z => n570);
   U707 : HS65_LH_AOI212X4 port map( A => registers_11_27_port, B => n2683, C 
                           => registers_10_27_port, D => n2680, E => n555, Z =>
                           n552);
   U708 : HS65_LH_OAI22X6 port map( A => n2677, B => n229, C => n2674, D => 
                           n197, Z => n555);
   U709 : HS65_LH_AOI212X4 port map( A => registers_11_28_port, B => n2683, C 
                           => registers_10_28_port, D => n2680, E => n540, Z =>
                           n537);
   U710 : HS65_LH_OAI22X6 port map( A => n2677, B => n228, C => n2674, D => 
                           n196, Z => n540);
   U711 : HS65_LH_AOI212X4 port map( A => registers_11_29_port, B => n2683, C 
                           => registers_10_29_port, D => n2680, E => n525, Z =>
                           n522);
   U712 : HS65_LH_OAI22X6 port map( A => n2677, B => n227, C => n2674, D => 
                           n195, Z => n525);
   U713 : HS65_LH_AOI212X4 port map( A => registers_11_30_port, B => n2683, C 
                           => registers_10_30_port, D => n2680, E => n495, Z =>
                           n492);
   U714 : HS65_LH_OAI22X6 port map( A => n2677, B => n226, C => n2674, D => 
                           n194, Z => n495);
   U715 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_0_port, C =>
                           n2586, D => registers_10_0_port, E => n1372, Z => 
                           n1365);
   U716 : HS65_LH_OAI22X6 port map( A => n256, B => n2583, C => n224, D => 
                           n2580, Z => n1372);
   U717 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_1_port, C =>
                           n2586, D => registers_10_1_port, E => n1203, Z => 
                           n1200);
   U718 : HS65_LH_OAI22X6 port map( A => n255, B => n2583, C => n223, D => 
                           n2580, Z => n1203);
   U719 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_2_port, C =>
                           n2587, D => registers_10_2_port, E => n1038, Z => 
                           n1035);
   U720 : HS65_LH_OAI22X6 port map( A => n254, B => n2584, C => n222, D => 
                           n2581, Z => n1038);
   U721 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_3_port, C =>
                           n2587, D => registers_10_3_port, E => n993, Z => 
                           n990);
   U722 : HS65_LH_OAI22X6 port map( A => n253, B => n2585, C => n221, D => 
                           n2581, Z => n993);
   U723 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_4_port, C =>
                           n2588, D => registers_10_4_port, E => n978, Z => 
                           n975);
   U724 : HS65_LH_OAI22X6 port map( A => n252, B => n2585, C => n220, D => 
                           n2582, Z => n978);
   U725 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_5_port, C =>
                           n2588, D => registers_10_5_port, E => n963, Z => 
                           n960);
   U726 : HS65_LH_OAI22X6 port map( A => n251, B => n2585, C => n219, D => 
                           n2582, Z => n963);
   U727 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_6_port, C =>
                           n2588, D => registers_10_6_port, E => n948, Z => 
                           n945);
   U728 : HS65_LH_OAI22X6 port map( A => n250, B => n2585, C => n218, D => 
                           n2582, Z => n948);
   U729 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_7_port, C =>
                           n2588, D => registers_10_7_port, E => n933, Z => 
                           n930);
   U730 : HS65_LH_OAI22X6 port map( A => n249, B => n2585, C => n217, D => 
                           n2582, Z => n933);
   U731 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_8_port, C =>
                           n2588, D => registers_10_8_port, E => n918, Z => 
                           n915);
   U732 : HS65_LH_OAI22X6 port map( A => n248, B => n2585, C => n216, D => 
                           n2582, Z => n918);
   U733 : HS65_LH_AOI212X4 port map( A => n2591, B => registers_11_9_port, C =>
                           n2588, D => registers_10_9_port, E => n877, Z => 
                           n868);
   U734 : HS65_LH_OAI22X6 port map( A => n247, B => n2585, C => n215, D => 
                           n2582, Z => n877);
   U735 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_10_port, C 
                           => n2586, D => registers_10_10_port, E => n1353, Z 
                           => n1350);
   U736 : HS65_LH_OAI22X6 port map( A => n246, B => n2583, C => n214, D => 
                           n2580, Z => n1353);
   U737 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_11_port, C 
                           => n2586, D => registers_10_11_port, E => n1338, Z 
                           => n1335);
   U738 : HS65_LH_OAI22X6 port map( A => n245, B => n2583, C => n213, D => 
                           n2580, Z => n1338);
   U739 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_12_port, C 
                           => n2586, D => registers_10_12_port, E => n1323, Z 
                           => n1320);
   U740 : HS65_LH_OAI22X6 port map( A => n244, B => n2583, C => n212, D => 
                           n2580, Z => n1323);
   U741 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_13_port, C 
                           => n2586, D => registers_10_13_port, E => n1308, Z 
                           => n1305);
   U742 : HS65_LH_OAI22X6 port map( A => n243, B => n2583, C => n211, D => 
                           n2580, Z => n1308);
   U743 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_14_port, C 
                           => n2586, D => registers_10_14_port, E => n1293, Z 
                           => n1290);
   U744 : HS65_LH_OAI22X6 port map( A => n242, B => n2583, C => n210, D => 
                           n2580, Z => n1293);
   U745 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_15_port, C 
                           => n2586, D => registers_10_15_port, E => n1278, Z 
                           => n1275);
   U746 : HS65_LH_OAI22X6 port map( A => n241, B => n2583, C => n209, D => 
                           n2580, Z => n1278);
   U747 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_16_port, C 
                           => n2586, D => registers_10_16_port, E => n1263, Z 
                           => n1260);
   U748 : HS65_LH_OAI22X6 port map( A => n240, B => n2583, C => n208, D => 
                           n2580, Z => n1263);
   U749 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_17_port, C 
                           => n2586, D => registers_10_17_port, E => n1248, Z 
                           => n1245);
   U750 : HS65_LH_OAI22X6 port map( A => n239, B => n2583, C => n207, D => 
                           n2580, Z => n1248);
   U751 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_18_port, C 
                           => n2586, D => registers_10_18_port, E => n1233, Z 
                           => n1230);
   U752 : HS65_LH_OAI22X6 port map( A => n238, B => n2583, C => n206, D => 
                           n2580, Z => n1233);
   U753 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_19_port, C 
                           => n2586, D => registers_10_19_port, E => n1218, Z 
                           => n1215);
   U754 : HS65_LH_OAI22X6 port map( A => n237, B => n2583, C => n205, D => 
                           n2580, Z => n1218);
   U755 : HS65_LH_AOI212X4 port map( A => n2589, B => registers_11_20_port, C 
                           => n2586, D => registers_10_20_port, E => n1188, Z 
                           => n1185);
   U756 : HS65_LH_OAI22X6 port map( A => n236, B => n2584, C => n204, D => 
                           n2580, Z => n1188);
   U757 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_21_port, C 
                           => n2587, D => registers_10_21_port, E => n1173, Z 
                           => n1170);
   U758 : HS65_LH_OAI22X6 port map( A => n235, B => n2584, C => n203, D => 
                           n2581, Z => n1173);
   U759 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_22_port, C 
                           => n2587, D => registers_10_22_port, E => n1158, Z 
                           => n1155);
   U760 : HS65_LH_OAI22X6 port map( A => n234, B => n2584, C => n202, D => 
                           n2581, Z => n1158);
   U761 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_23_port, C 
                           => n2587, D => registers_10_23_port, E => n1143, Z 
                           => n1140);
   U762 : HS65_LH_OAI22X6 port map( A => n233, B => n2584, C => n201, D => 
                           n2581, Z => n1143);
   U763 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_24_port, C 
                           => n2587, D => registers_10_24_port, E => n1128, Z 
                           => n1125);
   U764 : HS65_LH_OAI22X6 port map( A => n232, B => n2584, C => n200, D => 
                           n2581, Z => n1128);
   U765 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_25_port, C 
                           => n2587, D => registers_10_25_port, E => n1113, Z 
                           => n1110);
   U766 : HS65_LH_OAI22X6 port map( A => n231, B => n2584, C => n199, D => 
                           n2581, Z => n1113);
   U767 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_26_port, C 
                           => n2587, D => registers_10_26_port, E => n1098, Z 
                           => n1095);
   U768 : HS65_LH_OAI22X6 port map( A => n230, B => n2584, C => n198, D => 
                           n2581, Z => n1098);
   U769 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_27_port, C 
                           => n2587, D => registers_10_27_port, E => n1083, Z 
                           => n1080);
   U770 : HS65_LH_OAI22X6 port map( A => n229, B => n2584, C => n197, D => 
                           n2581, Z => n1083);
   U771 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_28_port, C 
                           => n2587, D => registers_10_28_port, E => n1068, Z 
                           => n1065);
   U772 : HS65_LH_OAI22X6 port map( A => n228, B => n2584, C => n196, D => 
                           n2581, Z => n1068);
   U773 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_29_port, C 
                           => n2587, D => registers_10_29_port, E => n1053, Z 
                           => n1050);
   U774 : HS65_LH_OAI22X6 port map( A => n227, B => n2584, C => n195, D => 
                           n2581, Z => n1053);
   U775 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_30_port, C 
                           => n2587, D => registers_10_30_port, E => n1023, Z 
                           => n1020);
   U776 : HS65_LH_OAI22X6 port map( A => n226, B => n2584, C => n194, D => 
                           n2581, Z => n1023);
   U777 : HS65_LH_AOI212X4 port map( A => n2590, B => registers_11_31_port, C 
                           => n2587, D => registers_10_31_port, E => n1008, Z 
                           => n1005);
   U778 : HS65_LH_OAI22X6 port map( A => n225, B => n2585, C => n193, D => 
                           n2581, Z => n1008);
   U779 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_0_port, C =>
                           n2598, D => registers_12_0_port, E => n1367, Z => 
                           n1366);
   U780 : HS65_LH_OAI22X6 port map( A => n192, B => n2595, C => n160, D => 
                           n2592, Z => n1367);
   U781 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_1_port, C =>
                           n2598, D => registers_12_1_port, E => n1202, Z => 
                           n1201);
   U782 : HS65_LH_OAI22X6 port map( A => n191, B => n2595, C => n159, D => 
                           n2592, Z => n1202);
   U783 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_2_port, C =>
                           n2599, D => registers_12_2_port, E => n1037, Z => 
                           n1036);
   U784 : HS65_LH_OAI22X6 port map( A => n190, B => n2596, C => n158, D => 
                           n2593, Z => n1037);
   U785 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_3_port, C =>
                           n2599, D => registers_12_3_port, E => n992, Z => 
                           n991);
   U786 : HS65_LH_OAI22X6 port map( A => n189, B => n2597, C => n157, D => 
                           n2593, Z => n992);
   U787 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_10_port, C 
                           => n2598, D => registers_12_10_port, E => n1352, Z 
                           => n1351);
   U788 : HS65_LH_OAI22X6 port map( A => n182, B => n2595, C => n150, D => 
                           n2592, Z => n1352);
   U789 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_11_port, C 
                           => n2598, D => registers_12_11_port, E => n1337, Z 
                           => n1336);
   U790 : HS65_LH_OAI22X6 port map( A => n181, B => n2595, C => n149, D => 
                           n2592, Z => n1337);
   U791 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_12_port, C 
                           => n2598, D => registers_12_12_port, E => n1322, Z 
                           => n1321);
   U792 : HS65_LH_OAI22X6 port map( A => n180, B => n2595, C => n148, D => 
                           n2592, Z => n1322);
   U793 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_13_port, C 
                           => n2598, D => registers_12_13_port, E => n1307, Z 
                           => n1306);
   U794 : HS65_LH_OAI22X6 port map( A => n179, B => n2595, C => n147, D => 
                           n2592, Z => n1307);
   U795 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_14_port, C 
                           => n2598, D => registers_12_14_port, E => n1292, Z 
                           => n1291);
   U796 : HS65_LH_OAI22X6 port map( A => n178, B => n2595, C => n146, D => 
                           n2592, Z => n1292);
   U797 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_15_port, C 
                           => n2598, D => registers_12_15_port, E => n1277, Z 
                           => n1276);
   U798 : HS65_LH_OAI22X6 port map( A => n177, B => n2595, C => n145, D => 
                           n2592, Z => n1277);
   U799 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_16_port, C 
                           => n2598, D => registers_12_16_port, E => n1262, Z 
                           => n1261);
   U800 : HS65_LH_OAI22X6 port map( A => n176, B => n2595, C => n144, D => 
                           n2592, Z => n1262);
   U801 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_17_port, C 
                           => n2598, D => registers_12_17_port, E => n1247, Z 
                           => n1246);
   U802 : HS65_LH_OAI22X6 port map( A => n175, B => n2595, C => n143, D => 
                           n2592, Z => n1247);
   U803 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_18_port, C 
                           => n2598, D => registers_12_18_port, E => n1232, Z 
                           => n1231);
   U804 : HS65_LH_OAI22X6 port map( A => n174, B => n2595, C => n142, D => 
                           n2592, Z => n1232);
   U805 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_19_port, C 
                           => n2598, D => registers_12_19_port, E => n1217, Z 
                           => n1216);
   U806 : HS65_LH_OAI22X6 port map( A => n173, B => n2595, C => n141, D => 
                           n2592, Z => n1217);
   U807 : HS65_LH_AOI212X4 port map( A => n2601, B => registers_13_20_port, C 
                           => n2598, D => registers_12_20_port, E => n1187, Z 
                           => n1186);
   U808 : HS65_LH_OAI22X6 port map( A => n172, B => n2596, C => n140, D => 
                           n2592, Z => n1187);
   U809 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_21_port, C 
                           => n2599, D => registers_12_21_port, E => n1172, Z 
                           => n1171);
   U810 : HS65_LH_OAI22X6 port map( A => n171, B => n2596, C => n139, D => 
                           n2593, Z => n1172);
   U811 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_22_port, C 
                           => n2599, D => registers_12_22_port, E => n1157, Z 
                           => n1156);
   U812 : HS65_LH_OAI22X6 port map( A => n170, B => n2596, C => n138, D => 
                           n2593, Z => n1157);
   U813 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_23_port, C 
                           => n2599, D => registers_12_23_port, E => n1142, Z 
                           => n1141);
   U814 : HS65_LH_OAI22X6 port map( A => n169, B => n2596, C => n137, D => 
                           n2593, Z => n1142);
   U815 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_24_port, C 
                           => n2599, D => registers_12_24_port, E => n1127, Z 
                           => n1126);
   U816 : HS65_LH_OAI22X6 port map( A => n168, B => n2596, C => n136, D => 
                           n2593, Z => n1127);
   U817 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_25_port, C 
                           => n2599, D => registers_12_25_port, E => n1112, Z 
                           => n1111);
   U818 : HS65_LH_OAI22X6 port map( A => n167, B => n2596, C => n135, D => 
                           n2593, Z => n1112);
   U819 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_26_port, C 
                           => n2599, D => registers_12_26_port, E => n1097, Z 
                           => n1096);
   U820 : HS65_LH_OAI22X6 port map( A => n166, B => n2596, C => n134, D => 
                           n2593, Z => n1097);
   U821 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_27_port, C 
                           => n2599, D => registers_12_27_port, E => n1082, Z 
                           => n1081);
   U822 : HS65_LH_OAI22X6 port map( A => n165, B => n2596, C => n133, D => 
                           n2593, Z => n1082);
   U823 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_28_port, C 
                           => n2599, D => registers_12_28_port, E => n1067, Z 
                           => n1066);
   U824 : HS65_LH_OAI22X6 port map( A => n164, B => n2596, C => n132, D => 
                           n2593, Z => n1067);
   U825 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_29_port, C 
                           => n2599, D => registers_12_29_port, E => n1052, Z 
                           => n1051);
   U826 : HS65_LH_OAI22X6 port map( A => n163, B => n2596, C => n131, D => 
                           n2593, Z => n1052);
   U827 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_30_port, C 
                           => n2599, D => registers_12_30_port, E => n1022, Z 
                           => n1021);
   U828 : HS65_LH_OAI22X6 port map( A => n162, B => n2596, C => n130, D => 
                           n2593, Z => n1022);
   U829 : HS65_LH_AOI212X4 port map( A => n2602, B => registers_13_31_port, C 
                           => n2599, D => registers_12_31_port, E => n1007, Z 
                           => n1006);
   U830 : HS65_LH_OAI22X6 port map( A => n161, B => n2597, C => n129, D => 
                           n2593, Z => n1007);
   U831 : HS65_LH_OAI22X6 port map( A => n2631, B => n128, C => n2628, D => n96
                           , Z => n858);
   U832 : HS65_LH_OAI22X6 port map( A => n2631, B => n127, C => n2628, D => n95
                           , Z => n681);
   U833 : HS65_LH_OAI22X6 port map( A => n2632, B => n126, C => n2629, D => n94
                           , Z => n516);
   U834 : HS65_LH_OAI22X6 port map( A => n2631, B => n118, C => n2628, D => n86
                           , Z => n831);
   U835 : HS65_LH_OAI22X6 port map( A => n2631, B => n117, C => n2628, D => n85
                           , Z => n816);
   U836 : HS65_LH_OAI22X6 port map( A => n2631, B => n116, C => n2628, D => n84
                           , Z => n801);
   U837 : HS65_LH_OAI22X6 port map( A => n2631, B => n115, C => n2628, D => n83
                           , Z => n786);
   U838 : HS65_LH_OAI22X6 port map( A => n2631, B => n114, C => n2628, D => n82
                           , Z => n771);
   U839 : HS65_LH_OAI22X6 port map( A => n2631, B => n113, C => n2628, D => n81
                           , Z => n756);
   U840 : HS65_LH_OAI22X6 port map( A => n2631, B => n112, C => n2628, D => n80
                           , Z => n741);
   U841 : HS65_LH_OAI22X6 port map( A => n2631, B => n111, C => n2628, D => n79
                           , Z => n726);
   U842 : HS65_LH_OAI22X6 port map( A => n2631, B => n110, C => n2628, D => n78
                           , Z => n711);
   U843 : HS65_LH_OAI22X6 port map( A => n2631, B => n109, C => n2628, D => n77
                           , Z => n696);
   U844 : HS65_LH_OAI22X6 port map( A => n2632, B => n108, C => n2628, D => n76
                           , Z => n666);
   U845 : HS65_LH_OAI22X6 port map( A => n2632, B => n107, C => n2629, D => n75
                           , Z => n651);
   U846 : HS65_LH_OAI22X6 port map( A => n2632, B => n106, C => n2629, D => n74
                           , Z => n636);
   U847 : HS65_LH_OAI22X6 port map( A => n2632, B => n105, C => n2629, D => n73
                           , Z => n621);
   U848 : HS65_LH_OAI22X6 port map( A => n2632, B => n104, C => n2629, D => n72
                           , Z => n606);
   U849 : HS65_LH_OAI22X6 port map( A => n2632, B => n103, C => n2629, D => n71
                           , Z => n591);
   U850 : HS65_LH_OAI22X6 port map( A => n2632, B => n102, C => n2629, D => n70
                           , Z => n576);
   U851 : HS65_LH_OAI22X6 port map( A => n2632, B => n101, C => n2629, D => n69
                           , Z => n561);
   U852 : HS65_LH_OAI22X6 port map( A => n2632, B => n100, C => n2629, D => n68
                           , Z => n546);
   U853 : HS65_LH_OAI22X6 port map( A => n2632, B => n99, C => n2629, D => n67,
                           Z => n531);
   U854 : HS65_LH_OAI22X6 port map( A => n2632, B => n98, C => n2629, D => n66,
                           Z => n501);
   U855 : HS65_LH_NAND4ABX3 port map( A => n851, B => n852, C => n853, D => 
                           n854, Z => n833);
   U856 : HS65_LH_AOI212X4 port map( A => registers_31_0_port, B => n2649, C =>
                           registers_30_0_port, D => n2646, E => n855, Z => 
                           n854);
   U857 : HS65_LH_AOI212X4 port map( A => registers_25_0_port, B => n2637, C =>
                           registers_24_0_port, D => n2634, E => n858, Z => 
                           n853);
   U858 : HS65_LH_MX41X7 port map( D0 => registers_16_0_port, S0 => n2625, D1 
                           => registers_17_0_port, S1 => n2622, D2 => 
                           registers_18_0_port, S2 => n2619, D3 => 
                           registers_19_0_port, S3 => n2616, Z => n852);
   U859 : HS65_LH_NAND4ABX3 port map( A => n676, B => n677, C => n678, D => 
                           n679, Z => n668);
   U860 : HS65_LH_AOI212X4 port map( A => registers_31_1_port, B => n2649, C =>
                           registers_30_1_port, D => n2646, E => n680, Z => 
                           n679);
   U861 : HS65_LH_AOI212X4 port map( A => registers_25_1_port, B => n2637, C =>
                           registers_24_1_port, D => n2634, E => n681, Z => 
                           n678);
   U862 : HS65_LH_MX41X7 port map( D0 => registers_16_1_port, S0 => n2625, D1 
                           => registers_17_1_port, S1 => n2622, D2 => 
                           registers_18_1_port, S2 => n2619, D3 => 
                           registers_19_1_port, S3 => n2616, Z => n677);
   U863 : HS65_LH_NAND4ABX3 port map( A => n511, B => n512, C => n513, D => 
                           n514, Z => n503);
   U864 : HS65_LH_AOI212X4 port map( A => registers_31_2_port, B => n2650, C =>
                           registers_30_2_port, D => n2647, E => n515, Z => 
                           n514);
   U865 : HS65_LH_AOI212X4 port map( A => registers_25_2_port, B => n2638, C =>
                           registers_24_2_port, D => n2635, E => n516, Z => 
                           n513);
   U866 : HS65_LH_MX41X7 port map( D0 => registers_16_2_port, S0 => n2626, D1 
                           => registers_17_2_port, S1 => n2623, D2 => 
                           registers_18_2_port, S2 => n2620, D3 => 
                           registers_19_2_port, S3 => n2617, Z => n512);
   U867 : HS65_LH_NAND4ABX3 port map( A => n466, B => n467, C => n468, D => 
                           n469, Z => n458);
   U868 : HS65_LH_AOI212X4 port map( A => registers_31_3_port, B => n2651, C =>
                           registers_30_3_port, D => n2647, E => n470, Z => 
                           n469);
   U869 : HS65_LH_AOI212X4 port map( A => registers_25_3_port, B => n2639, C =>
                           registers_24_3_port, D => n2635, E => n471, Z => 
                           n468);
   U870 : HS65_LH_MX41X7 port map( D0 => registers_16_3_port, S0 => n2627, D1 
                           => registers_17_3_port, S1 => n2624, D2 => 
                           registers_18_3_port, S2 => n2621, D3 => 
                           registers_19_3_port, S3 => n2618, Z => n467);
   U871 : HS65_LH_NAND4ABX3 port map( A => n451, B => n452, C => n453, D => 
                           n454, Z => n443);
   U872 : HS65_LH_AOI212X4 port map( A => registers_31_4_port, B => n2651, C =>
                           registers_30_4_port, D => n2648, E => n455, Z => 
                           n454);
   U873 : HS65_LH_AOI212X4 port map( A => registers_25_4_port, B => n2639, C =>
                           registers_24_4_port, D => n2636, E => n456, Z => 
                           n453);
   U874 : HS65_LH_MX41X7 port map( D0 => registers_16_4_port, S0 => n2627, D1 
                           => registers_17_4_port, S1 => n2624, D2 => 
                           registers_18_4_port, S2 => n2621, D3 => 
                           registers_19_4_port, S3 => n2618, Z => n452);
   U875 : HS65_LH_NAND4ABX3 port map( A => n436, B => n437, C => n438, D => 
                           n439, Z => n428);
   U876 : HS65_LH_AOI212X4 port map( A => registers_31_5_port, B => n2651, C =>
                           registers_30_5_port, D => n2648, E => n440, Z => 
                           n439);
   U877 : HS65_LH_AOI212X4 port map( A => registers_25_5_port, B => n2639, C =>
                           registers_24_5_port, D => n2636, E => n441, Z => 
                           n438);
   U878 : HS65_LH_MX41X7 port map( D0 => registers_16_5_port, S0 => n2627, D1 
                           => registers_17_5_port, S1 => n2624, D2 => 
                           registers_18_5_port, S2 => n2621, D3 => 
                           registers_19_5_port, S3 => n2618, Z => n437);
   U879 : HS65_LH_NAND4ABX3 port map( A => n421, B => n422, C => n423, D => 
                           n424, Z => n413);
   U880 : HS65_LH_AOI212X4 port map( A => registers_31_6_port, B => n2651, C =>
                           registers_30_6_port, D => n2648, E => n425, Z => 
                           n424);
   U881 : HS65_LH_AOI212X4 port map( A => registers_25_6_port, B => n2639, C =>
                           registers_24_6_port, D => n2636, E => n426, Z => 
                           n423);
   U882 : HS65_LH_MX41X7 port map( D0 => registers_16_6_port, S0 => n2627, D1 
                           => registers_17_6_port, S1 => n2624, D2 => 
                           registers_18_6_port, S2 => n2621, D3 => 
                           registers_19_6_port, S3 => n2618, Z => n422);
   U883 : HS65_LH_NAND4ABX3 port map( A => n406, B => n407, C => n408, D => 
                           n409, Z => n398);
   U884 : HS65_LH_AOI212X4 port map( A => registers_31_7_port, B => n2651, C =>
                           registers_30_7_port, D => n2648, E => n410, Z => 
                           n409);
   U885 : HS65_LH_AOI212X4 port map( A => registers_25_7_port, B => n2639, C =>
                           registers_24_7_port, D => n2636, E => n411, Z => 
                           n408);
   U886 : HS65_LH_MX41X7 port map( D0 => registers_16_7_port, S0 => n2627, D1 
                           => registers_17_7_port, S1 => n2624, D2 => 
                           registers_18_7_port, S2 => n2621, D3 => 
                           registers_19_7_port, S3 => n2618, Z => n407);
   U887 : HS65_LH_NAND4ABX3 port map( A => n391, B => n392, C => n393, D => 
                           n394, Z => n383);
   U888 : HS65_LH_AOI212X4 port map( A => registers_31_8_port, B => n2651, C =>
                           registers_30_8_port, D => n2648, E => n395, Z => 
                           n394);
   U889 : HS65_LH_AOI212X4 port map( A => registers_25_8_port, B => n2639, C =>
                           registers_24_8_port, D => n2636, E => n396, Z => 
                           n393);
   U890 : HS65_LH_MX41X7 port map( D0 => registers_16_8_port, S0 => n2627, D1 
                           => registers_17_8_port, S1 => n2624, D2 => 
                           registers_18_8_port, S2 => n2621, D3 => 
                           registers_19_8_port, S3 => n2618, Z => n392);
   U891 : HS65_LH_NAND4ABX3 port map( A => n360, B => n361, C => n362, D => 
                           n363, Z => n336);
   U892 : HS65_LH_AOI212X4 port map( A => registers_31_9_port, B => n2651, C =>
                           registers_30_9_port, D => n2648, E => n366, Z => 
                           n363);
   U893 : HS65_LH_AOI212X4 port map( A => registers_25_9_port, B => n2639, C =>
                           registers_24_9_port, D => n2636, E => n371, Z => 
                           n362);
   U894 : HS65_LH_MX41X7 port map( D0 => registers_16_9_port, S0 => n2627, D1 
                           => registers_17_9_port, S1 => n2624, D2 => 
                           registers_18_9_port, S2 => n2621, D3 => 
                           registers_19_9_port, S3 => n2618, Z => n361);
   U895 : HS65_LH_NAND4ABX3 port map( A => n826, B => n827, C => n828, D => 
                           n829, Z => n818);
   U896 : HS65_LH_AOI212X4 port map( A => registers_31_10_port, B => n2649, C 
                           => registers_30_10_port, D => n2646, E => n830, Z =>
                           n829);
   U897 : HS65_LH_AOI212X4 port map( A => registers_25_10_port, B => n2637, C 
                           => registers_24_10_port, D => n2634, E => n831, Z =>
                           n828);
   U898 : HS65_LH_MX41X7 port map( D0 => registers_16_10_port, S0 => n2625, D1 
                           => registers_17_10_port, S1 => n2622, D2 => 
                           registers_18_10_port, S2 => n2619, D3 => 
                           registers_19_10_port, S3 => n2616, Z => n827);
   U899 : HS65_LH_NAND4ABX3 port map( A => n811, B => n812, C => n813, D => 
                           n814, Z => n803);
   U900 : HS65_LH_AOI212X4 port map( A => registers_31_11_port, B => n2649, C 
                           => registers_30_11_port, D => n2646, E => n815, Z =>
                           n814);
   U901 : HS65_LH_AOI212X4 port map( A => registers_25_11_port, B => n2637, C 
                           => registers_24_11_port, D => n2634, E => n816, Z =>
                           n813);
   U902 : HS65_LH_MX41X7 port map( D0 => registers_16_11_port, S0 => n2625, D1 
                           => registers_17_11_port, S1 => n2622, D2 => 
                           registers_18_11_port, S2 => n2619, D3 => 
                           registers_19_11_port, S3 => n2616, Z => n812);
   U903 : HS65_LH_NAND4ABX3 port map( A => n796, B => n797, C => n798, D => 
                           n799, Z => n788);
   U904 : HS65_LH_AOI212X4 port map( A => registers_31_12_port, B => n2649, C 
                           => registers_30_12_port, D => n2646, E => n800, Z =>
                           n799);
   U905 : HS65_LH_AOI212X4 port map( A => registers_25_12_port, B => n2637, C 
                           => registers_24_12_port, D => n2634, E => n801, Z =>
                           n798);
   U906 : HS65_LH_MX41X7 port map( D0 => registers_16_12_port, S0 => n2625, D1 
                           => registers_17_12_port, S1 => n2622, D2 => 
                           registers_18_12_port, S2 => n2619, D3 => 
                           registers_19_12_port, S3 => n2616, Z => n797);
   U907 : HS65_LH_NAND4ABX3 port map( A => n781, B => n782, C => n783, D => 
                           n784, Z => n773);
   U908 : HS65_LH_AOI212X4 port map( A => registers_31_13_port, B => n2649, C 
                           => registers_30_13_port, D => n2646, E => n785, Z =>
                           n784);
   U909 : HS65_LH_AOI212X4 port map( A => registers_25_13_port, B => n2637, C 
                           => registers_24_13_port, D => n2634, E => n786, Z =>
                           n783);
   U910 : HS65_LH_MX41X7 port map( D0 => registers_16_13_port, S0 => n2625, D1 
                           => registers_17_13_port, S1 => n2622, D2 => 
                           registers_18_13_port, S2 => n2619, D3 => 
                           registers_19_13_port, S3 => n2616, Z => n782);
   U911 : HS65_LH_NAND4ABX3 port map( A => n766, B => n767, C => n768, D => 
                           n769, Z => n758);
   U912 : HS65_LH_AOI212X4 port map( A => registers_31_14_port, B => n2649, C 
                           => registers_30_14_port, D => n2646, E => n770, Z =>
                           n769);
   U913 : HS65_LH_AOI212X4 port map( A => registers_25_14_port, B => n2637, C 
                           => registers_24_14_port, D => n2634, E => n771, Z =>
                           n768);
   U914 : HS65_LH_MX41X7 port map( D0 => registers_16_14_port, S0 => n2625, D1 
                           => registers_17_14_port, S1 => n2622, D2 => 
                           registers_18_14_port, S2 => n2619, D3 => 
                           registers_19_14_port, S3 => n2616, Z => n767);
   U915 : HS65_LH_NAND4ABX3 port map( A => n751, B => n752, C => n753, D => 
                           n754, Z => n743);
   U916 : HS65_LH_AOI212X4 port map( A => registers_31_15_port, B => n2649, C 
                           => registers_30_15_port, D => n2646, E => n755, Z =>
                           n754);
   U917 : HS65_LH_AOI212X4 port map( A => registers_25_15_port, B => n2637, C 
                           => registers_24_15_port, D => n2634, E => n756, Z =>
                           n753);
   U918 : HS65_LH_MX41X7 port map( D0 => registers_16_15_port, S0 => n2625, D1 
                           => registers_17_15_port, S1 => n2622, D2 => 
                           registers_18_15_port, S2 => n2619, D3 => 
                           registers_19_15_port, S3 => n2616, Z => n752);
   U919 : HS65_LH_NAND4ABX3 port map( A => n736, B => n737, C => n738, D => 
                           n739, Z => n728);
   U920 : HS65_LH_AOI212X4 port map( A => registers_31_16_port, B => n2649, C 
                           => registers_30_16_port, D => n2646, E => n740, Z =>
                           n739);
   U921 : HS65_LH_AOI212X4 port map( A => registers_25_16_port, B => n2637, C 
                           => registers_24_16_port, D => n2634, E => n741, Z =>
                           n738);
   U922 : HS65_LH_MX41X7 port map( D0 => registers_16_16_port, S0 => n2625, D1 
                           => registers_17_16_port, S1 => n2622, D2 => 
                           registers_18_16_port, S2 => n2619, D3 => 
                           registers_19_16_port, S3 => n2616, Z => n737);
   U923 : HS65_LH_NAND4ABX3 port map( A => n721, B => n722, C => n723, D => 
                           n724, Z => n713);
   U924 : HS65_LH_AOI212X4 port map( A => registers_31_17_port, B => n2649, C 
                           => registers_30_17_port, D => n2646, E => n725, Z =>
                           n724);
   U925 : HS65_LH_AOI212X4 port map( A => registers_25_17_port, B => n2637, C 
                           => registers_24_17_port, D => n2634, E => n726, Z =>
                           n723);
   U926 : HS65_LH_MX41X7 port map( D0 => registers_16_17_port, S0 => n2625, D1 
                           => registers_17_17_port, S1 => n2622, D2 => 
                           registers_18_17_port, S2 => n2619, D3 => 
                           registers_19_17_port, S3 => n2616, Z => n722);
   U927 : HS65_LH_NAND4ABX3 port map( A => n706, B => n707, C => n708, D => 
                           n709, Z => n698);
   U928 : HS65_LH_AOI212X4 port map( A => registers_31_18_port, B => n2649, C 
                           => registers_30_18_port, D => n2646, E => n710, Z =>
                           n709);
   U929 : HS65_LH_AOI212X4 port map( A => registers_25_18_port, B => n2637, C 
                           => registers_24_18_port, D => n2634, E => n711, Z =>
                           n708);
   U930 : HS65_LH_MX41X7 port map( D0 => registers_16_18_port, S0 => n2625, D1 
                           => registers_17_18_port, S1 => n2622, D2 => 
                           registers_18_18_port, S2 => n2619, D3 => 
                           registers_19_18_port, S3 => n2616, Z => n707);
   U931 : HS65_LH_NAND4ABX3 port map( A => n691, B => n692, C => n693, D => 
                           n694, Z => n683);
   U932 : HS65_LH_AOI212X4 port map( A => registers_31_19_port, B => n2649, C 
                           => registers_30_19_port, D => n2646, E => n695, Z =>
                           n694);
   U933 : HS65_LH_AOI212X4 port map( A => registers_25_19_port, B => n2637, C 
                           => registers_24_19_port, D => n2634, E => n696, Z =>
                           n693);
   U934 : HS65_LH_MX41X7 port map( D0 => registers_16_19_port, S0 => n2625, D1 
                           => registers_17_19_port, S1 => n2622, D2 => 
                           registers_18_19_port, S2 => n2619, D3 => 
                           registers_19_19_port, S3 => n2616, Z => n692);
   U935 : HS65_LH_NAND4ABX3 port map( A => n661, B => n662, C => n663, D => 
                           n664, Z => n653);
   U936 : HS65_LH_AOI212X4 port map( A => registers_31_20_port, B => n2650, C 
                           => registers_30_20_port, D => n2646, E => n665, Z =>
                           n664);
   U937 : HS65_LH_AOI212X4 port map( A => registers_25_20_port, B => n2638, C 
                           => registers_24_20_port, D => n2634, E => n666, Z =>
                           n663);
   U938 : HS65_LH_MX41X7 port map( D0 => registers_16_20_port, S0 => n2626, D1 
                           => registers_17_20_port, S1 => n2623, D2 => 
                           registers_18_20_port, S2 => n2620, D3 => 
                           registers_19_20_port, S3 => n2617, Z => n662);
   U939 : HS65_LH_NAND4ABX3 port map( A => n646, B => n647, C => n648, D => 
                           n649, Z => n638);
   U940 : HS65_LH_AOI212X4 port map( A => registers_31_21_port, B => n2650, C 
                           => registers_30_21_port, D => n2647, E => n650, Z =>
                           n649);
   U941 : HS65_LH_AOI212X4 port map( A => registers_25_21_port, B => n2638, C 
                           => registers_24_21_port, D => n2635, E => n651, Z =>
                           n648);
   U942 : HS65_LH_MX41X7 port map( D0 => registers_16_21_port, S0 => n2626, D1 
                           => registers_17_21_port, S1 => n2623, D2 => 
                           registers_18_21_port, S2 => n2620, D3 => 
                           registers_19_21_port, S3 => n2617, Z => n647);
   U943 : HS65_LH_NAND4ABX3 port map( A => n631, B => n632, C => n633, D => 
                           n634, Z => n623);
   U944 : HS65_LH_AOI212X4 port map( A => registers_31_22_port, B => n2650, C 
                           => registers_30_22_port, D => n2647, E => n635, Z =>
                           n634);
   U945 : HS65_LH_AOI212X4 port map( A => registers_25_22_port, B => n2638, C 
                           => registers_24_22_port, D => n2635, E => n636, Z =>
                           n633);
   U946 : HS65_LH_MX41X7 port map( D0 => registers_16_22_port, S0 => n2626, D1 
                           => registers_17_22_port, S1 => n2623, D2 => 
                           registers_18_22_port, S2 => n2620, D3 => 
                           registers_19_22_port, S3 => n2617, Z => n632);
   U947 : HS65_LH_NAND4ABX3 port map( A => n616, B => n617, C => n618, D => 
                           n619, Z => n608);
   U948 : HS65_LH_AOI212X4 port map( A => registers_31_23_port, B => n2650, C 
                           => registers_30_23_port, D => n2647, E => n620, Z =>
                           n619);
   U949 : HS65_LH_AOI212X4 port map( A => registers_25_23_port, B => n2638, C 
                           => registers_24_23_port, D => n2635, E => n621, Z =>
                           n618);
   U950 : HS65_LH_MX41X7 port map( D0 => registers_16_23_port, S0 => n2626, D1 
                           => registers_17_23_port, S1 => n2623, D2 => 
                           registers_18_23_port, S2 => n2620, D3 => 
                           registers_19_23_port, S3 => n2617, Z => n617);
   U951 : HS65_LH_NAND4ABX3 port map( A => n601, B => n602, C => n603, D => 
                           n604, Z => n593);
   U952 : HS65_LH_AOI212X4 port map( A => registers_31_24_port, B => n2650, C 
                           => registers_30_24_port, D => n2647, E => n605, Z =>
                           n604);
   U953 : HS65_LH_AOI212X4 port map( A => registers_25_24_port, B => n2638, C 
                           => registers_24_24_port, D => n2635, E => n606, Z =>
                           n603);
   U954 : HS65_LH_MX41X7 port map( D0 => registers_16_24_port, S0 => n2626, D1 
                           => registers_17_24_port, S1 => n2623, D2 => 
                           registers_18_24_port, S2 => n2620, D3 => 
                           registers_19_24_port, S3 => n2617, Z => n602);
   U955 : HS65_LH_NAND4ABX3 port map( A => n586, B => n587, C => n588, D => 
                           n589, Z => n578);
   U956 : HS65_LH_AOI212X4 port map( A => registers_31_25_port, B => n2650, C 
                           => registers_30_25_port, D => n2647, E => n590, Z =>
                           n589);
   U957 : HS65_LH_AOI212X4 port map( A => registers_25_25_port, B => n2638, C 
                           => registers_24_25_port, D => n2635, E => n591, Z =>
                           n588);
   U958 : HS65_LH_MX41X7 port map( D0 => registers_16_25_port, S0 => n2626, D1 
                           => registers_17_25_port, S1 => n2623, D2 => 
                           registers_18_25_port, S2 => n2620, D3 => 
                           registers_19_25_port, S3 => n2617, Z => n587);
   U959 : HS65_LH_NAND4ABX3 port map( A => n571, B => n572, C => n573, D => 
                           n574, Z => n563);
   U960 : HS65_LH_AOI212X4 port map( A => registers_31_26_port, B => n2650, C 
                           => registers_30_26_port, D => n2647, E => n575, Z =>
                           n574);
   U961 : HS65_LH_AOI212X4 port map( A => registers_25_26_port, B => n2638, C 
                           => registers_24_26_port, D => n2635, E => n576, Z =>
                           n573);
   U962 : HS65_LH_MX41X7 port map( D0 => registers_16_26_port, S0 => n2626, D1 
                           => registers_17_26_port, S1 => n2623, D2 => 
                           registers_18_26_port, S2 => n2620, D3 => 
                           registers_19_26_port, S3 => n2617, Z => n572);
   U963 : HS65_LH_NAND4ABX3 port map( A => n556, B => n557, C => n558, D => 
                           n559, Z => n548);
   U964 : HS65_LH_AOI212X4 port map( A => registers_31_27_port, B => n2650, C 
                           => registers_30_27_port, D => n2647, E => n560, Z =>
                           n559);
   U965 : HS65_LH_AOI212X4 port map( A => registers_25_27_port, B => n2638, C 
                           => registers_24_27_port, D => n2635, E => n561, Z =>
                           n558);
   U966 : HS65_LH_MX41X7 port map( D0 => registers_16_27_port, S0 => n2626, D1 
                           => registers_17_27_port, S1 => n2623, D2 => 
                           registers_18_27_port, S2 => n2620, D3 => 
                           registers_19_27_port, S3 => n2617, Z => n557);
   U967 : HS65_LH_NAND4ABX3 port map( A => n541, B => n542, C => n543, D => 
                           n544, Z => n533);
   U968 : HS65_LH_AOI212X4 port map( A => registers_31_28_port, B => n2650, C 
                           => registers_30_28_port, D => n2647, E => n545, Z =>
                           n544);
   U969 : HS65_LH_AOI212X4 port map( A => registers_25_28_port, B => n2638, C 
                           => registers_24_28_port, D => n2635, E => n546, Z =>
                           n543);
   U970 : HS65_LH_MX41X7 port map( D0 => registers_16_28_port, S0 => n2626, D1 
                           => registers_17_28_port, S1 => n2623, D2 => 
                           registers_18_28_port, S2 => n2620, D3 => 
                           registers_19_28_port, S3 => n2617, Z => n542);
   U971 : HS65_LH_NAND4ABX3 port map( A => n526, B => n527, C => n528, D => 
                           n529, Z => n518);
   U972 : HS65_LH_AOI212X4 port map( A => registers_31_29_port, B => n2650, C 
                           => registers_30_29_port, D => n2647, E => n530, Z =>
                           n529);
   U973 : HS65_LH_AOI212X4 port map( A => registers_25_29_port, B => n2638, C 
                           => registers_24_29_port, D => n2635, E => n531, Z =>
                           n528);
   U974 : HS65_LH_MX41X7 port map( D0 => registers_16_29_port, S0 => n2626, D1 
                           => registers_17_29_port, S1 => n2623, D2 => 
                           registers_18_29_port, S2 => n2620, D3 => 
                           registers_19_29_port, S3 => n2617, Z => n527);
   U975 : HS65_LH_NAND4ABX3 port map( A => n496, B => n497, C => n498, D => 
                           n499, Z => n488);
   U976 : HS65_LH_AOI212X4 port map( A => registers_31_30_port, B => n2650, C 
                           => registers_30_30_port, D => n2647, E => n500, Z =>
                           n499);
   U977 : HS65_LH_AOI212X4 port map( A => registers_25_30_port, B => n2638, C 
                           => registers_24_30_port, D => n2635, E => n501, Z =>
                           n498);
   U978 : HS65_LH_MX41X7 port map( D0 => registers_16_30_port, S0 => n2626, D1 
                           => registers_17_30_port, S1 => n2623, D2 => 
                           registers_18_30_port, S2 => n2620, D3 => 
                           registers_19_30_port, S3 => n2617, Z => n497);
   U979 : HS65_LH_NAND4ABX3 port map( A => n481, B => n482, C => n483, D => 
                           n484, Z => n473);
   U980 : HS65_LH_AOI212X4 port map( A => registers_31_31_port, B => n2651, C 
                           => registers_30_31_port, D => n2647, E => n485, Z =>
                           n484);
   U981 : HS65_LH_AOI212X4 port map( A => registers_25_31_port, B => n2639, C 
                           => registers_24_31_port, D => n2635, E => n486, Z =>
                           n483);
   U982 : HS65_LH_MX41X7 port map( D0 => registers_16_31_port, S0 => n2627, D1 
                           => registers_17_31_port, S1 => n2624, D2 => 
                           registers_18_31_port, S2 => n2621, D3 => 
                           registers_19_31_port, S3 => n2618, Z => n482);
   U983 : HS65_LH_NAND4ABX3 port map( A => n1379, B => n1380, C => n1381, D => 
                           n1382, Z => n1361);
   U984 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_0_port, C =>
                           n2553, D => registers_30_0_port, E => n1383, Z => 
                           n1382);
   U985 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_0_port, C =>
                           n2541, D => registers_24_0_port, E => n1386, Z => 
                           n1381);
   U986 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_0_port, D1 
                           => n2529, S1 => registers_17_0_port, D2 => n2526, S2
                           => registers_18_0_port, D3 => n2523, S3 => 
                           registers_19_0_port, Z => n1380);
   U987 : HS65_LH_NAND4ABX3 port map( A => n1204, B => n1205, C => n1206, D => 
                           n1207, Z => n1196);
   U988 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_1_port, C =>
                           n2553, D => registers_30_1_port, E => n1208, Z => 
                           n1207);
   U989 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_1_port, C =>
                           n2541, D => registers_24_1_port, E => n1209, Z => 
                           n1206);
   U990 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_1_port, D1 
                           => n2529, S1 => registers_17_1_port, D2 => n2526, S2
                           => registers_18_1_port, D3 => n2523, S3 => 
                           registers_19_1_port, Z => n1205);
   U991 : HS65_LH_NAND4ABX3 port map( A => n1039, B => n1040, C => n1041, D => 
                           n1042, Z => n1031);
   U992 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_2_port, C =>
                           n2554, D => registers_30_2_port, E => n1043, Z => 
                           n1042);
   U993 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_2_port, C =>
                           n2542, D => registers_24_2_port, E => n1044, Z => 
                           n1041);
   U994 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_2_port, D1 
                           => n2530, S1 => registers_17_2_port, D2 => n2527, S2
                           => registers_18_2_port, D3 => n2524, S3 => 
                           registers_19_2_port, Z => n1040);
   U995 : HS65_LH_NAND4ABX3 port map( A => n994, B => n995, C => n996, D => 
                           n997, Z => n986);
   U996 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_3_port, C =>
                           n2554, D => registers_30_3_port, E => n998, Z => 
                           n997);
   U997 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_3_port, C =>
                           n2542, D => registers_24_3_port, E => n999, Z => 
                           n996);
   U998 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_3_port, D1 
                           => n2531, S1 => registers_17_3_port, D2 => n2527, S2
                           => registers_18_3_port, D3 => n2525, S3 => 
                           registers_19_3_port, Z => n995);
   U999 : HS65_LH_NAND4ABX3 port map( A => n979, B => n980, C => n981, D => 
                           n982, Z => n971);
   U1000 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_4_port, C 
                           => n2555, D => registers_30_4_port, E => n983, Z => 
                           n982);
   U1001 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_4_port, C 
                           => n2543, D => registers_24_4_port, E => n984, Z => 
                           n981);
   U1002 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_4_port, D1 
                           => n2531, S1 => registers_17_4_port, D2 => n2528, S2
                           => registers_18_4_port, D3 => n2525, S3 => 
                           registers_19_4_port, Z => n980);
   U1003 : HS65_LH_NAND4ABX3 port map( A => n964, B => n965, C => n966, D => 
                           n967, Z => n956);
   U1004 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_5_port, C 
                           => n2555, D => registers_30_5_port, E => n968, Z => 
                           n967);
   U1005 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_5_port, C 
                           => n2543, D => registers_24_5_port, E => n969, Z => 
                           n966);
   U1006 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_5_port, D1 
                           => n2531, S1 => registers_17_5_port, D2 => n2528, S2
                           => registers_18_5_port, D3 => n2525, S3 => 
                           registers_19_5_port, Z => n965);
   U1007 : HS65_LH_NAND4ABX3 port map( A => n949, B => n950, C => n951, D => 
                           n952, Z => n941);
   U1008 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_6_port, C 
                           => n2555, D => registers_30_6_port, E => n953, Z => 
                           n952);
   U1009 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_6_port, C 
                           => n2543, D => registers_24_6_port, E => n954, Z => 
                           n951);
   U1010 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_6_port, D1 
                           => n2531, S1 => registers_17_6_port, D2 => n2528, S2
                           => registers_18_6_port, D3 => n2525, S3 => 
                           registers_19_6_port, Z => n950);
   U1011 : HS65_LH_NAND4ABX3 port map( A => n934, B => n935, C => n936, D => 
                           n937, Z => n926);
   U1012 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_7_port, C 
                           => n2555, D => registers_30_7_port, E => n938, Z => 
                           n937);
   U1013 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_7_port, C 
                           => n2543, D => registers_24_7_port, E => n939, Z => 
                           n936);
   U1014 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_7_port, D1 
                           => n2531, S1 => registers_17_7_port, D2 => n2528, S2
                           => registers_18_7_port, D3 => n2525, S3 => 
                           registers_19_7_port, Z => n935);
   U1015 : HS65_LH_NAND4ABX3 port map( A => n919, B => n920, C => n921, D => 
                           n922, Z => n911);
   U1016 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_8_port, C 
                           => n2555, D => registers_30_8_port, E => n923, Z => 
                           n922);
   U1017 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_8_port, C 
                           => n2543, D => registers_24_8_port, E => n924, Z => 
                           n921);
   U1018 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_8_port, D1 
                           => n2531, S1 => registers_17_8_port, D2 => n2528, S2
                           => registers_18_8_port, D3 => n2525, S3 => 
                           registers_19_8_port, Z => n920);
   U1019 : HS65_LH_NAND4ABX3 port map( A => n888, B => n889, C => n890, D => 
                           n891, Z => n864);
   U1020 : HS65_LH_AOI212X4 port map( A => n2558, B => registers_31_9_port, C 
                           => n2555, D => registers_30_9_port, E => n894, Z => 
                           n891);
   U1021 : HS65_LH_AOI212X4 port map( A => n2546, B => registers_25_9_port, C 
                           => n2543, D => registers_24_9_port, E => n899, Z => 
                           n890);
   U1022 : HS65_LH_MX41X7 port map( D0 => n2534, S0 => registers_16_9_port, D1 
                           => n2531, S1 => registers_17_9_port, D2 => n2528, S2
                           => registers_18_9_port, D3 => n2525, S3 => 
                           registers_19_9_port, Z => n889);
   U1023 : HS65_LH_NAND4ABX3 port map( A => n1354, B => n1355, C => n1356, D =>
                           n1357, Z => n1346);
   U1024 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_10_port, C 
                           => n2553, D => registers_30_10_port, E => n1358, Z 
                           => n1357);
   U1025 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_10_port, C 
                           => n2541, D => registers_24_10_port, E => n1359, Z 
                           => n1356);
   U1026 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_10_port, D1
                           => n2529, S1 => registers_17_10_port, D2 => n2526, 
                           S2 => registers_18_10_port, D3 => n2523, S3 => 
                           registers_19_10_port, Z => n1355);
   U1027 : HS65_LH_NAND4ABX3 port map( A => n1339, B => n1340, C => n1341, D =>
                           n1342, Z => n1331);
   U1028 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_11_port, C 
                           => n2553, D => registers_30_11_port, E => n1343, Z 
                           => n1342);
   U1029 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_11_port, C 
                           => n2541, D => registers_24_11_port, E => n1344, Z 
                           => n1341);
   U1030 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_11_port, D1
                           => n2529, S1 => registers_17_11_port, D2 => n2526, 
                           S2 => registers_18_11_port, D3 => n2523, S3 => 
                           registers_19_11_port, Z => n1340);
   U1031 : HS65_LH_NAND4ABX3 port map( A => n1324, B => n1325, C => n1326, D =>
                           n1327, Z => n1316);
   U1032 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_12_port, C 
                           => n2553, D => registers_30_12_port, E => n1328, Z 
                           => n1327);
   U1033 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_12_port, C 
                           => n2541, D => registers_24_12_port, E => n1329, Z 
                           => n1326);
   U1034 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_12_port, D1
                           => n2529, S1 => registers_17_12_port, D2 => n2526, 
                           S2 => registers_18_12_port, D3 => n2523, S3 => 
                           registers_19_12_port, Z => n1325);
   U1035 : HS65_LH_NAND4ABX3 port map( A => n1309, B => n1310, C => n1311, D =>
                           n1312, Z => n1301);
   U1036 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_13_port, C 
                           => n2553, D => registers_30_13_port, E => n1313, Z 
                           => n1312);
   U1037 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_13_port, C 
                           => n2541, D => registers_24_13_port, E => n1314, Z 
                           => n1311);
   U1038 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_13_port, D1
                           => n2529, S1 => registers_17_13_port, D2 => n2526, 
                           S2 => registers_18_13_port, D3 => n2523, S3 => 
                           registers_19_13_port, Z => n1310);
   U1039 : HS65_LH_NAND4ABX3 port map( A => n1294, B => n1295, C => n1296, D =>
                           n1297, Z => n1286);
   U1040 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_14_port, C 
                           => n2553, D => registers_30_14_port, E => n1298, Z 
                           => n1297);
   U1041 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_14_port, C 
                           => n2541, D => registers_24_14_port, E => n1299, Z 
                           => n1296);
   U1042 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_14_port, D1
                           => n2529, S1 => registers_17_14_port, D2 => n2526, 
                           S2 => registers_18_14_port, D3 => n2523, S3 => 
                           registers_19_14_port, Z => n1295);
   U1043 : HS65_LH_NAND4ABX3 port map( A => n1279, B => n1280, C => n1281, D =>
                           n1282, Z => n1271);
   U1044 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_15_port, C 
                           => n2553, D => registers_30_15_port, E => n1283, Z 
                           => n1282);
   U1045 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_15_port, C 
                           => n2541, D => registers_24_15_port, E => n1284, Z 
                           => n1281);
   U1046 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_15_port, D1
                           => n2529, S1 => registers_17_15_port, D2 => n2526, 
                           S2 => registers_18_15_port, D3 => n2523, S3 => 
                           registers_19_15_port, Z => n1280);
   U1047 : HS65_LH_NAND4ABX3 port map( A => n1264, B => n1265, C => n1266, D =>
                           n1267, Z => n1256);
   U1048 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_16_port, C 
                           => n2553, D => registers_30_16_port, E => n1268, Z 
                           => n1267);
   U1049 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_16_port, C 
                           => n2541, D => registers_24_16_port, E => n1269, Z 
                           => n1266);
   U1050 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_16_port, D1
                           => n2529, S1 => registers_17_16_port, D2 => n2526, 
                           S2 => registers_18_16_port, D3 => n2523, S3 => 
                           registers_19_16_port, Z => n1265);
   U1051 : HS65_LH_NAND4ABX3 port map( A => n1249, B => n1250, C => n1251, D =>
                           n1252, Z => n1241);
   U1052 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_17_port, C 
                           => n2553, D => registers_30_17_port, E => n1253, Z 
                           => n1252);
   U1053 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_17_port, C 
                           => n2541, D => registers_24_17_port, E => n1254, Z 
                           => n1251);
   U1054 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_17_port, D1
                           => n2529, S1 => registers_17_17_port, D2 => n2526, 
                           S2 => registers_18_17_port, D3 => n2523, S3 => 
                           registers_19_17_port, Z => n1250);
   U1055 : HS65_LH_NAND4ABX3 port map( A => n1234, B => n1235, C => n1236, D =>
                           n1237, Z => n1226);
   U1056 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_18_port, C 
                           => n2553, D => registers_30_18_port, E => n1238, Z 
                           => n1237);
   U1057 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_18_port, C 
                           => n2541, D => registers_24_18_port, E => n1239, Z 
                           => n1236);
   U1058 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_18_port, D1
                           => n2529, S1 => registers_17_18_port, D2 => n2526, 
                           S2 => registers_18_18_port, D3 => n2523, S3 => 
                           registers_19_18_port, Z => n1235);
   U1059 : HS65_LH_NAND4ABX3 port map( A => n1219, B => n1220, C => n1221, D =>
                           n1222, Z => n1211);
   U1060 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_19_port, C 
                           => n2553, D => registers_30_19_port, E => n1223, Z 
                           => n1222);
   U1061 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_19_port, C 
                           => n2541, D => registers_24_19_port, E => n1224, Z 
                           => n1221);
   U1062 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_19_port, D1
                           => n2529, S1 => registers_17_19_port, D2 => n2526, 
                           S2 => registers_18_19_port, D3 => n2523, S3 => 
                           registers_19_19_port, Z => n1220);
   U1063 : HS65_LH_NAND4ABX3 port map( A => n1189, B => n1190, C => n1191, D =>
                           n1192, Z => n1181);
   U1064 : HS65_LH_AOI212X4 port map( A => n2556, B => registers_31_20_port, C 
                           => n2553, D => registers_30_20_port, E => n1193, Z 
                           => n1192);
   U1065 : HS65_LH_AOI212X4 port map( A => n2544, B => registers_25_20_port, C 
                           => n2541, D => registers_24_20_port, E => n1194, Z 
                           => n1191);
   U1066 : HS65_LH_MX41X7 port map( D0 => n2532, S0 => registers_16_20_port, D1
                           => n2530, S1 => registers_17_20_port, D2 => n2526, 
                           S2 => registers_18_20_port, D3 => n2524, S3 => 
                           registers_19_20_port, Z => n1190);
   U1067 : HS65_LH_NAND4ABX3 port map( A => n1174, B => n1175, C => n1176, D =>
                           n1177, Z => n1166);
   U1068 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_21_port, C 
                           => n2554, D => registers_30_21_port, E => n1178, Z 
                           => n1177);
   U1069 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_21_port, C 
                           => n2542, D => registers_24_21_port, E => n1179, Z 
                           => n1176);
   U1070 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_21_port, D1
                           => n2530, S1 => registers_17_21_port, D2 => n2527, 
                           S2 => registers_18_21_port, D3 => n2524, S3 => 
                           registers_19_21_port, Z => n1175);
   U1071 : HS65_LH_NAND4ABX3 port map( A => n1159, B => n1160, C => n1161, D =>
                           n1162, Z => n1151);
   U1072 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_22_port, C 
                           => n2554, D => registers_30_22_port, E => n1163, Z 
                           => n1162);
   U1073 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_22_port, C 
                           => n2542, D => registers_24_22_port, E => n1164, Z 
                           => n1161);
   U1074 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_22_port, D1
                           => n2530, S1 => registers_17_22_port, D2 => n2527, 
                           S2 => registers_18_22_port, D3 => n2524, S3 => 
                           registers_19_22_port, Z => n1160);
   U1075 : HS65_LH_NAND4ABX3 port map( A => n1144, B => n1145, C => n1146, D =>
                           n1147, Z => n1136);
   U1076 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_23_port, C 
                           => n2554, D => registers_30_23_port, E => n1148, Z 
                           => n1147);
   U1077 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_23_port, C 
                           => n2542, D => registers_24_23_port, E => n1149, Z 
                           => n1146);
   U1078 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_23_port, D1
                           => n2530, S1 => registers_17_23_port, D2 => n2527, 
                           S2 => registers_18_23_port, D3 => n2524, S3 => 
                           registers_19_23_port, Z => n1145);
   U1079 : HS65_LH_NAND4ABX3 port map( A => n1129, B => n1130, C => n1131, D =>
                           n1132, Z => n1121);
   U1080 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_24_port, C 
                           => n2554, D => registers_30_24_port, E => n1133, Z 
                           => n1132);
   U1081 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_24_port, C 
                           => n2542, D => registers_24_24_port, E => n1134, Z 
                           => n1131);
   U1082 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_24_port, D1
                           => n2530, S1 => registers_17_24_port, D2 => n2527, 
                           S2 => registers_18_24_port, D3 => n2524, S3 => 
                           registers_19_24_port, Z => n1130);
   U1083 : HS65_LH_NAND4ABX3 port map( A => n1114, B => n1115, C => n1116, D =>
                           n1117, Z => n1106);
   U1084 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_25_port, C 
                           => n2554, D => registers_30_25_port, E => n1118, Z 
                           => n1117);
   U1085 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_25_port, C 
                           => n2542, D => registers_24_25_port, E => n1119, Z 
                           => n1116);
   U1086 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_25_port, D1
                           => n2530, S1 => registers_17_25_port, D2 => n2527, 
                           S2 => registers_18_25_port, D3 => n2524, S3 => 
                           registers_19_25_port, Z => n1115);
   U1087 : HS65_LH_NAND4ABX3 port map( A => n1099, B => n1100, C => n1101, D =>
                           n1102, Z => n1091);
   U1088 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_26_port, C 
                           => n2554, D => registers_30_26_port, E => n1103, Z 
                           => n1102);
   U1089 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_26_port, C 
                           => n2542, D => registers_24_26_port, E => n1104, Z 
                           => n1101);
   U1090 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_26_port, D1
                           => n2530, S1 => registers_17_26_port, D2 => n2527, 
                           S2 => registers_18_26_port, D3 => n2524, S3 => 
                           registers_19_26_port, Z => n1100);
   U1091 : HS65_LH_NAND4ABX3 port map( A => n1084, B => n1085, C => n1086, D =>
                           n1087, Z => n1076);
   U1092 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_27_port, C 
                           => n2554, D => registers_30_27_port, E => n1088, Z 
                           => n1087);
   U1093 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_27_port, C 
                           => n2542, D => registers_24_27_port, E => n1089, Z 
                           => n1086);
   U1094 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_27_port, D1
                           => n2530, S1 => registers_17_27_port, D2 => n2527, 
                           S2 => registers_18_27_port, D3 => n2524, S3 => 
                           registers_19_27_port, Z => n1085);
   U1095 : HS65_LH_NAND4ABX3 port map( A => n1069, B => n1070, C => n1071, D =>
                           n1072, Z => n1061);
   U1096 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_28_port, C 
                           => n2554, D => registers_30_28_port, E => n1073, Z 
                           => n1072);
   U1097 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_28_port, C 
                           => n2542, D => registers_24_28_port, E => n1074, Z 
                           => n1071);
   U1098 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_28_port, D1
                           => n2530, S1 => registers_17_28_port, D2 => n2527, 
                           S2 => registers_18_28_port, D3 => n2524, S3 => 
                           registers_19_28_port, Z => n1070);
   U1099 : HS65_LH_NAND4ABX3 port map( A => n1054, B => n1055, C => n1056, D =>
                           n1057, Z => n1046);
   U1100 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_29_port, C 
                           => n2554, D => registers_30_29_port, E => n1058, Z 
                           => n1057);
   U1101 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_29_port, C 
                           => n2542, D => registers_24_29_port, E => n1059, Z 
                           => n1056);
   U1102 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_29_port, D1
                           => n2530, S1 => registers_17_29_port, D2 => n2527, 
                           S2 => registers_18_29_port, D3 => n2524, S3 => 
                           registers_19_29_port, Z => n1055);
   U1103 : HS65_LH_NAND4ABX3 port map( A => n1024, B => n1025, C => n1026, D =>
                           n1027, Z => n1016);
   U1104 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_30_port, C 
                           => n2554, D => registers_30_30_port, E => n1028, Z 
                           => n1027);
   U1105 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_30_port, C 
                           => n2542, D => registers_24_30_port, E => n1029, Z 
                           => n1026);
   U1106 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_30_port, D1
                           => n2530, S1 => registers_17_30_port, D2 => n2527, 
                           S2 => registers_18_30_port, D3 => n2524, S3 => 
                           registers_19_30_port, Z => n1025);
   U1107 : HS65_LH_NAND4ABX3 port map( A => n1009, B => n1010, C => n1011, D =>
                           n1012, Z => n1001);
   U1108 : HS65_LH_AOI212X4 port map( A => n2557, B => registers_31_31_port, C 
                           => n2554, D => registers_30_31_port, E => n1013, Z 
                           => n1012);
   U1109 : HS65_LH_AOI212X4 port map( A => n2545, B => registers_25_31_port, C 
                           => n2542, D => registers_24_31_port, E => n1014, Z 
                           => n1011);
   U1110 : HS65_LH_MX41X7 port map( D0 => n2533, S0 => registers_16_31_port, D1
                           => n2531, S1 => registers_17_31_port, D2 => n2527, 
                           S2 => registers_18_31_port, D3 => n2525, S3 => 
                           registers_19_31_port, Z => n1010);
   U1111 : HS65_LH_NAND4ABX3 port map( A => n820, B => n821, C => n822, D => 
                           n823, Z => n819);
   U1112 : HS65_LH_NAND3X5 port map( A => n2968, B => n2969, C => n2970, Z => 
                           n821);
   U1113 : HS65_LH_AOI212X4 port map( A => registers_13_10_port, B => n2694, C 
                           => registers_12_10_port, D => n2691, E => n824, Z =>
                           n823);
   U1114 : HS65_LH_AOI212X4 port map( A => registers_11_10_port, B => n2682, C 
                           => registers_10_10_port, D => n2679, E => n825, Z =>
                           n822);
   U1115 : HS65_LH_AND2X4 port map( A => n847, B => regfile_i(40), Z => n840);
   U1116 : HS65_LH_AND2X4 port map( A => n1375, B => regfile_i(45), Z => n1368)
                           ;
   U1117 : HS65_LH_AND2X4 port map( A => n859, B => regfile_i(40), Z => n856);
   U1118 : HS65_LH_AND2X4 port map( A => n1387, B => regfile_i(45), Z => n1384)
                           ;
   U1119 : HS65_LH_AND2X4 port map( A => n862, B => regfile_i(40), Z => n860);
   U1120 : HS65_LH_AND2X4 port map( A => n850, B => regfile_i(40), Z => n848);
   U1121 : HS65_LH_AND2X4 port map( A => n1390, B => regfile_i(45), Z => n1388)
                           ;
   U1122 : HS65_LH_AND2X4 port map( A => n1378, B => regfile_i(45), Z => n1376)
                           ;
   U1123 : HS65_LH_NOR2X6 port map( A => n2902, B => regfile_i(43), Z => n862);
   U1124 : HS65_LH_NOR2X6 port map( A => n2907, B => regfile_i(48), Z => n1390)
                           ;
   U1125 : HS65_LH_NOR2X6 port map( A => regfile_i(43), B => regfile_i(44), Z 
                           => n850);
   U1126 : HS65_LH_NOR2X6 port map( A => n2901, B => regfile_i(44), Z => n847);
   U1127 : HS65_LH_NOR2X6 port map( A => regfile_i(48), B => regfile_i(49), Z 
                           => n1378);
   U1128 : HS65_LH_NOR2X6 port map( A => n2906, B => regfile_i(49), Z => n1375)
                           ;
   U1129 : HS65_LH_MX41X7 port map( D0 => registers_20_0_port, S0 => n2613, D1 
                           => registers_21_0_port, S1 => n2610, D2 => 
                           registers_22_0_port, S2 => n2607, D3 => 
                           registers_23_0_port, S3 => n2604, Z => n851);
   U1130 : HS65_LH_MX41X7 port map( D0 => registers_4_0_port, S0 => n2661, D1 
                           => registers_5_0_port, S1 => n2658, D2 => 
                           registers_6_0_port, S2 => n2655, D3 => 
                           registers_7_0_port, S3 => n2652, Z => n835);
   U1131 : HS65_LH_MX41X7 port map( D0 => registers_20_1_port, S0 => n2613, D1 
                           => registers_21_1_port, S1 => n2610, D2 => 
                           registers_22_1_port, S2 => n2607, D3 => 
                           registers_23_1_port, S3 => n2604, Z => n676);
   U1132 : HS65_LH_MX41X7 port map( D0 => registers_4_1_port, S0 => n2661, D1 
                           => registers_5_1_port, S1 => n2658, D2 => 
                           registers_6_1_port, S2 => n2655, D3 => 
                           registers_7_1_port, S3 => n2652, Z => n670);
   U1133 : HS65_LH_MX41X7 port map( D0 => registers_20_2_port, S0 => n2614, D1 
                           => registers_21_2_port, S1 => n2611, D2 => 
                           registers_22_2_port, S2 => n2608, D3 => 
                           registers_23_2_port, S3 => n2605, Z => n511);
   U1134 : HS65_LH_MX41X7 port map( D0 => registers_4_2_port, S0 => n2662, D1 
                           => registers_5_2_port, S1 => n2659, D2 => 
                           registers_6_2_port, S2 => n2656, D3 => 
                           registers_7_2_port, S3 => n2653, Z => n505);
   U1135 : HS65_LH_MX41X7 port map( D0 => registers_20_3_port, S0 => n2615, D1 
                           => registers_21_3_port, S1 => n2612, D2 => 
                           registers_22_3_port, S2 => n2609, D3 => 
                           registers_23_3_port, S3 => n2606, Z => n466);
   U1136 : HS65_LH_MX41X7 port map( D0 => registers_4_3_port, S0 => n2663, D1 
                           => registers_5_3_port, S1 => n2660, D2 => 
                           registers_6_3_port, S2 => n2657, D3 => 
                           registers_7_3_port, S3 => n2654, Z => n460);
   U1137 : HS65_LH_MX41X7 port map( D0 => registers_20_4_port, S0 => n2615, D1 
                           => registers_21_4_port, S1 => n2612, D2 => 
                           registers_22_4_port, S2 => n2609, D3 => 
                           registers_23_4_port, S3 => n2606, Z => n451);
   U1138 : HS65_LH_MX41X7 port map( D0 => registers_4_4_port, S0 => n2663, D1 
                           => registers_5_4_port, S1 => n2660, D2 => 
                           registers_6_4_port, S2 => n2657, D3 => 
                           registers_7_4_port, S3 => n2654, Z => n445);
   U1139 : HS65_LH_MX41X7 port map( D0 => registers_20_5_port, S0 => n2615, D1 
                           => registers_21_5_port, S1 => n2612, D2 => 
                           registers_22_5_port, S2 => n2609, D3 => 
                           registers_23_5_port, S3 => n2606, Z => n436);
   U1140 : HS65_LH_MX41X7 port map( D0 => registers_4_5_port, S0 => n2663, D1 
                           => registers_5_5_port, S1 => n2660, D2 => 
                           registers_6_5_port, S2 => n2657, D3 => 
                           registers_7_5_port, S3 => n2654, Z => n430);
   U1141 : HS65_LH_MX41X7 port map( D0 => registers_20_6_port, S0 => n2615, D1 
                           => registers_21_6_port, S1 => n2612, D2 => 
                           registers_22_6_port, S2 => n2609, D3 => 
                           registers_23_6_port, S3 => n2606, Z => n421);
   U1142 : HS65_LH_MX41X7 port map( D0 => registers_4_6_port, S0 => n2663, D1 
                           => registers_5_6_port, S1 => n2660, D2 => 
                           registers_6_6_port, S2 => n2657, D3 => 
                           registers_7_6_port, S3 => n2654, Z => n415);
   U1143 : HS65_LH_MX41X7 port map( D0 => registers_20_7_port, S0 => n2615, D1 
                           => registers_21_7_port, S1 => n2612, D2 => 
                           registers_22_7_port, S2 => n2609, D3 => 
                           registers_23_7_port, S3 => n2606, Z => n406);
   U1144 : HS65_LH_MX41X7 port map( D0 => registers_4_7_port, S0 => n2663, D1 
                           => registers_5_7_port, S1 => n2660, D2 => 
                           registers_6_7_port, S2 => n2657, D3 => 
                           registers_7_7_port, S3 => n2654, Z => n400);
   U1145 : HS65_LH_MX41X7 port map( D0 => registers_20_8_port, S0 => n2615, D1 
                           => registers_21_8_port, S1 => n2612, D2 => 
                           registers_22_8_port, S2 => n2609, D3 => 
                           registers_23_8_port, S3 => n2606, Z => n391);
   U1146 : HS65_LH_MX41X7 port map( D0 => registers_4_8_port, S0 => n2663, D1 
                           => registers_5_8_port, S1 => n2660, D2 => 
                           registers_6_8_port, S2 => n2657, D3 => 
                           registers_7_8_port, S3 => n2654, Z => n385);
   U1147 : HS65_LH_MX41X7 port map( D0 => registers_20_9_port, S0 => n2615, D1 
                           => registers_21_9_port, S1 => n2612, D2 => 
                           registers_22_9_port, S2 => n2609, D3 => 
                           registers_23_9_port, S3 => n2606, Z => n360);
   U1148 : HS65_LH_MX41X7 port map( D0 => registers_4_9_port, S0 => n2663, D1 
                           => registers_5_9_port, S1 => n2660, D2 => 
                           registers_6_9_port, S2 => n2657, D3 => 
                           registers_7_9_port, S3 => n2654, Z => n338);
   U1149 : HS65_LH_MX41X7 port map( D0 => registers_20_10_port, S0 => n2613, D1
                           => registers_21_10_port, S1 => n2610, D2 => 
                           registers_22_10_port, S2 => n2607, D3 => 
                           registers_23_10_port, S3 => n2604, Z => n826);
   U1150 : HS65_LH_MX41X7 port map( D0 => registers_4_10_port, S0 => n2661, D1 
                           => registers_5_10_port, S1 => n2658, D2 => 
                           registers_6_10_port, S2 => n2655, D3 => 
                           registers_7_10_port, S3 => n2652, Z => n820);
   U1151 : HS65_LH_MX41X7 port map( D0 => registers_20_11_port, S0 => n2613, D1
                           => registers_21_11_port, S1 => n2610, D2 => 
                           registers_22_11_port, S2 => n2607, D3 => 
                           registers_23_11_port, S3 => n2604, Z => n811);
   U1152 : HS65_LH_MX41X7 port map( D0 => registers_4_11_port, S0 => n2661, D1 
                           => registers_5_11_port, S1 => n2658, D2 => 
                           registers_6_11_port, S2 => n2655, D3 => 
                           registers_7_11_port, S3 => n2652, Z => n805);
   U1153 : HS65_LH_MX41X7 port map( D0 => registers_20_12_port, S0 => n2613, D1
                           => registers_21_12_port, S1 => n2610, D2 => 
                           registers_22_12_port, S2 => n2607, D3 => 
                           registers_23_12_port, S3 => n2604, Z => n796);
   U1154 : HS65_LH_MX41X7 port map( D0 => registers_4_12_port, S0 => n2661, D1 
                           => registers_5_12_port, S1 => n2658, D2 => 
                           registers_6_12_port, S2 => n2655, D3 => 
                           registers_7_12_port, S3 => n2652, Z => n790);
   U1155 : HS65_LH_MX41X7 port map( D0 => registers_20_13_port, S0 => n2613, D1
                           => registers_21_13_port, S1 => n2610, D2 => 
                           registers_22_13_port, S2 => n2607, D3 => 
                           registers_23_13_port, S3 => n2604, Z => n781);
   U1156 : HS65_LH_MX41X7 port map( D0 => registers_4_13_port, S0 => n2661, D1 
                           => registers_5_13_port, S1 => n2658, D2 => 
                           registers_6_13_port, S2 => n2655, D3 => 
                           registers_7_13_port, S3 => n2652, Z => n775);
   U1157 : HS65_LH_MX41X7 port map( D0 => registers_20_14_port, S0 => n2613, D1
                           => registers_21_14_port, S1 => n2610, D2 => 
                           registers_22_14_port, S2 => n2607, D3 => 
                           registers_23_14_port, S3 => n2604, Z => n766);
   U1158 : HS65_LH_MX41X7 port map( D0 => registers_4_14_port, S0 => n2661, D1 
                           => registers_5_14_port, S1 => n2658, D2 => 
                           registers_6_14_port, S2 => n2655, D3 => 
                           registers_7_14_port, S3 => n2652, Z => n760);
   U1159 : HS65_LH_MX41X7 port map( D0 => registers_20_15_port, S0 => n2613, D1
                           => registers_21_15_port, S1 => n2610, D2 => 
                           registers_22_15_port, S2 => n2607, D3 => 
                           registers_23_15_port, S3 => n2604, Z => n751);
   U1160 : HS65_LH_MX41X7 port map( D0 => registers_4_15_port, S0 => n2661, D1 
                           => registers_5_15_port, S1 => n2658, D2 => 
                           registers_6_15_port, S2 => n2655, D3 => 
                           registers_7_15_port, S3 => n2652, Z => n745);
   U1161 : HS65_LH_MX41X7 port map( D0 => registers_20_16_port, S0 => n2613, D1
                           => registers_21_16_port, S1 => n2610, D2 => 
                           registers_22_16_port, S2 => n2607, D3 => 
                           registers_23_16_port, S3 => n2604, Z => n736);
   U1162 : HS65_LH_MX41X7 port map( D0 => registers_4_16_port, S0 => n2661, D1 
                           => registers_5_16_port, S1 => n2658, D2 => 
                           registers_6_16_port, S2 => n2655, D3 => 
                           registers_7_16_port, S3 => n2652, Z => n730);
   U1163 : HS65_LH_MX41X7 port map( D0 => registers_20_17_port, S0 => n2613, D1
                           => registers_21_17_port, S1 => n2610, D2 => 
                           registers_22_17_port, S2 => n2607, D3 => 
                           registers_23_17_port, S3 => n2604, Z => n721);
   U1164 : HS65_LH_MX41X7 port map( D0 => registers_4_17_port, S0 => n2661, D1 
                           => registers_5_17_port, S1 => n2658, D2 => 
                           registers_6_17_port, S2 => n2655, D3 => 
                           registers_7_17_port, S3 => n2652, Z => n715);
   U1165 : HS65_LH_MX41X7 port map( D0 => registers_20_18_port, S0 => n2613, D1
                           => registers_21_18_port, S1 => n2610, D2 => 
                           registers_22_18_port, S2 => n2607, D3 => 
                           registers_23_18_port, S3 => n2604, Z => n706);
   U1166 : HS65_LH_MX41X7 port map( D0 => registers_4_18_port, S0 => n2661, D1 
                           => registers_5_18_port, S1 => n2658, D2 => 
                           registers_6_18_port, S2 => n2655, D3 => 
                           registers_7_18_port, S3 => n2652, Z => n700);
   U1167 : HS65_LH_MX41X7 port map( D0 => registers_20_19_port, S0 => n2613, D1
                           => registers_21_19_port, S1 => n2610, D2 => 
                           registers_22_19_port, S2 => n2607, D3 => 
                           registers_23_19_port, S3 => n2604, Z => n691);
   U1168 : HS65_LH_MX41X7 port map( D0 => registers_4_19_port, S0 => n2661, D1 
                           => registers_5_19_port, S1 => n2658, D2 => 
                           registers_6_19_port, S2 => n2655, D3 => 
                           registers_7_19_port, S3 => n2652, Z => n685);
   U1169 : HS65_LH_MX41X7 port map( D0 => registers_20_20_port, S0 => n2614, D1
                           => registers_21_20_port, S1 => n2611, D2 => 
                           registers_22_20_port, S2 => n2608, D3 => 
                           registers_23_20_port, S3 => n2605, Z => n661);
   U1170 : HS65_LH_MX41X7 port map( D0 => registers_4_20_port, S0 => n2662, D1 
                           => registers_5_20_port, S1 => n2659, D2 => 
                           registers_6_20_port, S2 => n2656, D3 => 
                           registers_7_20_port, S3 => n2653, Z => n655);
   U1171 : HS65_LH_MX41X7 port map( D0 => registers_20_21_port, S0 => n2614, D1
                           => registers_21_21_port, S1 => n2611, D2 => 
                           registers_22_21_port, S2 => n2608, D3 => 
                           registers_23_21_port, S3 => n2605, Z => n646);
   U1172 : HS65_LH_MX41X7 port map( D0 => registers_4_21_port, S0 => n2662, D1 
                           => registers_5_21_port, S1 => n2659, D2 => 
                           registers_6_21_port, S2 => n2656, D3 => 
                           registers_7_21_port, S3 => n2653, Z => n640);
   U1173 : HS65_LH_MX41X7 port map( D0 => registers_20_22_port, S0 => n2614, D1
                           => registers_21_22_port, S1 => n2611, D2 => 
                           registers_22_22_port, S2 => n2608, D3 => 
                           registers_23_22_port, S3 => n2605, Z => n631);
   U1174 : HS65_LH_MX41X7 port map( D0 => registers_4_22_port, S0 => n2662, D1 
                           => registers_5_22_port, S1 => n2659, D2 => 
                           registers_6_22_port, S2 => n2656, D3 => 
                           registers_7_22_port, S3 => n2653, Z => n625);
   U1175 : HS65_LH_MX41X7 port map( D0 => registers_20_23_port, S0 => n2614, D1
                           => registers_21_23_port, S1 => n2611, D2 => 
                           registers_22_23_port, S2 => n2608, D3 => 
                           registers_23_23_port, S3 => n2605, Z => n616);
   U1176 : HS65_LH_MX41X7 port map( D0 => registers_4_23_port, S0 => n2662, D1 
                           => registers_5_23_port, S1 => n2659, D2 => 
                           registers_6_23_port, S2 => n2656, D3 => 
                           registers_7_23_port, S3 => n2653, Z => n610);
   U1177 : HS65_LH_MX41X7 port map( D0 => registers_20_24_port, S0 => n2614, D1
                           => registers_21_24_port, S1 => n2611, D2 => 
                           registers_22_24_port, S2 => n2608, D3 => 
                           registers_23_24_port, S3 => n2605, Z => n601);
   U1178 : HS65_LH_MX41X7 port map( D0 => registers_4_24_port, S0 => n2662, D1 
                           => registers_5_24_port, S1 => n2659, D2 => 
                           registers_6_24_port, S2 => n2656, D3 => 
                           registers_7_24_port, S3 => n2653, Z => n595);
   U1179 : HS65_LH_MX41X7 port map( D0 => registers_20_25_port, S0 => n2614, D1
                           => registers_21_25_port, S1 => n2611, D2 => 
                           registers_22_25_port, S2 => n2608, D3 => 
                           registers_23_25_port, S3 => n2605, Z => n586);
   U1180 : HS65_LH_MX41X7 port map( D0 => registers_4_25_port, S0 => n2662, D1 
                           => registers_5_25_port, S1 => n2659, D2 => 
                           registers_6_25_port, S2 => n2656, D3 => 
                           registers_7_25_port, S3 => n2653, Z => n580);
   U1181 : HS65_LH_MX41X7 port map( D0 => registers_20_26_port, S0 => n2614, D1
                           => registers_21_26_port, S1 => n2611, D2 => 
                           registers_22_26_port, S2 => n2608, D3 => 
                           registers_23_26_port, S3 => n2605, Z => n571);
   U1182 : HS65_LH_MX41X7 port map( D0 => registers_4_26_port, S0 => n2662, D1 
                           => registers_5_26_port, S1 => n2659, D2 => 
                           registers_6_26_port, S2 => n2656, D3 => 
                           registers_7_26_port, S3 => n2653, Z => n565);
   U1183 : HS65_LH_MX41X7 port map( D0 => registers_20_27_port, S0 => n2614, D1
                           => registers_21_27_port, S1 => n2611, D2 => 
                           registers_22_27_port, S2 => n2608, D3 => 
                           registers_23_27_port, S3 => n2605, Z => n556);
   U1184 : HS65_LH_MX41X7 port map( D0 => registers_4_27_port, S0 => n2662, D1 
                           => registers_5_27_port, S1 => n2659, D2 => 
                           registers_6_27_port, S2 => n2656, D3 => 
                           registers_7_27_port, S3 => n2653, Z => n550);
   U1185 : HS65_LH_MX41X7 port map( D0 => registers_20_28_port, S0 => n2614, D1
                           => registers_21_28_port, S1 => n2611, D2 => 
                           registers_22_28_port, S2 => n2608, D3 => 
                           registers_23_28_port, S3 => n2605, Z => n541);
   U1186 : HS65_LH_MX41X7 port map( D0 => registers_4_28_port, S0 => n2662, D1 
                           => registers_5_28_port, S1 => n2659, D2 => 
                           registers_6_28_port, S2 => n2656, D3 => 
                           registers_7_28_port, S3 => n2653, Z => n535);
   U1187 : HS65_LH_MX41X7 port map( D0 => registers_20_29_port, S0 => n2614, D1
                           => registers_21_29_port, S1 => n2611, D2 => 
                           registers_22_29_port, S2 => n2608, D3 => 
                           registers_23_29_port, S3 => n2605, Z => n526);
   U1188 : HS65_LH_MX41X7 port map( D0 => registers_4_29_port, S0 => n2662, D1 
                           => registers_5_29_port, S1 => n2659, D2 => 
                           registers_6_29_port, S2 => n2656, D3 => 
                           registers_7_29_port, S3 => n2653, Z => n520);
   U1189 : HS65_LH_MX41X7 port map( D0 => registers_20_30_port, S0 => n2614, D1
                           => registers_21_30_port, S1 => n2611, D2 => 
                           registers_22_30_port, S2 => n2608, D3 => 
                           registers_23_30_port, S3 => n2605, Z => n496);
   U1190 : HS65_LH_MX41X7 port map( D0 => registers_4_30_port, S0 => n2662, D1 
                           => registers_5_30_port, S1 => n2659, D2 => 
                           registers_6_30_port, S2 => n2656, D3 => 
                           registers_7_30_port, S3 => n2653, Z => n490);
   U1191 : HS65_LH_MX41X7 port map( D0 => registers_20_31_port, S0 => n2615, D1
                           => registers_21_31_port, S1 => n2612, D2 => 
                           registers_22_31_port, S2 => n2609, D3 => 
                           registers_23_31_port, S3 => n2606, Z => n481);
   U1192 : HS65_LH_MX41X7 port map( D0 => registers_4_31_port, S0 => n2663, D1 
                           => registers_5_31_port, S1 => n2660, D2 => 
                           registers_6_31_port, S2 => n2657, D3 => 
                           registers_7_31_port, S3 => n2654, Z => n475);
   U1193 : HS65_LH_IVX9 port map( A => regfile_i(40), Z => n2898);
   U1194 : HS65_LH_IVX9 port map( A => regfile_i(45), Z => n2903);
   U1195 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_0_port, D1 
                           => n2517, S1 => registers_21_0_port, D2 => n2514, S2
                           => registers_22_0_port, D3 => n2511, S3 => 
                           registers_23_0_port, Z => n1379);
   U1196 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_0_port, D1 
                           => n2565, S1 => registers_5_0_port, D2 => n2562, S2 
                           => registers_6_0_port, D3 => n2559, S3 => 
                           registers_7_0_port, Z => n1363);
   U1197 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_1_port, D1 
                           => n2517, S1 => registers_21_1_port, D2 => n2514, S2
                           => registers_22_1_port, D3 => n2511, S3 => 
                           registers_23_1_port, Z => n1204);
   U1198 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_1_port, D1 
                           => n2565, S1 => registers_5_1_port, D2 => n2562, S2 
                           => registers_6_1_port, D3 => n2559, S3 => 
                           registers_7_1_port, Z => n1198);
   U1199 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_2_port, D1 
                           => n2518, S1 => registers_21_2_port, D2 => n2515, S2
                           => registers_22_2_port, D3 => n2512, S3 => 
                           registers_23_2_port, Z => n1039);
   U1200 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_2_port, D1 
                           => n2566, S1 => registers_5_2_port, D2 => n2563, S2 
                           => registers_6_2_port, D3 => n2560, S3 => 
                           registers_7_2_port, Z => n1033);
   U1201 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_3_port, D1 
                           => n2519, S1 => registers_21_3_port, D2 => n2515, S2
                           => registers_22_3_port, D3 => n2513, S3 => 
                           registers_23_3_port, Z => n994);
   U1202 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_3_port, D1 
                           => n2567, S1 => registers_5_3_port, D2 => n2563, S2 
                           => registers_6_3_port, D3 => n2561, S3 => 
                           registers_7_3_port, Z => n988);
   U1203 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_4_port, D1 
                           => n2519, S1 => registers_21_4_port, D2 => n2516, S2
                           => registers_22_4_port, D3 => n2513, S3 => 
                           registers_23_4_port, Z => n979);
   U1204 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_4_port, D1 
                           => n2567, S1 => registers_5_4_port, D2 => n2564, S2 
                           => registers_6_4_port, D3 => n2561, S3 => 
                           registers_7_4_port, Z => n973);
   U1205 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_5_port, D1 
                           => n2519, S1 => registers_21_5_port, D2 => n2516, S2
                           => registers_22_5_port, D3 => n2513, S3 => 
                           registers_23_5_port, Z => n964);
   U1206 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_5_port, D1 
                           => n2567, S1 => registers_5_5_port, D2 => n2564, S2 
                           => registers_6_5_port, D3 => n2561, S3 => 
                           registers_7_5_port, Z => n958);
   U1207 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_6_port, D1 
                           => n2519, S1 => registers_21_6_port, D2 => n2516, S2
                           => registers_22_6_port, D3 => n2513, S3 => 
                           registers_23_6_port, Z => n949);
   U1208 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_6_port, D1 
                           => n2567, S1 => registers_5_6_port, D2 => n2564, S2 
                           => registers_6_6_port, D3 => n2561, S3 => 
                           registers_7_6_port, Z => n943);
   U1209 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_7_port, D1 
                           => n2519, S1 => registers_21_7_port, D2 => n2516, S2
                           => registers_22_7_port, D3 => n2513, S3 => 
                           registers_23_7_port, Z => n934);
   U1210 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_7_port, D1 
                           => n2567, S1 => registers_5_7_port, D2 => n2564, S2 
                           => registers_6_7_port, D3 => n2561, S3 => 
                           registers_7_7_port, Z => n928);
   U1211 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_8_port, D1 
                           => n2519, S1 => registers_21_8_port, D2 => n2516, S2
                           => registers_22_8_port, D3 => n2513, S3 => 
                           registers_23_8_port, Z => n919);
   U1212 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_8_port, D1 
                           => n2567, S1 => registers_5_8_port, D2 => n2564, S2 
                           => registers_6_8_port, D3 => n2561, S3 => 
                           registers_7_8_port, Z => n913);
   U1213 : HS65_LH_MX41X7 port map( D0 => n2522, S0 => registers_20_9_port, D1 
                           => n2519, S1 => registers_21_9_port, D2 => n2516, S2
                           => registers_22_9_port, D3 => n2513, S3 => 
                           registers_23_9_port, Z => n888);
   U1214 : HS65_LH_MX41X7 port map( D0 => n2570, S0 => registers_4_9_port, D1 
                           => n2567, S1 => registers_5_9_port, D2 => n2564, S2 
                           => registers_6_9_port, D3 => n2561, S3 => 
                           registers_7_9_port, Z => n866);
   U1215 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_10_port, D1
                           => n2517, S1 => registers_21_10_port, D2 => n2514, 
                           S2 => registers_22_10_port, D3 => n2511, S3 => 
                           registers_23_10_port, Z => n1354);
   U1216 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_10_port, D1 
                           => n2565, S1 => registers_5_10_port, D2 => n2562, S2
                           => registers_6_10_port, D3 => n2559, S3 => 
                           registers_7_10_port, Z => n1348);
   U1217 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_11_port, D1
                           => n2517, S1 => registers_21_11_port, D2 => n2514, 
                           S2 => registers_22_11_port, D3 => n2511, S3 => 
                           registers_23_11_port, Z => n1339);
   U1218 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_11_port, D1 
                           => n2565, S1 => registers_5_11_port, D2 => n2562, S2
                           => registers_6_11_port, D3 => n2559, S3 => 
                           registers_7_11_port, Z => n1333);
   U1219 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_12_port, D1
                           => n2517, S1 => registers_21_12_port, D2 => n2514, 
                           S2 => registers_22_12_port, D3 => n2511, S3 => 
                           registers_23_12_port, Z => n1324);
   U1220 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_12_port, D1 
                           => n2565, S1 => registers_5_12_port, D2 => n2562, S2
                           => registers_6_12_port, D3 => n2559, S3 => 
                           registers_7_12_port, Z => n1318);
   U1221 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_13_port, D1
                           => n2517, S1 => registers_21_13_port, D2 => n2514, 
                           S2 => registers_22_13_port, D3 => n2511, S3 => 
                           registers_23_13_port, Z => n1309);
   U1222 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_13_port, D1 
                           => n2565, S1 => registers_5_13_port, D2 => n2562, S2
                           => registers_6_13_port, D3 => n2559, S3 => 
                           registers_7_13_port, Z => n1303);
   U1223 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_14_port, D1
                           => n2517, S1 => registers_21_14_port, D2 => n2514, 
                           S2 => registers_22_14_port, D3 => n2511, S3 => 
                           registers_23_14_port, Z => n1294);
   U1224 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_14_port, D1 
                           => n2565, S1 => registers_5_14_port, D2 => n2562, S2
                           => registers_6_14_port, D3 => n2559, S3 => 
                           registers_7_14_port, Z => n1288);
   U1225 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_15_port, D1
                           => n2517, S1 => registers_21_15_port, D2 => n2514, 
                           S2 => registers_22_15_port, D3 => n2511, S3 => 
                           registers_23_15_port, Z => n1279);
   U1226 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_15_port, D1 
                           => n2565, S1 => registers_5_15_port, D2 => n2562, S2
                           => registers_6_15_port, D3 => n2559, S3 => 
                           registers_7_15_port, Z => n1273);
   U1227 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_16_port, D1
                           => n2517, S1 => registers_21_16_port, D2 => n2514, 
                           S2 => registers_22_16_port, D3 => n2511, S3 => 
                           registers_23_16_port, Z => n1264);
   U1228 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_16_port, D1 
                           => n2565, S1 => registers_5_16_port, D2 => n2562, S2
                           => registers_6_16_port, D3 => n2559, S3 => 
                           registers_7_16_port, Z => n1258);
   U1229 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_17_port, D1
                           => n2517, S1 => registers_21_17_port, D2 => n2514, 
                           S2 => registers_22_17_port, D3 => n2511, S3 => 
                           registers_23_17_port, Z => n1249);
   U1230 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_17_port, D1 
                           => n2565, S1 => registers_5_17_port, D2 => n2562, S2
                           => registers_6_17_port, D3 => n2559, S3 => 
                           registers_7_17_port, Z => n1243);
   U1231 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_18_port, D1
                           => n2517, S1 => registers_21_18_port, D2 => n2514, 
                           S2 => registers_22_18_port, D3 => n2511, S3 => 
                           registers_23_18_port, Z => n1234);
   U1232 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_18_port, D1 
                           => n2565, S1 => registers_5_18_port, D2 => n2562, S2
                           => registers_6_18_port, D3 => n2559, S3 => 
                           registers_7_18_port, Z => n1228);
   U1233 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_19_port, D1
                           => n2517, S1 => registers_21_19_port, D2 => n2514, 
                           S2 => registers_22_19_port, D3 => n2511, S3 => 
                           registers_23_19_port, Z => n1219);
   U1234 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_19_port, D1 
                           => n2565, S1 => registers_5_19_port, D2 => n2562, S2
                           => registers_6_19_port, D3 => n2559, S3 => 
                           registers_7_19_port, Z => n1213);
   U1235 : HS65_LH_MX41X7 port map( D0 => n2520, S0 => registers_20_20_port, D1
                           => n2518, S1 => registers_21_20_port, D2 => n2514, 
                           S2 => registers_22_20_port, D3 => n2512, S3 => 
                           registers_23_20_port, Z => n1189);
   U1236 : HS65_LH_MX41X7 port map( D0 => n2568, S0 => registers_4_20_port, D1 
                           => n2566, S1 => registers_5_20_port, D2 => n2562, S2
                           => registers_6_20_port, D3 => n2560, S3 => 
                           registers_7_20_port, Z => n1183);
   U1237 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_21_port, D1
                           => n2518, S1 => registers_21_21_port, D2 => n2515, 
                           S2 => registers_22_21_port, D3 => n2512, S3 => 
                           registers_23_21_port, Z => n1174);
   U1238 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_21_port, D1 
                           => n2566, S1 => registers_5_21_port, D2 => n2563, S2
                           => registers_6_21_port, D3 => n2560, S3 => 
                           registers_7_21_port, Z => n1168);
   U1239 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_22_port, D1
                           => n2518, S1 => registers_21_22_port, D2 => n2515, 
                           S2 => registers_22_22_port, D3 => n2512, S3 => 
                           registers_23_22_port, Z => n1159);
   U1240 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_22_port, D1 
                           => n2566, S1 => registers_5_22_port, D2 => n2563, S2
                           => registers_6_22_port, D3 => n2560, S3 => 
                           registers_7_22_port, Z => n1153);
   U1241 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_23_port, D1
                           => n2518, S1 => registers_21_23_port, D2 => n2515, 
                           S2 => registers_22_23_port, D3 => n2512, S3 => 
                           registers_23_23_port, Z => n1144);
   U1242 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_23_port, D1 
                           => n2566, S1 => registers_5_23_port, D2 => n2563, S2
                           => registers_6_23_port, D3 => n2560, S3 => 
                           registers_7_23_port, Z => n1138);
   U1243 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_24_port, D1
                           => n2518, S1 => registers_21_24_port, D2 => n2515, 
                           S2 => registers_22_24_port, D3 => n2512, S3 => 
                           registers_23_24_port, Z => n1129);
   U1244 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_24_port, D1 
                           => n2566, S1 => registers_5_24_port, D2 => n2563, S2
                           => registers_6_24_port, D3 => n2560, S3 => 
                           registers_7_24_port, Z => n1123);
   U1245 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_25_port, D1
                           => n2518, S1 => registers_21_25_port, D2 => n2515, 
                           S2 => registers_22_25_port, D3 => n2512, S3 => 
                           registers_23_25_port, Z => n1114);
   U1246 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_25_port, D1 
                           => n2566, S1 => registers_5_25_port, D2 => n2563, S2
                           => registers_6_25_port, D3 => n2560, S3 => 
                           registers_7_25_port, Z => n1108);
   U1247 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_26_port, D1
                           => n2518, S1 => registers_21_26_port, D2 => n2515, 
                           S2 => registers_22_26_port, D3 => n2512, S3 => 
                           registers_23_26_port, Z => n1099);
   U1248 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_26_port, D1 
                           => n2566, S1 => registers_5_26_port, D2 => n2563, S2
                           => registers_6_26_port, D3 => n2560, S3 => 
                           registers_7_26_port, Z => n1093);
   U1249 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_27_port, D1
                           => n2518, S1 => registers_21_27_port, D2 => n2515, 
                           S2 => registers_22_27_port, D3 => n2512, S3 => 
                           registers_23_27_port, Z => n1084);
   U1250 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_27_port, D1 
                           => n2566, S1 => registers_5_27_port, D2 => n2563, S2
                           => registers_6_27_port, D3 => n2560, S3 => 
                           registers_7_27_port, Z => n1078);
   U1251 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_28_port, D1
                           => n2518, S1 => registers_21_28_port, D2 => n2515, 
                           S2 => registers_22_28_port, D3 => n2512, S3 => 
                           registers_23_28_port, Z => n1069);
   U1252 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_28_port, D1 
                           => n2566, S1 => registers_5_28_port, D2 => n2563, S2
                           => registers_6_28_port, D3 => n2560, S3 => 
                           registers_7_28_port, Z => n1063);
   U1253 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_29_port, D1
                           => n2518, S1 => registers_21_29_port, D2 => n2515, 
                           S2 => registers_22_29_port, D3 => n2512, S3 => 
                           registers_23_29_port, Z => n1054);
   U1254 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_29_port, D1 
                           => n2566, S1 => registers_5_29_port, D2 => n2563, S2
                           => registers_6_29_port, D3 => n2560, S3 => 
                           registers_7_29_port, Z => n1048);
   U1255 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_30_port, D1
                           => n2518, S1 => registers_21_30_port, D2 => n2515, 
                           S2 => registers_22_30_port, D3 => n2512, S3 => 
                           registers_23_30_port, Z => n1024);
   U1256 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_30_port, D1 
                           => n2566, S1 => registers_5_30_port, D2 => n2563, S2
                           => registers_6_30_port, D3 => n2560, S3 => 
                           registers_7_30_port, Z => n1018);
   U1257 : HS65_LH_MX41X7 port map( D0 => n2521, S0 => registers_20_31_port, D1
                           => n2519, S1 => registers_21_31_port, D2 => n2515, 
                           S2 => registers_22_31_port, D3 => n2513, S3 => 
                           registers_23_31_port, Z => n1009);
   U1258 : HS65_LH_MX41X7 port map( D0 => n2569, S0 => registers_4_31_port, D1 
                           => n2567, S1 => registers_5_31_port, D2 => n2563, S2
                           => registers_6_31_port, D3 => n2561, S3 => 
                           registers_7_31_port, Z => n1003);
   U1259 : HS65_LH_IVX9 port map( A => regfile_i(44), Z => n2902);
   U1260 : HS65_LH_IVX9 port map( A => regfile_i(49), Z => n2907);
   U1261 : HS65_LH_IVX9 port map( A => regfile_i(42), Z => n2900);
   U1262 : HS65_LH_IVX9 port map( A => regfile_i(47), Z => n2905);
   U1263 : HS65_LH_IVX9 port map( A => regfile_i(43), Z => n2901);
   U1264 : HS65_LH_IVX9 port map( A => regfile_i(48), Z => n2906);
   U1265 : HS65_LH_IVX9 port map( A => regfile_i(41), Z => n2899);
   U1266 : HS65_LH_IVX9 port map( A => regfile_i(46), Z => n2904);
   U1267 : HS65_LH_OAI21X3 port map( A => n2698, B => n280, C => n1360, Z => 
                           regfile_o(32));
   U1268 : HS65_LH_OAI21X3 port map( A => n1361, B => n1362, C => n278, Z => 
                           n1360);
   U1269 : HS65_LH_NAND4ABX3 port map( A => n1363, B => n1364, C => n1365, D =>
                           n1366, Z => n1362);
   U1270 : HS65_LH_OAI21X3 port map( A => n2700, B => n282, C => n1195, Z => 
                           regfile_o(33));
   U1271 : HS65_LH_OAI21X3 port map( A => n1196, B => n1197, C => n279, Z => 
                           n1195);
   U1272 : HS65_LH_NAND4ABX3 port map( A => n1198, B => n1199, C => n1200, D =>
                           n1201, Z => n1197);
   U1273 : HS65_LH_OAI21X3 port map( A => n2702, B => n281, C => n1030, Z => 
                           regfile_o(34));
   U1274 : HS65_LH_OAI21X3 port map( A => n1031, B => n1032, C => n280, Z => 
                           n1030);
   U1275 : HS65_LH_NAND4ABX3 port map( A => n1033, B => n1034, C => n1035, D =>
                           n1036, Z => n1032);
   U1276 : HS65_LH_OAI21X3 port map( A => n2704, B => n280, C => n985, Z => 
                           regfile_o(35));
   U1277 : HS65_LH_OAI21X3 port map( A => n986, B => n987, C => n279, Z => n985
                           );
   U1278 : HS65_LH_NAND4ABX3 port map( A => n988, B => n989, C => n990, D => 
                           n991, Z => n987);
   U1279 : HS65_LH_OAI21X3 port map( A => n2706, B => n281, C => n970, Z => 
                           regfile_o(36));
   U1280 : HS65_LH_OAI21X3 port map( A => n971, B => n972, C => n279, Z => n970
                           );
   U1281 : HS65_LH_NAND4ABX3 port map( A => n973, B => n974, C => n975, D => 
                           n976, Z => n972);
   U1282 : HS65_LH_OAI21X3 port map( A => n2708, B => n280, C => n955, Z => 
                           regfile_o(37));
   U1283 : HS65_LH_OAI21X3 port map( A => n956, B => n957, C => n279, Z => n955
                           );
   U1284 : HS65_LH_NAND4ABX3 port map( A => n958, B => n959, C => n960, D => 
                           n961, Z => n957);
   U1285 : HS65_LH_OAI21X3 port map( A => n2710, B => n280, C => n940, Z => 
                           regfile_o(38));
   U1286 : HS65_LH_OAI21X3 port map( A => n941, B => n942, C => n278, Z => n940
                           );
   U1287 : HS65_LH_NAND4ABX3 port map( A => n943, B => n944, C => n945, D => 
                           n946, Z => n942);
   U1288 : HS65_LH_OAI21X3 port map( A => n2712, B => n281, C => n925, Z => 
                           regfile_o(39));
   U1289 : HS65_LH_OAI21X3 port map( A => n926, B => n927, C => n278, Z => n925
                           );
   U1290 : HS65_LH_NAND4ABX3 port map( A => n928, B => n929, C => n930, D => 
                           n931, Z => n927);
   U1291 : HS65_LH_OAI21X3 port map( A => n2714, B => n280, C => n910, Z => 
                           regfile_o(40));
   U1292 : HS65_LH_OAI21X3 port map( A => n911, B => n912, C => n278, Z => n910
                           );
   U1293 : HS65_LH_NAND4ABX3 port map( A => n913, B => n914, C => n915, D => 
                           n916, Z => n912);
   U1294 : HS65_LH_OAI21X3 port map( A => n2716, B => n281, C => n863, Z => 
                           regfile_o(41));
   U1295 : HS65_LH_OAI21X3 port map( A => n864, B => n865, C => n278, Z => n863
                           );
   U1296 : HS65_LH_NAND4ABX3 port map( A => n866, B => n867, C => n868, D => 
                           n869, Z => n865);
   U1297 : HS65_LH_OAI21X3 port map( A => n2718, B => n282, C => n1345, Z => 
                           regfile_o(42));
   U1298 : HS65_LH_OAI21X3 port map( A => n1346, B => n1347, C => n278, Z => 
                           n1345);
   U1299 : HS65_LH_NAND4ABX3 port map( A => n1348, B => n1349, C => n1350, D =>
                           n1351, Z => n1347);
   U1300 : HS65_LH_OAI21X3 port map( A => n2720, B => n282, C => n1330, Z => 
                           regfile_o(43));
   U1301 : HS65_LH_OAI21X3 port map( A => n1331, B => n1332, C => n278, Z => 
                           n1330);
   U1302 : HS65_LH_NAND4ABX3 port map( A => n1333, B => n1334, C => n1335, D =>
                           n1336, Z => n1332);
   U1303 : HS65_LH_OAI21X3 port map( A => n2722, B => n282, C => n1315, Z => 
                           regfile_o(44));
   U1304 : HS65_LH_OAI21X3 port map( A => n1316, B => n1317, C => n278, Z => 
                           n1315);
   U1305 : HS65_LH_NAND4ABX3 port map( A => n1318, B => n1319, C => n1320, D =>
                           n1321, Z => n1317);
   U1306 : HS65_LH_OAI21X3 port map( A => n2724, B => n282, C => n1300, Z => 
                           regfile_o(45));
   U1307 : HS65_LH_OAI21X3 port map( A => n1301, B => n1302, C => n278, Z => 
                           n1300);
   U1308 : HS65_LH_NAND4ABX3 port map( A => n1303, B => n1304, C => n1305, D =>
                           n1306, Z => n1302);
   U1309 : HS65_LH_OAI21X3 port map( A => n2726, B => n282, C => n1285, Z => 
                           regfile_o(46));
   U1310 : HS65_LH_OAI21X3 port map( A => n1286, B => n1287, C => n278, Z => 
                           n1285);
   U1311 : HS65_LH_NAND4ABX3 port map( A => n1288, B => n1289, C => n1290, D =>
                           n1291, Z => n1287);
   U1312 : HS65_LH_OAI21X3 port map( A => n2728, B => n282, C => n1270, Z => 
                           regfile_o(47));
   U1313 : HS65_LH_OAI21X3 port map( A => n1271, B => n1272, C => n278, Z => 
                           n1270);
   U1314 : HS65_LH_NAND4ABX3 port map( A => n1273, B => n1274, C => n1275, D =>
                           n1276, Z => n1272);
   U1315 : HS65_LH_OAI21X3 port map( A => n2730, B => n282, C => n1255, Z => 
                           regfile_o(48));
   U1316 : HS65_LH_OAI21X3 port map( A => n1256, B => n1257, C => n278, Z => 
                           n1255);
   U1317 : HS65_LH_NAND4ABX3 port map( A => n1258, B => n1259, C => n1260, D =>
                           n1261, Z => n1257);
   U1318 : HS65_LH_OAI21X3 port map( A => n2732, B => n282, C => n1240, Z => 
                           regfile_o(49));
   U1319 : HS65_LH_OAI21X3 port map( A => n1241, B => n1242, C => n279, Z => 
                           n1240);
   U1320 : HS65_LH_NAND4ABX3 port map( A => n1243, B => n1244, C => n1245, D =>
                           n1246, Z => n1242);
   U1321 : HS65_LH_OAI21X3 port map( A => n2734, B => n282, C => n1225, Z => 
                           regfile_o(50));
   U1322 : HS65_LH_OAI21X3 port map( A => n1226, B => n1227, C => n279, Z => 
                           n1225);
   U1323 : HS65_LH_NAND4ABX3 port map( A => n1228, B => n1229, C => n1230, D =>
                           n1231, Z => n1227);
   U1324 : HS65_LH_OAI21X3 port map( A => n2736, B => n282, C => n1210, Z => 
                           regfile_o(51));
   U1325 : HS65_LH_OAI21X3 port map( A => n1211, B => n1212, C => n279, Z => 
                           n1210);
   U1326 : HS65_LH_NAND4ABX3 port map( A => n1213, B => n1214, C => n1215, D =>
                           n1216, Z => n1212);
   U1327 : HS65_LH_OAI21X3 port map( A => n2738, B => n282, C => n1180, Z => 
                           regfile_o(52));
   U1328 : HS65_LH_OAI21X3 port map( A => n1181, B => n1182, C => n279, Z => 
                           n1180);
   U1329 : HS65_LH_NAND4ABX3 port map( A => n1183, B => n1184, C => n1185, D =>
                           n1186, Z => n1182);
   U1330 : HS65_LH_OAI21X3 port map( A => n2740, B => n282, C => n1165, Z => 
                           regfile_o(53));
   U1331 : HS65_LH_OAI21X3 port map( A => n1166, B => n1167, C => n279, Z => 
                           n1165);
   U1332 : HS65_LH_NAND4ABX3 port map( A => n1168, B => n1169, C => n1170, D =>
                           n1171, Z => n1167);
   U1333 : HS65_LH_OAI21X3 port map( A => n2742, B => n281, C => n1150, Z => 
                           regfile_o(54));
   U1334 : HS65_LH_OAI21X3 port map( A => n1151, B => n1152, C => n279, Z => 
                           n1150);
   U1335 : HS65_LH_NAND4ABX3 port map( A => n1153, B => n1154, C => n1155, D =>
                           n1156, Z => n1152);
   U1336 : HS65_LH_OAI21X3 port map( A => n2744, B => n281, C => n1135, Z => 
                           regfile_o(55));
   U1337 : HS65_LH_OAI21X3 port map( A => n1136, B => n1137, C => n279, Z => 
                           n1135);
   U1338 : HS65_LH_NAND4ABX3 port map( A => n1138, B => n1139, C => n1140, D =>
                           n1141, Z => n1137);
   U1339 : HS65_LH_OAI21X3 port map( A => n2746, B => n281, C => n1120, Z => 
                           regfile_o(56));
   U1340 : HS65_LH_OAI21X3 port map( A => n1121, B => n1122, C => n280, Z => 
                           n1120);
   U1341 : HS65_LH_NAND4ABX3 port map( A => n1123, B => n1124, C => n1125, D =>
                           n1126, Z => n1122);
   U1342 : HS65_LH_OAI21X3 port map( A => n2748, B => n281, C => n1105, Z => 
                           regfile_o(57));
   U1343 : HS65_LH_OAI21X3 port map( A => n1106, B => n1107, C => n280, Z => 
                           n1105);
   U1344 : HS65_LH_NAND4ABX3 port map( A => n1108, B => n1109, C => n1110, D =>
                           n1111, Z => n1107);
   U1345 : HS65_LH_OAI21X3 port map( A => n2750, B => n281, C => n1090, Z => 
                           regfile_o(58));
   U1346 : HS65_LH_OAI21X3 port map( A => n1091, B => n1092, C => n279, Z => 
                           n1090);
   U1347 : HS65_LH_NAND4ABX3 port map( A => n1093, B => n1094, C => n1095, D =>
                           n1096, Z => n1092);
   U1348 : HS65_LH_OAI21X3 port map( A => n2752, B => n281, C => n1075, Z => 
                           regfile_o(59));
   U1349 : HS65_LH_OAI21X3 port map( A => n1076, B => n1077, C => n280, Z => 
                           n1075);
   U1350 : HS65_LH_NAND4ABX3 port map( A => n1078, B => n1079, C => n1080, D =>
                           n1081, Z => n1077);
   U1351 : HS65_LH_OAI21X3 port map( A => n2754, B => n281, C => n1060, Z => 
                           regfile_o(60));
   U1352 : HS65_LH_OAI21X3 port map( A => n1061, B => n1062, C => n280, Z => 
                           n1060);
   U1353 : HS65_LH_NAND4ABX3 port map( A => n1063, B => n1064, C => n1065, D =>
                           n1066, Z => n1062);
   U1354 : HS65_LH_OAI21X3 port map( A => n2756, B => n281, C => n1045, Z => 
                           regfile_o(61));
   U1355 : HS65_LH_OAI21X3 port map( A => n1046, B => n1047, C => n280, Z => 
                           n1045);
   U1356 : HS65_LH_NAND4ABX3 port map( A => n1048, B => n1049, C => n1050, D =>
                           n1051, Z => n1047);
   U1357 : HS65_LH_OAI21X3 port map( A => n2758, B => n281, C => n1015, Z => 
                           regfile_o(62));
   U1358 : HS65_LH_OAI21X3 port map( A => n1016, B => n1017, C => n280, Z => 
                           n1015);
   U1359 : HS65_LH_NAND4ABX3 port map( A => n1018, B => n1019, C => n1020, D =>
                           n1021, Z => n1017);
   U1360 : HS65_LH_OAI21X3 port map( A => n2760, B => n281, C => n1000, Z => 
                           regfile_o(63));
   U1361 : HS65_LH_OAI21X3 port map( A => n1001, B => n1002, C => n280, Z => 
                           n1000);
   U1362 : HS65_LH_NAND4ABX3 port map( A => n1003, B => n1004, C => n1005, D =>
                           n1006, Z => n1002);
   U1363 : HS65_LH_OAI21X3 port map( A => n285, B => n2698, C => n832, Z => 
                           regfile_o(0));
   U1364 : HS65_LH_OAI21X3 port map( A => n833, B => n834, C => n283, Z => n832
                           );
   U1365 : HS65_LH_NAND4ABX3 port map( A => n835, B => n836, C => n837, D => 
                           n838, Z => n834);
   U1366 : HS65_LH_OAI21X3 port map( A => n287, B => n2700, C => n667, Z => 
                           regfile_o(1));
   U1367 : HS65_LH_OAI21X3 port map( A => n668, B => n669, C => n284, Z => n667
                           );
   U1368 : HS65_LH_NAND4ABX3 port map( A => n670, B => n671, C => n672, D => 
                           n673, Z => n669);
   U1369 : HS65_LH_OAI21X3 port map( A => n286, B => n2702, C => n502, Z => 
                           regfile_o(2));
   U1370 : HS65_LH_OAI21X3 port map( A => n503, B => n504, C => n285, Z => n502
                           );
   U1371 : HS65_LH_NAND4ABX3 port map( A => n505, B => n506, C => n507, D => 
                           n508, Z => n504);
   U1372 : HS65_LH_OAI21X3 port map( A => n285, B => n2704, C => n457, Z => 
                           regfile_o(3));
   U1373 : HS65_LH_OAI21X3 port map( A => n458, B => n459, C => n284, Z => n457
                           );
   U1374 : HS65_LH_NAND4ABX3 port map( A => n460, B => n461, C => n462, D => 
                           n463, Z => n459);
   U1375 : HS65_LH_OAI21X3 port map( A => n286, B => n2706, C => n442, Z => 
                           regfile_o(4));
   U1376 : HS65_LH_OAI21X3 port map( A => n443, B => n444, C => n284, Z => n442
                           );
   U1377 : HS65_LH_NAND4ABX3 port map( A => n445, B => n446, C => n447, D => 
                           n448, Z => n444);
   U1378 : HS65_LH_OAI21X3 port map( A => n285, B => n2708, C => n427, Z => 
                           regfile_o(5));
   U1379 : HS65_LH_OAI21X3 port map( A => n428, B => n429, C => n284, Z => n427
                           );
   U1380 : HS65_LH_NAND4ABX3 port map( A => n430, B => n431, C => n432, D => 
                           n433, Z => n429);
   U1381 : HS65_LH_OAI21X3 port map( A => n285, B => n2710, C => n412, Z => 
                           regfile_o(6));
   U1382 : HS65_LH_OAI21X3 port map( A => n413, B => n414, C => n283, Z => n412
                           );
   U1383 : HS65_LH_NAND4ABX3 port map( A => n415, B => n416, C => n417, D => 
                           n418, Z => n414);
   U1384 : HS65_LH_OAI21X3 port map( A => n286, B => n2712, C => n397, Z => 
                           regfile_o(7));
   U1385 : HS65_LH_OAI21X3 port map( A => n398, B => n399, C => n283, Z => n397
                           );
   U1386 : HS65_LH_NAND4ABX3 port map( A => n400, B => n401, C => n402, D => 
                           n403, Z => n399);
   U1387 : HS65_LH_OAI21X3 port map( A => n285, B => n2714, C => n382, Z => 
                           regfile_o(8));
   U1388 : HS65_LH_OAI21X3 port map( A => n383, B => n384, C => n283, Z => n382
                           );
   U1389 : HS65_LH_NAND4ABX3 port map( A => n385, B => n386, C => n387, D => 
                           n388, Z => n384);
   U1390 : HS65_LH_OAI21X3 port map( A => n286, B => n2716, C => n335, Z => 
                           regfile_o(9));
   U1391 : HS65_LH_OAI21X3 port map( A => n336, B => n337, C => n283, Z => n335
                           );
   U1392 : HS65_LH_NAND4ABX3 port map( A => n338, B => n339, C => n340, D => 
                           n341, Z => n337);
   U1393 : HS65_LH_OAI21X3 port map( A => n287, B => n2720, C => n802, Z => 
                           regfile_o(11));
   U1394 : HS65_LH_OAI21X3 port map( A => n803, B => n804, C => n283, Z => n802
                           );
   U1395 : HS65_LH_NAND4ABX3 port map( A => n805, B => n806, C => n807, D => 
                           n808, Z => n804);
   U1396 : HS65_LH_OAI21X3 port map( A => n287, B => n2722, C => n787, Z => 
                           regfile_o(12));
   U1397 : HS65_LH_OAI21X3 port map( A => n788, B => n789, C => n283, Z => n787
                           );
   U1398 : HS65_LH_NAND4ABX3 port map( A => n790, B => n791, C => n792, D => 
                           n793, Z => n789);
   U1399 : HS65_LH_OAI21X3 port map( A => n287, B => n2724, C => n772, Z => 
                           regfile_o(13));
   U1400 : HS65_LH_OAI21X3 port map( A => n773, B => n774, C => n283, Z => n772
                           );
   U1401 : HS65_LH_NAND4ABX3 port map( A => n775, B => n776, C => n777, D => 
                           n778, Z => n774);
   U1402 : HS65_LH_OAI21X3 port map( A => n287, B => n2726, C => n757, Z => 
                           regfile_o(14));
   U1403 : HS65_LH_OAI21X3 port map( A => n758, B => n759, C => n283, Z => n757
                           );
   U1404 : HS65_LH_NAND4ABX3 port map( A => n760, B => n761, C => n762, D => 
                           n763, Z => n759);
   U1405 : HS65_LH_OAI21X3 port map( A => n287, B => n2728, C => n742, Z => 
                           regfile_o(15));
   U1406 : HS65_LH_OAI21X3 port map( A => n743, B => n744, C => n283, Z => n742
                           );
   U1407 : HS65_LH_NAND4ABX3 port map( A => n745, B => n746, C => n747, D => 
                           n748, Z => n744);
   U1408 : HS65_LH_OAI21X3 port map( A => n287, B => n2730, C => n727, Z => 
                           regfile_o(16));
   U1409 : HS65_LH_OAI21X3 port map( A => n728, B => n729, C => n283, Z => n727
                           );
   U1410 : HS65_LH_NAND4ABX3 port map( A => n730, B => n731, C => n732, D => 
                           n733, Z => n729);
   U1411 : HS65_LH_OAI21X3 port map( A => n287, B => n2732, C => n712, Z => 
                           regfile_o(17));
   U1412 : HS65_LH_OAI21X3 port map( A => n713, B => n714, C => n284, Z => n712
                           );
   U1413 : HS65_LH_NAND4ABX3 port map( A => n715, B => n716, C => n717, D => 
                           n718, Z => n714);
   U1414 : HS65_LH_OAI21X3 port map( A => n287, B => n2734, C => n697, Z => 
                           regfile_o(18));
   U1415 : HS65_LH_OAI21X3 port map( A => n698, B => n699, C => n284, Z => n697
                           );
   U1416 : HS65_LH_NAND4ABX3 port map( A => n700, B => n701, C => n702, D => 
                           n703, Z => n699);
   U1417 : HS65_LH_OAI21X3 port map( A => n287, B => n2736, C => n682, Z => 
                           regfile_o(19));
   U1418 : HS65_LH_OAI21X3 port map( A => n683, B => n684, C => n284, Z => n682
                           );
   U1419 : HS65_LH_NAND4ABX3 port map( A => n685, B => n686, C => n687, D => 
                           n688, Z => n684);
   U1420 : HS65_LH_OAI21X3 port map( A => n287, B => n2738, C => n652, Z => 
                           regfile_o(20));
   U1421 : HS65_LH_OAI21X3 port map( A => n653, B => n654, C => n284, Z => n652
                           );
   U1422 : HS65_LH_NAND4ABX3 port map( A => n655, B => n656, C => n657, D => 
                           n658, Z => n654);
   U1423 : HS65_LH_OAI21X3 port map( A => n287, B => n2740, C => n637, Z => 
                           regfile_o(21));
   U1424 : HS65_LH_OAI21X3 port map( A => n638, B => n639, C => n284, Z => n637
                           );
   U1425 : HS65_LH_NAND4ABX3 port map( A => n640, B => n641, C => n642, D => 
                           n643, Z => n639);
   U1426 : HS65_LH_OAI21X3 port map( A => n287, B => n2742, C => n622, Z => 
                           regfile_o(22));
   U1427 : HS65_LH_OAI21X3 port map( A => n623, B => n624, C => n284, Z => n622
                           );
   U1428 : HS65_LH_NAND4ABX3 port map( A => n625, B => n626, C => n627, D => 
                           n628, Z => n624);
   U1429 : HS65_LH_OAI21X3 port map( A => n286, B => n2744, C => n607, Z => 
                           regfile_o(23));
   U1430 : HS65_LH_OAI21X3 port map( A => n608, B => n609, C => n284, Z => n607
                           );
   U1431 : HS65_LH_NAND4ABX3 port map( A => n610, B => n611, C => n612, D => 
                           n613, Z => n609);
   U1432 : HS65_LH_OAI21X3 port map( A => n286, B => n2746, C => n592, Z => 
                           regfile_o(24));
   U1433 : HS65_LH_OAI21X3 port map( A => n593, B => n594, C => n285, Z => n592
                           );
   U1434 : HS65_LH_NAND4ABX3 port map( A => n595, B => n596, C => n597, D => 
                           n598, Z => n594);
   U1435 : HS65_LH_OAI21X3 port map( A => n286, B => n2748, C => n577, Z => 
                           regfile_o(25));
   U1436 : HS65_LH_OAI21X3 port map( A => n578, B => n579, C => n285, Z => n577
                           );
   U1437 : HS65_LH_NAND4ABX3 port map( A => n580, B => n581, C => n582, D => 
                           n583, Z => n579);
   U1438 : HS65_LH_OAI21X3 port map( A => n286, B => n2750, C => n562, Z => 
                           regfile_o(26));
   U1439 : HS65_LH_OAI21X3 port map( A => n563, B => n564, C => n284, Z => n562
                           );
   U1440 : HS65_LH_NAND4ABX3 port map( A => n565, B => n566, C => n567, D => 
                           n568, Z => n564);
   U1441 : HS65_LH_OAI21X3 port map( A => n286, B => n2752, C => n547, Z => 
                           regfile_o(27));
   U1442 : HS65_LH_OAI21X3 port map( A => n548, B => n549, C => n285, Z => n547
                           );
   U1443 : HS65_LH_NAND4ABX3 port map( A => n550, B => n551, C => n552, D => 
                           n553, Z => n549);
   U1444 : HS65_LH_OAI21X3 port map( A => n286, B => n2754, C => n532, Z => 
                           regfile_o(28));
   U1445 : HS65_LH_OAI21X3 port map( A => n533, B => n534, C => n285, Z => n532
                           );
   U1446 : HS65_LH_NAND4ABX3 port map( A => n535, B => n536, C => n537, D => 
                           n538, Z => n534);
   U1447 : HS65_LH_OAI21X3 port map( A => n286, B => n2756, C => n517, Z => 
                           regfile_o(29));
   U1448 : HS65_LH_OAI21X3 port map( A => n518, B => n519, C => n285, Z => n517
                           );
   U1449 : HS65_LH_NAND4ABX3 port map( A => n520, B => n521, C => n522, D => 
                           n523, Z => n519);
   U1450 : HS65_LH_OAI21X3 port map( A => n286, B => n2758, C => n487, Z => 
                           regfile_o(30));
   U1451 : HS65_LH_OAI21X3 port map( A => n488, B => n489, C => n285, Z => n487
                           );
   U1452 : HS65_LH_NAND4ABX3 port map( A => n490, B => n491, C => n492, D => 
                           n493, Z => n489);
   U1453 : HS65_LH_OAI21X3 port map( A => n286, B => n2760, C => n472, Z => 
                           regfile_o(31));
   U1454 : HS65_LH_OAI21X3 port map( A => n473, B => n474, C => n285, Z => n472
                           );
   U1455 : HS65_LH_NAND4ABX3 port map( A => n475, B => n476, C => n477, D => 
                           n478, Z => n474);
   U1456 : HS65_LH_OAI21X3 port map( A => n287, B => n2718, C => n817, Z => 
                           regfile_o(10));
   U1457 : HS65_LH_OAI21X3 port map( A => n818, B => n819, C => n283, Z => n817
                           );
   U1458 : HS65_LH_AOI212X4 port map( A => registers_11_3_port, B => n2684, C 
                           => registers_10_3_port, D => n2680, E => n465, Z => 
                           n462);
   U1459 : HS65_LH_OAI22X6 port map( A => n2678, B => n253, C => n2674, D => 
                           n221, Z => n465);
   U1460 : HS65_LH_AOI212X4 port map( A => registers_11_4_port, B => n2684, C 
                           => registers_10_4_port, D => n2681, E => n450, Z => 
                           n447);
   U1461 : HS65_LH_OAI22X6 port map( A => n2678, B => n252, C => n2675, D => 
                           n220, Z => n450);
   U1462 : HS65_LH_AOI212X4 port map( A => registers_11_5_port, B => n2684, C 
                           => registers_10_5_port, D => n2681, E => n435, Z => 
                           n432);
   U1463 : HS65_LH_OAI22X6 port map( A => n2678, B => n251, C => n2675, D => 
                           n219, Z => n435);
   U1464 : HS65_LH_AOI212X4 port map( A => registers_11_6_port, B => n2684, C 
                           => registers_10_6_port, D => n2681, E => n420, Z => 
                           n417);
   U1465 : HS65_LH_OAI22X6 port map( A => n2678, B => n250, C => n2675, D => 
                           n218, Z => n420);
   U1466 : HS65_LH_AOI212X4 port map( A => registers_11_7_port, B => n2684, C 
                           => registers_10_7_port, D => n2681, E => n405, Z => 
                           n402);
   U1467 : HS65_LH_OAI22X6 port map( A => n2678, B => n249, C => n2675, D => 
                           n217, Z => n405);
   U1468 : HS65_LH_AOI212X4 port map( A => registers_11_8_port, B => n2684, C 
                           => registers_10_8_port, D => n2681, E => n390, Z => 
                           n387);
   U1469 : HS65_LH_OAI22X6 port map( A => n2678, B => n248, C => n2675, D => 
                           n216, Z => n390);
   U1470 : HS65_LH_AOI212X4 port map( A => registers_11_9_port, B => n2684, C 
                           => registers_10_9_port, D => n2681, E => n349, Z => 
                           n340);
   U1471 : HS65_LH_OAI22X6 port map( A => n2678, B => n247, C => n2675, D => 
                           n215, Z => n349);
   U1472 : HS65_LH_AOI212X4 port map( A => registers_11_31_port, B => n2684, C 
                           => registers_10_31_port, D => n2680, E => n480, Z =>
                           n477);
   U1473 : HS65_LH_OAI22X6 port map( A => n2678, B => n225, C => n2674, D => 
                           n193, Z => n480);
   U1474 : HS65_LH_AOI212X4 port map( A => registers_13_0_port, B => n2694, C 
                           => registers_12_0_port, D => n2691, E => n839, Z => 
                           n838);
   U1475 : HS65_LH_OAI22X6 port map( A => n2688, B => n192, C => n2685, D => 
                           n160, Z => n839);
   U1476 : HS65_LH_AOI212X4 port map( A => registers_13_1_port, B => n2694, C 
                           => registers_12_1_port, D => n2691, E => n674, Z => 
                           n673);
   U1477 : HS65_LH_OAI22X6 port map( A => n2688, B => n191, C => n2685, D => 
                           n159, Z => n674);
   U1478 : HS65_LH_AOI212X4 port map( A => registers_13_2_port, B => n2695, C 
                           => registers_12_2_port, D => n2692, E => n509, Z => 
                           n508);
   U1479 : HS65_LH_OAI22X6 port map( A => n2689, B => n190, C => n2686, D => 
                           n158, Z => n509);
   U1480 : HS65_LH_AOI212X4 port map( A => registers_13_3_port, B => n2696, C 
                           => registers_12_3_port, D => n2692, E => n464, Z => 
                           n463);
   U1481 : HS65_LH_OAI22X6 port map( A => n2690, B => n189, C => n2686, D => 
                           n157, Z => n464);
   U1482 : HS65_LH_AOI212X4 port map( A => registers_13_4_port, B => n2696, C 
                           => registers_12_4_port, D => n2693, E => n449, Z => 
                           n448);
   U1483 : HS65_LH_OAI22X6 port map( A => n2690, B => n188, C => n2687, D => 
                           n156, Z => n449);
   U1484 : HS65_LH_AOI212X4 port map( A => registers_13_5_port, B => n2696, C 
                           => registers_12_5_port, D => n2693, E => n434, Z => 
                           n433);
   U1485 : HS65_LH_OAI22X6 port map( A => n2690, B => n187, C => n2687, D => 
                           n155, Z => n434);
   U1486 : HS65_LH_AOI212X4 port map( A => registers_13_6_port, B => n2696, C 
                           => registers_12_6_port, D => n2693, E => n419, Z => 
                           n418);
   U1487 : HS65_LH_OAI22X6 port map( A => n2690, B => n186, C => n2687, D => 
                           n154, Z => n419);
   U1488 : HS65_LH_AOI212X4 port map( A => registers_13_7_port, B => n2696, C 
                           => registers_12_7_port, D => n2693, E => n404, Z => 
                           n403);
   U1489 : HS65_LH_OAI22X6 port map( A => n2690, B => n185, C => n2687, D => 
                           n153, Z => n404);
   U1490 : HS65_LH_AOI212X4 port map( A => registers_13_8_port, B => n2696, C 
                           => registers_12_8_port, D => n2693, E => n389, Z => 
                           n388);
   U1491 : HS65_LH_OAI22X6 port map( A => n2690, B => n184, C => n2687, D => 
                           n152, Z => n389);
   U1492 : HS65_LH_AOI212X4 port map( A => registers_13_9_port, B => n2696, C 
                           => registers_12_9_port, D => n2693, E => n344, Z => 
                           n341);
   U1493 : HS65_LH_OAI22X6 port map( A => n2690, B => n183, C => n2687, D => 
                           n151, Z => n344);
   U1494 : HS65_LH_AOI212X4 port map( A => registers_13_11_port, B => n2694, C 
                           => registers_12_11_port, D => n2691, E => n809, Z =>
                           n808);
   U1495 : HS65_LH_OAI22X6 port map( A => n2688, B => n181, C => n2685, D => 
                           n149, Z => n809);
   U1496 : HS65_LH_AOI212X4 port map( A => registers_13_12_port, B => n2694, C 
                           => registers_12_12_port, D => n2691, E => n794, Z =>
                           n793);
   U1497 : HS65_LH_OAI22X6 port map( A => n2688, B => n180, C => n2685, D => 
                           n148, Z => n794);
   U1498 : HS65_LH_AOI212X4 port map( A => registers_13_13_port, B => n2694, C 
                           => registers_12_13_port, D => n2691, E => n779, Z =>
                           n778);
   U1499 : HS65_LH_OAI22X6 port map( A => n2688, B => n179, C => n2685, D => 
                           n147, Z => n779);
   U1500 : HS65_LH_AOI212X4 port map( A => registers_13_14_port, B => n2694, C 
                           => registers_12_14_port, D => n2691, E => n764, Z =>
                           n763);
   U1501 : HS65_LH_OAI22X6 port map( A => n2688, B => n178, C => n2685, D => 
                           n146, Z => n764);
   U1502 : HS65_LH_AOI212X4 port map( A => registers_13_15_port, B => n2694, C 
                           => registers_12_15_port, D => n2691, E => n749, Z =>
                           n748);
   U1503 : HS65_LH_OAI22X6 port map( A => n2688, B => n177, C => n2685, D => 
                           n145, Z => n749);
   U1504 : HS65_LH_AOI212X4 port map( A => registers_13_16_port, B => n2694, C 
                           => registers_12_16_port, D => n2691, E => n734, Z =>
                           n733);
   U1505 : HS65_LH_OAI22X6 port map( A => n2688, B => n176, C => n2685, D => 
                           n144, Z => n734);
   U1506 : HS65_LH_AOI212X4 port map( A => registers_13_17_port, B => n2694, C 
                           => registers_12_17_port, D => n2691, E => n719, Z =>
                           n718);
   U1507 : HS65_LH_OAI22X6 port map( A => n2688, B => n175, C => n2685, D => 
                           n143, Z => n719);
   U1508 : HS65_LH_AOI212X4 port map( A => registers_13_18_port, B => n2694, C 
                           => registers_12_18_port, D => n2691, E => n704, Z =>
                           n703);
   U1509 : HS65_LH_OAI22X6 port map( A => n2688, B => n174, C => n2685, D => 
                           n142, Z => n704);
   U1510 : HS65_LH_AOI212X4 port map( A => registers_13_19_port, B => n2694, C 
                           => registers_12_19_port, D => n2691, E => n689, Z =>
                           n688);
   U1511 : HS65_LH_OAI22X6 port map( A => n2688, B => n173, C => n2685, D => 
                           n141, Z => n689);
   U1512 : HS65_LH_AOI212X4 port map( A => registers_13_20_port, B => n2695, C 
                           => registers_12_20_port, D => n2691, E => n659, Z =>
                           n658);
   U1513 : HS65_LH_OAI22X6 port map( A => n2689, B => n172, C => n2685, D => 
                           n140, Z => n659);
   U1514 : HS65_LH_AOI212X4 port map( A => registers_13_21_port, B => n2695, C 
                           => registers_12_21_port, D => n2692, E => n644, Z =>
                           n643);
   U1515 : HS65_LH_OAI22X6 port map( A => n2689, B => n171, C => n2686, D => 
                           n139, Z => n644);
   U1516 : HS65_LH_AOI212X4 port map( A => registers_13_22_port, B => n2695, C 
                           => registers_12_22_port, D => n2692, E => n629, Z =>
                           n628);
   U1517 : HS65_LH_OAI22X6 port map( A => n2689, B => n170, C => n2686, D => 
                           n138, Z => n629);
   U1518 : HS65_LH_AOI212X4 port map( A => registers_13_23_port, B => n2695, C 
                           => registers_12_23_port, D => n2692, E => n614, Z =>
                           n613);
   U1519 : HS65_LH_OAI22X6 port map( A => n2689, B => n169, C => n2686, D => 
                           n137, Z => n614);
   U1520 : HS65_LH_AOI212X4 port map( A => registers_13_24_port, B => n2695, C 
                           => registers_12_24_port, D => n2692, E => n599, Z =>
                           n598);
   U1521 : HS65_LH_OAI22X6 port map( A => n2689, B => n168, C => n2686, D => 
                           n136, Z => n599);
   U1522 : HS65_LH_AOI212X4 port map( A => registers_13_25_port, B => n2695, C 
                           => registers_12_25_port, D => n2692, E => n584, Z =>
                           n583);
   U1523 : HS65_LH_OAI22X6 port map( A => n2689, B => n167, C => n2686, D => 
                           n135, Z => n584);
   U1524 : HS65_LH_AOI212X4 port map( A => registers_13_26_port, B => n2695, C 
                           => registers_12_26_port, D => n2692, E => n569, Z =>
                           n568);
   U1525 : HS65_LH_OAI22X6 port map( A => n2689, B => n166, C => n2686, D => 
                           n134, Z => n569);
   U1526 : HS65_LH_AOI212X4 port map( A => registers_13_27_port, B => n2695, C 
                           => registers_12_27_port, D => n2692, E => n554, Z =>
                           n553);
   U1527 : HS65_LH_OAI22X6 port map( A => n2689, B => n165, C => n2686, D => 
                           n133, Z => n554);
   U1528 : HS65_LH_AOI212X4 port map( A => registers_13_28_port, B => n2695, C 
                           => registers_12_28_port, D => n2692, E => n539, Z =>
                           n538);
   U1529 : HS65_LH_OAI22X6 port map( A => n2689, B => n164, C => n2686, D => 
                           n132, Z => n539);
   U1530 : HS65_LH_AOI212X4 port map( A => registers_13_29_port, B => n2695, C 
                           => registers_12_29_port, D => n2692, E => n524, Z =>
                           n523);
   U1531 : HS65_LH_OAI22X6 port map( A => n2689, B => n163, C => n2686, D => 
                           n131, Z => n524);
   U1532 : HS65_LH_AOI212X4 port map( A => registers_13_30_port, B => n2695, C 
                           => registers_12_30_port, D => n2692, E => n494, Z =>
                           n493);
   U1533 : HS65_LH_OAI22X6 port map( A => n2689, B => n162, C => n2686, D => 
                           n130, Z => n494);
   U1534 : HS65_LH_AOI212X4 port map( A => registers_13_31_port, B => n2696, C 
                           => registers_12_31_port, D => n2692, E => n479, Z =>
                           n478);
   U1535 : HS65_LH_OAI22X6 port map( A => n2690, B => n161, C => n2686, D => 
                           n129, Z => n479);
   U1536 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_4_port, C 
                           => n2600, D => registers_12_4_port, E => n977, Z => 
                           n976);
   U1537 : HS65_LH_OAI22X6 port map( A => n188, B => n2597, C => n156, D => 
                           n2594, Z => n977);
   U1538 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_5_port, C 
                           => n2600, D => registers_12_5_port, E => n962, Z => 
                           n961);
   U1539 : HS65_LH_OAI22X6 port map( A => n187, B => n2597, C => n155, D => 
                           n2594, Z => n962);
   U1540 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_6_port, C 
                           => n2600, D => registers_12_6_port, E => n947, Z => 
                           n946);
   U1541 : HS65_LH_OAI22X6 port map( A => n186, B => n2597, C => n154, D => 
                           n2594, Z => n947);
   U1542 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_7_port, C 
                           => n2600, D => registers_12_7_port, E => n932, Z => 
                           n931);
   U1543 : HS65_LH_OAI22X6 port map( A => n185, B => n2597, C => n153, D => 
                           n2594, Z => n932);
   U1544 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_8_port, C 
                           => n2600, D => registers_12_8_port, E => n917, Z => 
                           n916);
   U1545 : HS65_LH_OAI22X6 port map( A => n184, B => n2597, C => n152, D => 
                           n2594, Z => n917);
   U1546 : HS65_LH_AOI212X4 port map( A => n2603, B => registers_13_9_port, C 
                           => n2600, D => registers_12_9_port, E => n872, Z => 
                           n869);
   U1547 : HS65_LH_OAI22X6 port map( A => n183, B => n2597, C => n151, D => 
                           n2594, Z => n872);
   U1548 : HS65_LH_OAI22X6 port map( A => n2643, B => n64, C => n2640, D => n32
                           , Z => n855);
   U1549 : HS65_LH_OAI22X6 port map( A => n2643, B => n63, C => n2640, D => n31
                           , Z => n680);
   U1550 : HS65_LH_OAI22X6 port map( A => n2644, B => n62, C => n2641, D => n30
                           , Z => n515);
   U1551 : HS65_LH_OAI22X6 port map( A => n2633, B => n125, C => n2629, D => 
                           n93, Z => n471);
   U1552 : HS65_LH_OAI22X6 port map( A => n2645, B => n61, C => n2641, D => n29
                           , Z => n470);
   U1553 : HS65_LH_OAI22X6 port map( A => n2633, B => n124, C => n2630, D => 
                           n92, Z => n456);
   U1554 : HS65_LH_OAI22X6 port map( A => n2645, B => n60, C => n2642, D => n28
                           , Z => n455);
   U1555 : HS65_LH_OAI22X6 port map( A => n2633, B => n123, C => n2630, D => 
                           n91, Z => n441);
   U1556 : HS65_LH_OAI22X6 port map( A => n2645, B => n59, C => n2642, D => n27
                           , Z => n440);
   U1557 : HS65_LH_OAI22X6 port map( A => n2633, B => n122, C => n2630, D => 
                           n90, Z => n426);
   U1558 : HS65_LH_OAI22X6 port map( A => n2645, B => n58, C => n2642, D => n26
                           , Z => n425);
   U1559 : HS65_LH_OAI22X6 port map( A => n2633, B => n121, C => n2630, D => 
                           n89, Z => n411);
   U1560 : HS65_LH_OAI22X6 port map( A => n2645, B => n57, C => n2642, D => n25
                           , Z => n410);
   U1561 : HS65_LH_OAI22X6 port map( A => n2633, B => n120, C => n2630, D => 
                           n88, Z => n396);
   U1562 : HS65_LH_OAI22X6 port map( A => n2645, B => n56, C => n2642, D => n24
                           , Z => n395);
   U1563 : HS65_LH_OAI22X6 port map( A => n2633, B => n119, C => n2630, D => 
                           n87, Z => n371);
   U1564 : HS65_LH_OAI22X6 port map( A => n2645, B => n55, C => n2642, D => n23
                           , Z => n366);
   U1565 : HS65_LH_OAI22X6 port map( A => n2643, B => n54, C => n2640, D => n22
                           , Z => n830);
   U1566 : HS65_LH_OAI22X6 port map( A => n2676, B => n246, C => n2673, D => 
                           n214, Z => n825);
   U1567 : HS65_LH_OAI22X6 port map( A => n2688, B => n182, C => n2685, D => 
                           n150, Z => n824);
   U1568 : HS65_LH_OAI22X6 port map( A => n2643, B => n53, C => n2640, D => n21
                           , Z => n815);
   U1569 : HS65_LH_OAI22X6 port map( A => n2643, B => n52, C => n2640, D => n20
                           , Z => n800);
   U1570 : HS65_LH_OAI22X6 port map( A => n2643, B => n51, C => n2640, D => n19
                           , Z => n785);
   U1571 : HS65_LH_OAI22X6 port map( A => n2643, B => n50, C => n2640, D => n18
                           , Z => n770);
   U1572 : HS65_LH_OAI22X6 port map( A => n2643, B => n49, C => n2640, D => n17
                           , Z => n755);
   U1573 : HS65_LH_OAI22X6 port map( A => n2643, B => n48, C => n2640, D => n16
                           , Z => n740);
   U1574 : HS65_LH_OAI22X6 port map( A => n2643, B => n47, C => n2640, D => n15
                           , Z => n725);
   U1575 : HS65_LH_OAI22X6 port map( A => n2643, B => n46, C => n2640, D => n14
                           , Z => n710);
   U1576 : HS65_LH_OAI22X6 port map( A => n2643, B => n45, C => n2640, D => n13
                           , Z => n695);
   U1577 : HS65_LH_OAI22X6 port map( A => n2644, B => n44, C => n2640, D => n12
                           , Z => n665);
   U1578 : HS65_LH_OAI22X6 port map( A => n2644, B => n43, C => n2641, D => n11
                           , Z => n650);
   U1579 : HS65_LH_OAI22X6 port map( A => n2644, B => n42, C => n2641, D => n10
                           , Z => n635);
   U1580 : HS65_LH_OAI22X6 port map( A => n2644, B => n41, C => n2641, D => n9,
                           Z => n620);
   U1581 : HS65_LH_OAI22X6 port map( A => n2644, B => n40, C => n2641, D => n8,
                           Z => n605);
   U1582 : HS65_LH_OAI22X6 port map( A => n2644, B => n39, C => n2641, D => n7,
                           Z => n590);
   U1583 : HS65_LH_OAI22X6 port map( A => n2644, B => n38, C => n2641, D => n6,
                           Z => n575);
   U1584 : HS65_LH_OAI22X6 port map( A => n2644, B => n37, C => n2641, D => n5,
                           Z => n560);
   U1585 : HS65_LH_OAI22X6 port map( A => n2644, B => n36, C => n2641, D => n4,
                           Z => n545);
   U1586 : HS65_LH_OAI22X6 port map( A => n2644, B => n35, C => n2641, D => n3,
                           Z => n530);
   U1587 : HS65_LH_OAI22X6 port map( A => n2644, B => n34, C => n2641, D => n2,
                           Z => n500);
   U1588 : HS65_LH_OAI22X6 port map( A => n2633, B => n97, C => n2629, D => n65
                           , Z => n486);
   U1589 : HS65_LH_OAI22X6 port map( A => n2645, B => n33, C => n2641, D => n1,
                           Z => n485);
   U1590 : HS65_LH_OAI22X6 port map( A => n128, B => n2538, C => n96, D => 
                           n2535, Z => n1386);
   U1591 : HS65_LH_OAI22X6 port map( A => n64, B => n2550, C => n32, D => n2547
                           , Z => n1383);
   U1592 : HS65_LH_OAI22X6 port map( A => n127, B => n2538, C => n95, D => 
                           n2535, Z => n1209);
   U1593 : HS65_LH_OAI22X6 port map( A => n63, B => n2550, C => n31, D => n2547
                           , Z => n1208);
   U1594 : HS65_LH_OAI22X6 port map( A => n126, B => n2539, C => n94, D => 
                           n2536, Z => n1044);
   U1595 : HS65_LH_OAI22X6 port map( A => n62, B => n2551, C => n30, D => n2548
                           , Z => n1043);
   U1596 : HS65_LH_OAI22X6 port map( A => n118, B => n2538, C => n86, D => 
                           n2535, Z => n1359);
   U1597 : HS65_LH_OAI22X6 port map( A => n54, B => n2550, C => n22, D => n2547
                           , Z => n1358);
   U1598 : HS65_LH_OAI22X6 port map( A => n117, B => n2538, C => n85, D => 
                           n2535, Z => n1344);
   U1599 : HS65_LH_OAI22X6 port map( A => n53, B => n2550, C => n21, D => n2547
                           , Z => n1343);
   U1600 : HS65_LH_OAI22X6 port map( A => n116, B => n2538, C => n84, D => 
                           n2535, Z => n1329);
   U1601 : HS65_LH_OAI22X6 port map( A => n52, B => n2550, C => n20, D => n2547
                           , Z => n1328);
   U1602 : HS65_LH_OAI22X6 port map( A => n115, B => n2538, C => n83, D => 
                           n2535, Z => n1314);
   U1603 : HS65_LH_OAI22X6 port map( A => n51, B => n2550, C => n19, D => n2547
                           , Z => n1313);
   U1604 : HS65_LH_OAI22X6 port map( A => n114, B => n2538, C => n82, D => 
                           n2535, Z => n1299);
   U1605 : HS65_LH_OAI22X6 port map( A => n50, B => n2550, C => n18, D => n2547
                           , Z => n1298);
   U1606 : HS65_LH_OAI22X6 port map( A => n113, B => n2538, C => n81, D => 
                           n2535, Z => n1284);
   U1607 : HS65_LH_OAI22X6 port map( A => n49, B => n2550, C => n17, D => n2547
                           , Z => n1283);
   U1608 : HS65_LH_OAI22X6 port map( A => n112, B => n2538, C => n80, D => 
                           n2535, Z => n1269);
   U1609 : HS65_LH_OAI22X6 port map( A => n48, B => n2550, C => n16, D => n2547
                           , Z => n1268);
   U1610 : HS65_LH_OAI22X6 port map( A => n111, B => n2538, C => n79, D => 
                           n2535, Z => n1254);
   U1611 : HS65_LH_OAI22X6 port map( A => n47, B => n2550, C => n15, D => n2547
                           , Z => n1253);
   U1612 : HS65_LH_OAI22X6 port map( A => n110, B => n2538, C => n78, D => 
                           n2535, Z => n1239);
   U1613 : HS65_LH_OAI22X6 port map( A => n46, B => n2550, C => n14, D => n2547
                           , Z => n1238);
   U1614 : HS65_LH_OAI22X6 port map( A => n109, B => n2538, C => n77, D => 
                           n2535, Z => n1224);
   U1615 : HS65_LH_OAI22X6 port map( A => n45, B => n2550, C => n13, D => n2547
                           , Z => n1223);
   U1616 : HS65_LH_OAI22X6 port map( A => n108, B => n2539, C => n76, D => 
                           n2535, Z => n1194);
   U1617 : HS65_LH_OAI22X6 port map( A => n44, B => n2551, C => n12, D => n2547
                           , Z => n1193);
   U1618 : HS65_LH_OAI22X6 port map( A => n107, B => n2539, C => n75, D => 
                           n2536, Z => n1179);
   U1619 : HS65_LH_OAI22X6 port map( A => n43, B => n2551, C => n11, D => n2548
                           , Z => n1178);
   U1620 : HS65_LH_OAI22X6 port map( A => n106, B => n2539, C => n74, D => 
                           n2536, Z => n1164);
   U1621 : HS65_LH_OAI22X6 port map( A => n42, B => n2551, C => n10, D => n2548
                           , Z => n1163);
   U1622 : HS65_LH_OAI22X6 port map( A => n105, B => n2539, C => n73, D => 
                           n2536, Z => n1149);
   U1623 : HS65_LH_OAI22X6 port map( A => n41, B => n2551, C => n9, D => n2548,
                           Z => n1148);
   U1624 : HS65_LH_OAI22X6 port map( A => n104, B => n2539, C => n72, D => 
                           n2536, Z => n1134);
   U1625 : HS65_LH_OAI22X6 port map( A => n40, B => n2551, C => n8, D => n2548,
                           Z => n1133);
   U1626 : HS65_LH_OAI22X6 port map( A => n103, B => n2539, C => n71, D => 
                           n2536, Z => n1119);
   U1627 : HS65_LH_OAI22X6 port map( A => n39, B => n2551, C => n7, D => n2548,
                           Z => n1118);
   U1628 : HS65_LH_OAI22X6 port map( A => n102, B => n2539, C => n70, D => 
                           n2536, Z => n1104);
   U1629 : HS65_LH_OAI22X6 port map( A => n38, B => n2551, C => n6, D => n2548,
                           Z => n1103);
   U1630 : HS65_LH_OAI22X6 port map( A => n101, B => n2539, C => n69, D => 
                           n2536, Z => n1089);
   U1631 : HS65_LH_OAI22X6 port map( A => n37, B => n2551, C => n5, D => n2548,
                           Z => n1088);
   U1632 : HS65_LH_OAI22X6 port map( A => n100, B => n2539, C => n68, D => 
                           n2536, Z => n1074);
   U1633 : HS65_LH_OAI22X6 port map( A => n36, B => n2551, C => n4, D => n2548,
                           Z => n1073);
   U1634 : HS65_LH_OAI22X6 port map( A => n99, B => n2539, C => n67, D => n2536
                           , Z => n1059);
   U1635 : HS65_LH_OAI22X6 port map( A => n35, B => n2551, C => n3, D => n2548,
                           Z => n1058);
   U1636 : HS65_LH_OAI22X6 port map( A => n98, B => n2539, C => n66, D => n2536
                           , Z => n1029);
   U1637 : HS65_LH_OAI22X6 port map( A => n34, B => n2551, C => n2, D => n2548,
                           Z => n1028);
   U1638 : HS65_LH_OAI22X6 port map( A => n125, B => n2540, C => n93, D => 
                           n2536, Z => n999);
   U1639 : HS65_LH_OAI22X6 port map( A => n61, B => n2552, C => n29, D => n2548
                           , Z => n998);
   U1640 : HS65_LH_OAI22X6 port map( A => n124, B => n2540, C => n92, D => 
                           n2537, Z => n984);
   U1641 : HS65_LH_OAI22X6 port map( A => n60, B => n2552, C => n28, D => n2549
                           , Z => n983);
   U1642 : HS65_LH_OAI22X6 port map( A => n123, B => n2540, C => n91, D => 
                           n2537, Z => n969);
   U1643 : HS65_LH_OAI22X6 port map( A => n59, B => n2552, C => n27, D => n2549
                           , Z => n968);
   U1644 : HS65_LH_OAI22X6 port map( A => n122, B => n2540, C => n90, D => 
                           n2537, Z => n954);
   U1645 : HS65_LH_OAI22X6 port map( A => n58, B => n2552, C => n26, D => n2549
                           , Z => n953);
   U1646 : HS65_LH_OAI22X6 port map( A => n121, B => n2540, C => n89, D => 
                           n2537, Z => n939);
   U1647 : HS65_LH_OAI22X6 port map( A => n57, B => n2552, C => n25, D => n2549
                           , Z => n938);
   U1648 : HS65_LH_OAI22X6 port map( A => n120, B => n2540, C => n88, D => 
                           n2537, Z => n924);
   U1649 : HS65_LH_OAI22X6 port map( A => n56, B => n2552, C => n24, D => n2549
                           , Z => n923);
   U1650 : HS65_LH_OAI22X6 port map( A => n119, B => n2540, C => n87, D => 
                           n2537, Z => n899);
   U1651 : HS65_LH_OAI22X6 port map( A => n55, B => n2552, C => n23, D => n2549
                           , Z => n894);
   U1652 : HS65_LH_OAI22X6 port map( A => n97, B => n2540, C => n65, D => n2536
                           , Z => n1014);
   U1653 : HS65_LH_OAI22X6 port map( A => n33, B => n2552, C => n1, D => n2548,
                           Z => n1013);
   U1654 : HS65_LH_OAI22X6 port map( A => n2760, B => n2473, C => n2471, D => 
                           n225, Z => n1689);
   U1655 : HS65_LH_OAI22X6 port map( A => n2760, B => n2468, C => n2466, D => 
                           n193, Z => n1721);
   U1656 : HS65_LH_OAI22X6 port map( A => n2760, B => n2443, C => n2441, D => 
                           n161, Z => n1881);
   U1657 : HS65_LH_OAI22X6 port map( A => n2760, B => n2438, C => n2436, D => 
                           n129, Z => n1913);
   U1658 : HS65_LH_OAI22X6 port map( A => n2760, B => n305, C => n303, D => n33
                           , Z => n2329);
   U1659 : HS65_LH_OAI22X6 port map( A => n2760, B => n300, C => n298, D => n1,
                           Z => n2361);
   U1660 : HS65_LH_OAI22X6 port map( A => n2760, B => n315, C => n313, D => n97
                           , Z => n2265);
   U1661 : HS65_LH_OAI22X6 port map( A => n2760, B => n310, C => n308, D => n65
                           , Z => n2297);
   U1662 : HS65_LH_OAI22X6 port map( A => n2724, B => n2474, C => n2472, D => 
                           n243, Z => n1671);
   U1663 : HS65_LH_OAI22X6 port map( A => n2726, B => n2474, C => n2472, D => 
                           n242, Z => n1672);
   U1664 : HS65_LH_OAI22X6 port map( A => n2728, B => n2474, C => n2472, D => 
                           n241, Z => n1673);
   U1665 : HS65_LH_OAI22X6 port map( A => n2730, B => n2474, C => n2472, D => 
                           n240, Z => n1674);
   U1666 : HS65_LH_OAI22X6 port map( A => n2732, B => n2474, C => n2472, D => 
                           n239, Z => n1675);
   U1667 : HS65_LH_OAI22X6 port map( A => n2734, B => n2474, C => n2472, D => 
                           n238, Z => n1676);
   U1668 : HS65_LH_OAI22X6 port map( A => n2736, B => n2474, C => n2471, D => 
                           n237, Z => n1677);
   U1669 : HS65_LH_OAI22X6 port map( A => n2738, B => n2474, C => n2471, D => 
                           n236, Z => n1678);
   U1670 : HS65_LH_OAI22X6 port map( A => n2740, B => n2474, C => n2471, D => 
                           n235, Z => n1679);
   U1671 : HS65_LH_OAI22X6 port map( A => n2742, B => n2474, C => n2471, D => 
                           n234, Z => n1680);
   U1672 : HS65_LH_OAI22X6 port map( A => n2744, B => n2474, C => n2471, D => 
                           n233, Z => n1681);
   U1673 : HS65_LH_OAI22X6 port map( A => n2746, B => n2474, C => n2471, D => 
                           n232, Z => n1682);
   U1674 : HS65_LH_OAI22X6 port map( A => n2748, B => n2474, C => n2471, D => 
                           n231, Z => n1683);
   U1675 : HS65_LH_OAI22X6 port map( A => n2750, B => n2474, C => n2471, D => 
                           n230, Z => n1684);
   U1676 : HS65_LH_OAI22X6 port map( A => n2752, B => n2474, C => n2471, D => 
                           n229, Z => n1685);
   U1677 : HS65_LH_OAI22X6 port map( A => n2754, B => n2474, C => n2471, D => 
                           n228, Z => n1686);
   U1678 : HS65_LH_OAI22X6 port map( A => n2756, B => n2474, C => n2471, D => 
                           n227, Z => n1687);
   U1679 : HS65_LH_OAI22X6 port map( A => n2758, B => n2474, C => n2471, D => 
                           n226, Z => n1688);
   U1680 : HS65_LH_OAI22X6 port map( A => n2724, B => n2469, C => n2467, D => 
                           n211, Z => n1703);
   U1681 : HS65_LH_OAI22X6 port map( A => n2726, B => n2469, C => n2467, D => 
                           n210, Z => n1704);
   U1682 : HS65_LH_OAI22X6 port map( A => n2728, B => n2469, C => n2467, D => 
                           n209, Z => n1705);
   U1683 : HS65_LH_OAI22X6 port map( A => n2730, B => n2469, C => n2467, D => 
                           n208, Z => n1706);
   U1684 : HS65_LH_OAI22X6 port map( A => n2732, B => n2469, C => n2467, D => 
                           n207, Z => n1707);
   U1685 : HS65_LH_OAI22X6 port map( A => n2734, B => n2469, C => n2467, D => 
                           n206, Z => n1708);
   U1686 : HS65_LH_OAI22X6 port map( A => n2736, B => n2469, C => n2466, D => 
                           n205, Z => n1709);
   U1687 : HS65_LH_OAI22X6 port map( A => n2738, B => n2469, C => n2466, D => 
                           n204, Z => n1710);
   U1688 : HS65_LH_OAI22X6 port map( A => n2740, B => n2469, C => n2466, D => 
                           n203, Z => n1711);
   U1689 : HS65_LH_OAI22X6 port map( A => n2742, B => n2469, C => n2466, D => 
                           n202, Z => n1712);
   U1690 : HS65_LH_OAI22X6 port map( A => n2744, B => n2469, C => n2466, D => 
                           n201, Z => n1713);
   U1691 : HS65_LH_OAI22X6 port map( A => n2746, B => n2469, C => n2466, D => 
                           n200, Z => n1714);
   U1692 : HS65_LH_OAI22X6 port map( A => n2748, B => n2469, C => n2466, D => 
                           n199, Z => n1715);
   U1693 : HS65_LH_OAI22X6 port map( A => n2750, B => n2469, C => n2466, D => 
                           n198, Z => n1716);
   U1694 : HS65_LH_OAI22X6 port map( A => n2752, B => n2469, C => n2466, D => 
                           n197, Z => n1717);
   U1695 : HS65_LH_OAI22X6 port map( A => n2754, B => n2469, C => n2466, D => 
                           n196, Z => n1718);
   U1696 : HS65_LH_OAI22X6 port map( A => n2756, B => n2469, C => n2466, D => 
                           n195, Z => n1719);
   U1697 : HS65_LH_OAI22X6 port map( A => n2758, B => n2469, C => n2466, D => 
                           n194, Z => n1720);
   U1698 : HS65_LH_OAI22X6 port map( A => n2724, B => n2444, C => n2442, D => 
                           n179, Z => n1863);
   U1699 : HS65_LH_OAI22X6 port map( A => n2726, B => n2444, C => n2442, D => 
                           n178, Z => n1864);
   U1700 : HS65_LH_OAI22X6 port map( A => n2728, B => n2444, C => n2442, D => 
                           n177, Z => n1865);
   U1701 : HS65_LH_OAI22X6 port map( A => n2730, B => n2444, C => n2442, D => 
                           n176, Z => n1866);
   U1702 : HS65_LH_OAI22X6 port map( A => n2732, B => n2444, C => n2442, D => 
                           n175, Z => n1867);
   U1703 : HS65_LH_OAI22X6 port map( A => n2734, B => n2444, C => n2442, D => 
                           n174, Z => n1868);
   U1704 : HS65_LH_OAI22X6 port map( A => n2736, B => n2444, C => n2441, D => 
                           n173, Z => n1869);
   U1705 : HS65_LH_OAI22X6 port map( A => n2738, B => n2444, C => n2441, D => 
                           n172, Z => n1870);
   U1706 : HS65_LH_OAI22X6 port map( A => n2740, B => n2444, C => n2441, D => 
                           n171, Z => n1871);
   U1707 : HS65_LH_OAI22X6 port map( A => n2742, B => n2444, C => n2441, D => 
                           n170, Z => n1872);
   U1708 : HS65_LH_OAI22X6 port map( A => n2744, B => n2444, C => n2441, D => 
                           n169, Z => n1873);
   U1709 : HS65_LH_OAI22X6 port map( A => n2746, B => n2444, C => n2441, D => 
                           n168, Z => n1874);
   U1710 : HS65_LH_OAI22X6 port map( A => n2748, B => n2444, C => n2441, D => 
                           n167, Z => n1875);
   U1711 : HS65_LH_OAI22X6 port map( A => n2750, B => n2444, C => n2441, D => 
                           n166, Z => n1876);
   U1712 : HS65_LH_OAI22X6 port map( A => n2752, B => n2444, C => n2441, D => 
                           n165, Z => n1877);
   U1713 : HS65_LH_OAI22X6 port map( A => n2754, B => n2444, C => n2441, D => 
                           n164, Z => n1878);
   U1714 : HS65_LH_OAI22X6 port map( A => n2756, B => n2444, C => n2441, D => 
                           n163, Z => n1879);
   U1715 : HS65_LH_OAI22X6 port map( A => n2758, B => n2444, C => n2441, D => 
                           n162, Z => n1880);
   U1716 : HS65_LH_OAI22X6 port map( A => n2724, B => n2439, C => n2437, D => 
                           n147, Z => n1895);
   U1717 : HS65_LH_OAI22X6 port map( A => n2726, B => n2439, C => n2437, D => 
                           n146, Z => n1896);
   U1718 : HS65_LH_OAI22X6 port map( A => n2728, B => n2439, C => n2437, D => 
                           n145, Z => n1897);
   U1719 : HS65_LH_OAI22X6 port map( A => n2730, B => n2439, C => n2437, D => 
                           n144, Z => n1898);
   U1720 : HS65_LH_OAI22X6 port map( A => n2732, B => n2439, C => n2437, D => 
                           n143, Z => n1899);
   U1721 : HS65_LH_OAI22X6 port map( A => n2734, B => n2439, C => n2437, D => 
                           n142, Z => n1900);
   U1722 : HS65_LH_OAI22X6 port map( A => n2736, B => n2439, C => n2436, D => 
                           n141, Z => n1901);
   U1723 : HS65_LH_OAI22X6 port map( A => n2738, B => n2439, C => n2436, D => 
                           n140, Z => n1902);
   U1724 : HS65_LH_OAI22X6 port map( A => n2740, B => n2439, C => n2436, D => 
                           n139, Z => n1903);
   U1725 : HS65_LH_OAI22X6 port map( A => n2742, B => n2439, C => n2436, D => 
                           n138, Z => n1904);
   U1726 : HS65_LH_OAI22X6 port map( A => n2744, B => n2439, C => n2436, D => 
                           n137, Z => n1905);
   U1727 : HS65_LH_OAI22X6 port map( A => n2746, B => n2439, C => n2436, D => 
                           n136, Z => n1906);
   U1728 : HS65_LH_OAI22X6 port map( A => n2748, B => n2439, C => n2436, D => 
                           n135, Z => n1907);
   U1729 : HS65_LH_OAI22X6 port map( A => n2750, B => n2439, C => n2436, D => 
                           n134, Z => n1908);
   U1730 : HS65_LH_OAI22X6 port map( A => n2752, B => n2439, C => n2436, D => 
                           n133, Z => n1909);
   U1731 : HS65_LH_OAI22X6 port map( A => n2754, B => n2439, C => n2436, D => 
                           n132, Z => n1910);
   U1732 : HS65_LH_OAI22X6 port map( A => n2756, B => n2439, C => n2436, D => 
                           n131, Z => n1911);
   U1733 : HS65_LH_OAI22X6 port map( A => n2758, B => n2439, C => n2436, D => 
                           n130, Z => n1912);
   U1734 : HS65_LH_OAI22X6 port map( A => n2724, B => n306, C => n304, D => n51
                           , Z => n2311);
   U1735 : HS65_LH_OAI22X6 port map( A => n2726, B => n306, C => n304, D => n50
                           , Z => n2312);
   U1736 : HS65_LH_OAI22X6 port map( A => n2728, B => n306, C => n304, D => n49
                           , Z => n2313);
   U1737 : HS65_LH_OAI22X6 port map( A => n2730, B => n306, C => n304, D => n48
                           , Z => n2314);
   U1738 : HS65_LH_OAI22X6 port map( A => n2732, B => n306, C => n304, D => n47
                           , Z => n2315);
   U1739 : HS65_LH_OAI22X6 port map( A => n2734, B => n306, C => n304, D => n46
                           , Z => n2316);
   U1740 : HS65_LH_OAI22X6 port map( A => n2736, B => n306, C => n303, D => n45
                           , Z => n2317);
   U1741 : HS65_LH_OAI22X6 port map( A => n2738, B => n306, C => n303, D => n44
                           , Z => n2318);
   U1742 : HS65_LH_OAI22X6 port map( A => n2740, B => n306, C => n303, D => n43
                           , Z => n2319);
   U1743 : HS65_LH_OAI22X6 port map( A => n2742, B => n306, C => n303, D => n42
                           , Z => n2320);
   U1744 : HS65_LH_OAI22X6 port map( A => n2744, B => n306, C => n303, D => n41
                           , Z => n2321);
   U1745 : HS65_LH_OAI22X6 port map( A => n2746, B => n306, C => n303, D => n40
                           , Z => n2322);
   U1746 : HS65_LH_OAI22X6 port map( A => n2748, B => n306, C => n303, D => n39
                           , Z => n2323);
   U1747 : HS65_LH_OAI22X6 port map( A => n2750, B => n306, C => n303, D => n38
                           , Z => n2324);
   U1748 : HS65_LH_OAI22X6 port map( A => n2752, B => n306, C => n303, D => n37
                           , Z => n2325);
   U1749 : HS65_LH_OAI22X6 port map( A => n2754, B => n306, C => n303, D => n36
                           , Z => n2326);
   U1750 : HS65_LH_OAI22X6 port map( A => n2756, B => n306, C => n303, D => n35
                           , Z => n2327);
   U1751 : HS65_LH_OAI22X6 port map( A => n2758, B => n306, C => n303, D => n34
                           , Z => n2328);
   U1752 : HS65_LH_OAI22X6 port map( A => n2724, B => n301, C => n299, D => n19
                           , Z => n2343);
   U1753 : HS65_LH_OAI22X6 port map( A => n2726, B => n301, C => n299, D => n18
                           , Z => n2344);
   U1754 : HS65_LH_OAI22X6 port map( A => n2728, B => n301, C => n299, D => n17
                           , Z => n2345);
   U1755 : HS65_LH_OAI22X6 port map( A => n2730, B => n301, C => n299, D => n16
                           , Z => n2346);
   U1756 : HS65_LH_OAI22X6 port map( A => n2732, B => n301, C => n299, D => n15
                           , Z => n2347);
   U1757 : HS65_LH_OAI22X6 port map( A => n2734, B => n301, C => n299, D => n14
                           , Z => n2348);
   U1758 : HS65_LH_OAI22X6 port map( A => n2736, B => n301, C => n298, D => n13
                           , Z => n2349);
   U1759 : HS65_LH_OAI22X6 port map( A => n2738, B => n301, C => n298, D => n12
                           , Z => n2350);
   U1760 : HS65_LH_OAI22X6 port map( A => n2740, B => n301, C => n298, D => n11
                           , Z => n2351);
   U1761 : HS65_LH_OAI22X6 port map( A => n2742, B => n301, C => n298, D => n10
                           , Z => n2352);
   U1762 : HS65_LH_OAI22X6 port map( A => n2744, B => n301, C => n298, D => n9,
                           Z => n2353);
   U1763 : HS65_LH_OAI22X6 port map( A => n2746, B => n301, C => n298, D => n8,
                           Z => n2354);
   U1764 : HS65_LH_OAI22X6 port map( A => n2748, B => n301, C => n298, D => n7,
                           Z => n2355);
   U1765 : HS65_LH_OAI22X6 port map( A => n2750, B => n301, C => n298, D => n6,
                           Z => n2356);
   U1766 : HS65_LH_OAI22X6 port map( A => n2752, B => n301, C => n298, D => n5,
                           Z => n2357);
   U1767 : HS65_LH_OAI22X6 port map( A => n2754, B => n301, C => n298, D => n4,
                           Z => n2358);
   U1768 : HS65_LH_OAI22X6 port map( A => n2756, B => n301, C => n298, D => n3,
                           Z => n2359);
   U1769 : HS65_LH_OAI22X6 port map( A => n2758, B => n301, C => n298, D => n2,
                           Z => n2360);
   U1770 : HS65_LH_OAI22X6 port map( A => n2724, B => n316, C => n314, D => 
                           n115, Z => n2247);
   U1771 : HS65_LH_OAI22X6 port map( A => n2726, B => n316, C => n314, D => 
                           n114, Z => n2248);
   U1772 : HS65_LH_OAI22X6 port map( A => n2728, B => n316, C => n314, D => 
                           n113, Z => n2249);
   U1773 : HS65_LH_OAI22X6 port map( A => n2730, B => n316, C => n314, D => 
                           n112, Z => n2250);
   U1774 : HS65_LH_OAI22X6 port map( A => n2732, B => n316, C => n314, D => 
                           n111, Z => n2251);
   U1775 : HS65_LH_OAI22X6 port map( A => n2734, B => n316, C => n314, D => 
                           n110, Z => n2252);
   U1776 : HS65_LH_OAI22X6 port map( A => n2736, B => n316, C => n313, D => 
                           n109, Z => n2253);
   U1777 : HS65_LH_OAI22X6 port map( A => n2738, B => n316, C => n313, D => 
                           n108, Z => n2254);
   U1778 : HS65_LH_OAI22X6 port map( A => n2740, B => n316, C => n313, D => 
                           n107, Z => n2255);
   U1779 : HS65_LH_OAI22X6 port map( A => n2742, B => n316, C => n313, D => 
                           n106, Z => n2256);
   U1780 : HS65_LH_OAI22X6 port map( A => n2744, B => n316, C => n313, D => 
                           n105, Z => n2257);
   U1781 : HS65_LH_OAI22X6 port map( A => n2746, B => n316, C => n313, D => 
                           n104, Z => n2258);
   U1782 : HS65_LH_OAI22X6 port map( A => n2748, B => n316, C => n313, D => 
                           n103, Z => n2259);
   U1783 : HS65_LH_OAI22X6 port map( A => n2750, B => n316, C => n313, D => 
                           n102, Z => n2260);
   U1784 : HS65_LH_OAI22X6 port map( A => n2752, B => n316, C => n313, D => 
                           n101, Z => n2261);
   U1785 : HS65_LH_OAI22X6 port map( A => n2754, B => n316, C => n313, D => 
                           n100, Z => n2262);
   U1786 : HS65_LH_OAI22X6 port map( A => n2756, B => n316, C => n313, D => n99
                           , Z => n2263);
   U1787 : HS65_LH_OAI22X6 port map( A => n2758, B => n316, C => n313, D => n98
                           , Z => n2264);
   U1788 : HS65_LH_OAI22X6 port map( A => n2724, B => n311, C => n309, D => n83
                           , Z => n2279);
   U1789 : HS65_LH_OAI22X6 port map( A => n2726, B => n311, C => n309, D => n82
                           , Z => n2280);
   U1790 : HS65_LH_OAI22X6 port map( A => n2728, B => n311, C => n309, D => n81
                           , Z => n2281);
   U1791 : HS65_LH_OAI22X6 port map( A => n2730, B => n311, C => n309, D => n80
                           , Z => n2282);
   U1792 : HS65_LH_OAI22X6 port map( A => n2732, B => n311, C => n309, D => n79
                           , Z => n2283);
   U1793 : HS65_LH_OAI22X6 port map( A => n2734, B => n311, C => n309, D => n78
                           , Z => n2284);
   U1794 : HS65_LH_OAI22X6 port map( A => n2736, B => n311, C => n308, D => n77
                           , Z => n2285);
   U1795 : HS65_LH_OAI22X6 port map( A => n2738, B => n311, C => n308, D => n76
                           , Z => n2286);
   U1796 : HS65_LH_OAI22X6 port map( A => n2740, B => n311, C => n308, D => n75
                           , Z => n2287);
   U1797 : HS65_LH_OAI22X6 port map( A => n2742, B => n311, C => n308, D => n74
                           , Z => n2288);
   U1798 : HS65_LH_OAI22X6 port map( A => n2744, B => n311, C => n308, D => n73
                           , Z => n2289);
   U1799 : HS65_LH_OAI22X6 port map( A => n2746, B => n311, C => n308, D => n72
                           , Z => n2290);
   U1800 : HS65_LH_OAI22X6 port map( A => n2748, B => n311, C => n308, D => n71
                           , Z => n2291);
   U1801 : HS65_LH_OAI22X6 port map( A => n2750, B => n311, C => n308, D => n70
                           , Z => n2292);
   U1802 : HS65_LH_OAI22X6 port map( A => n2752, B => n311, C => n308, D => n69
                           , Z => n2293);
   U1803 : HS65_LH_OAI22X6 port map( A => n2754, B => n311, C => n308, D => n68
                           , Z => n2294);
   U1804 : HS65_LH_OAI22X6 port map( A => n2756, B => n311, C => n308, D => n67
                           , Z => n2295);
   U1805 : HS65_LH_OAI22X6 port map( A => n2758, B => n311, C => n308, D => n66
                           , Z => n2296);
   U1806 : HS65_LH_OAI22X6 port map( A => n2698, B => n2475, C => n2472, D => 
                           n256, Z => n1658);
   U1807 : HS65_LH_OAI22X6 port map( A => n2700, B => n2475, C => n2471, D => 
                           n255, Z => n1659);
   U1808 : HS65_LH_OAI22X6 port map( A => n2702, B => n2475, C => n2472, D => 
                           n254, Z => n1660);
   U1809 : HS65_LH_OAI22X6 port map( A => n2704, B => n2475, C => n2471, D => 
                           n253, Z => n1661);
   U1810 : HS65_LH_OAI22X6 port map( A => n2706, B => n2475, C => n2472, D => 
                           n252, Z => n1662);
   U1811 : HS65_LH_OAI22X6 port map( A => n2708, B => n2475, C => n2471, D => 
                           n251, Z => n1663);
   U1812 : HS65_LH_OAI22X6 port map( A => n2710, B => n2475, C => n2472, D => 
                           n250, Z => n1664);
   U1813 : HS65_LH_OAI22X6 port map( A => n2712, B => n2475, C => n2472, D => 
                           n249, Z => n1665);
   U1814 : HS65_LH_OAI22X6 port map( A => n2714, B => n2475, C => n2472, D => 
                           n248, Z => n1666);
   U1815 : HS65_LH_OAI22X6 port map( A => n2716, B => n2475, C => n2472, D => 
                           n247, Z => n1667);
   U1816 : HS65_LH_OAI22X6 port map( A => n2718, B => n2475, C => n2472, D => 
                           n246, Z => n1668);
   U1817 : HS65_LH_OAI22X6 port map( A => n2720, B => n2475, C => n2472, D => 
                           n245, Z => n1669);
   U1818 : HS65_LH_OAI22X6 port map( A => n2722, B => n2475, C => n2472, D => 
                           n244, Z => n1670);
   U1819 : HS65_LH_OAI22X6 port map( A => n2698, B => n2470, C => n2467, D => 
                           n224, Z => n1690);
   U1820 : HS65_LH_OAI22X6 port map( A => n2700, B => n2470, C => n2466, D => 
                           n223, Z => n1691);
   U1821 : HS65_LH_OAI22X6 port map( A => n2702, B => n2470, C => n2467, D => 
                           n222, Z => n1692);
   U1822 : HS65_LH_OAI22X6 port map( A => n2704, B => n2470, C => n2466, D => 
                           n221, Z => n1693);
   U1823 : HS65_LH_OAI22X6 port map( A => n2706, B => n2470, C => n2467, D => 
                           n220, Z => n1694);
   U1824 : HS65_LH_OAI22X6 port map( A => n2708, B => n2470, C => n2466, D => 
                           n219, Z => n1695);
   U1825 : HS65_LH_OAI22X6 port map( A => n2710, B => n2470, C => n2467, D => 
                           n218, Z => n1696);
   U1826 : HS65_LH_OAI22X6 port map( A => n2712, B => n2470, C => n2467, D => 
                           n217, Z => n1697);
   U1827 : HS65_LH_OAI22X6 port map( A => n2714, B => n2470, C => n2467, D => 
                           n216, Z => n1698);
   U1828 : HS65_LH_OAI22X6 port map( A => n2716, B => n2470, C => n2467, D => 
                           n215, Z => n1699);
   U1829 : HS65_LH_OAI22X6 port map( A => n2718, B => n2470, C => n2467, D => 
                           n214, Z => n1700);
   U1830 : HS65_LH_OAI22X6 port map( A => n2720, B => n2470, C => n2467, D => 
                           n213, Z => n1701);
   U1831 : HS65_LH_OAI22X6 port map( A => n2722, B => n2470, C => n2467, D => 
                           n212, Z => n1702);
   U1832 : HS65_LH_OAI22X6 port map( A => n2698, B => n2445, C => n2442, D => 
                           n192, Z => n1850);
   U1833 : HS65_LH_OAI22X6 port map( A => n2700, B => n2445, C => n2441, D => 
                           n191, Z => n1851);
   U1834 : HS65_LH_OAI22X6 port map( A => n2702, B => n2445, C => n2442, D => 
                           n190, Z => n1852);
   U1835 : HS65_LH_OAI22X6 port map( A => n2704, B => n2445, C => n2441, D => 
                           n189, Z => n1853);
   U1836 : HS65_LH_OAI22X6 port map( A => n2706, B => n2445, C => n2442, D => 
                           n188, Z => n1854);
   U1837 : HS65_LH_OAI22X6 port map( A => n2708, B => n2445, C => n2441, D => 
                           n187, Z => n1855);
   U1838 : HS65_LH_OAI22X6 port map( A => n2710, B => n2445, C => n2442, D => 
                           n186, Z => n1856);
   U1839 : HS65_LH_OAI22X6 port map( A => n2712, B => n2445, C => n2442, D => 
                           n185, Z => n1857);
   U1840 : HS65_LH_OAI22X6 port map( A => n2714, B => n2445, C => n2442, D => 
                           n184, Z => n1858);
   U1841 : HS65_LH_OAI22X6 port map( A => n2716, B => n2445, C => n2442, D => 
                           n183, Z => n1859);
   U1842 : HS65_LH_OAI22X6 port map( A => n2718, B => n2445, C => n2442, D => 
                           n182, Z => n1860);
   U1843 : HS65_LH_OAI22X6 port map( A => n2720, B => n2445, C => n2442, D => 
                           n181, Z => n1861);
   U1844 : HS65_LH_OAI22X6 port map( A => n2722, B => n2445, C => n2442, D => 
                           n180, Z => n1862);
   U1845 : HS65_LH_OAI22X6 port map( A => n2698, B => n2440, C => n2437, D => 
                           n160, Z => n1882);
   U1846 : HS65_LH_OAI22X6 port map( A => n2700, B => n2440, C => n2436, D => 
                           n159, Z => n1883);
   U1847 : HS65_LH_OAI22X6 port map( A => n2702, B => n2440, C => n2437, D => 
                           n158, Z => n1884);
   U1848 : HS65_LH_OAI22X6 port map( A => n2704, B => n2440, C => n2436, D => 
                           n157, Z => n1885);
   U1849 : HS65_LH_OAI22X6 port map( A => n2706, B => n2440, C => n2437, D => 
                           n156, Z => n1886);
   U1850 : HS65_LH_OAI22X6 port map( A => n2708, B => n2440, C => n2436, D => 
                           n155, Z => n1887);
   U1851 : HS65_LH_OAI22X6 port map( A => n2710, B => n2440, C => n2437, D => 
                           n154, Z => n1888);
   U1852 : HS65_LH_OAI22X6 port map( A => n2712, B => n2440, C => n2437, D => 
                           n153, Z => n1889);
   U1853 : HS65_LH_OAI22X6 port map( A => n2714, B => n2440, C => n2437, D => 
                           n152, Z => n1890);
   U1854 : HS65_LH_OAI22X6 port map( A => n2716, B => n2440, C => n2437, D => 
                           n151, Z => n1891);
   U1855 : HS65_LH_OAI22X6 port map( A => n2718, B => n2440, C => n2437, D => 
                           n150, Z => n1892);
   U1856 : HS65_LH_OAI22X6 port map( A => n2720, B => n2440, C => n2437, D => 
                           n149, Z => n1893);
   U1857 : HS65_LH_OAI22X6 port map( A => n2722, B => n2440, C => n2437, D => 
                           n148, Z => n1894);
   U1858 : HS65_LH_OAI22X6 port map( A => n2698, B => n307, C => n304, D => n64
                           , Z => n2298);
   U1859 : HS65_LH_OAI22X6 port map( A => n2700, B => n307, C => n303, D => n63
                           , Z => n2299);
   U1860 : HS65_LH_OAI22X6 port map( A => n2702, B => n307, C => n304, D => n62
                           , Z => n2300);
   U1861 : HS65_LH_OAI22X6 port map( A => n2704, B => n307, C => n303, D => n61
                           , Z => n2301);
   U1862 : HS65_LH_OAI22X6 port map( A => n2706, B => n307, C => n304, D => n60
                           , Z => n2302);
   U1863 : HS65_LH_OAI22X6 port map( A => n2708, B => n307, C => n303, D => n59
                           , Z => n2303);
   U1864 : HS65_LH_OAI22X6 port map( A => n2710, B => n307, C => n304, D => n58
                           , Z => n2304);
   U1865 : HS65_LH_OAI22X6 port map( A => n2712, B => n307, C => n304, D => n57
                           , Z => n2305);
   U1866 : HS65_LH_OAI22X6 port map( A => n2714, B => n307, C => n304, D => n56
                           , Z => n2306);
   U1867 : HS65_LH_OAI22X6 port map( A => n2716, B => n307, C => n304, D => n55
                           , Z => n2307);
   U1868 : HS65_LH_OAI22X6 port map( A => n2718, B => n307, C => n304, D => n54
                           , Z => n2308);
   U1869 : HS65_LH_OAI22X6 port map( A => n2720, B => n307, C => n304, D => n53
                           , Z => n2309);
   U1870 : HS65_LH_OAI22X6 port map( A => n2722, B => n307, C => n304, D => n52
                           , Z => n2310);
   U1871 : HS65_LH_OAI22X6 port map( A => n2698, B => n302, C => n299, D => n32
                           , Z => n2330);
   U1872 : HS65_LH_OAI22X6 port map( A => n2700, B => n302, C => n298, D => n31
                           , Z => n2331);
   U1873 : HS65_LH_OAI22X6 port map( A => n2702, B => n302, C => n299, D => n30
                           , Z => n2332);
   U1874 : HS65_LH_OAI22X6 port map( A => n2704, B => n302, C => n298, D => n29
                           , Z => n2333);
   U1875 : HS65_LH_OAI22X6 port map( A => n2706, B => n302, C => n299, D => n28
                           , Z => n2334);
   U1876 : HS65_LH_OAI22X6 port map( A => n2708, B => n302, C => n298, D => n27
                           , Z => n2335);
   U1877 : HS65_LH_OAI22X6 port map( A => n2710, B => n302, C => n299, D => n26
                           , Z => n2336);
   U1878 : HS65_LH_OAI22X6 port map( A => n2712, B => n302, C => n299, D => n25
                           , Z => n2337);
   U1879 : HS65_LH_OAI22X6 port map( A => n2714, B => n302, C => n299, D => n24
                           , Z => n2338);
   U1880 : HS65_LH_OAI22X6 port map( A => n2716, B => n302, C => n299, D => n23
                           , Z => n2339);
   U1881 : HS65_LH_OAI22X6 port map( A => n2718, B => n302, C => n299, D => n22
                           , Z => n2340);
   U1882 : HS65_LH_OAI22X6 port map( A => n2720, B => n302, C => n299, D => n21
                           , Z => n2341);
   U1883 : HS65_LH_OAI22X6 port map( A => n2722, B => n302, C => n299, D => n20
                           , Z => n2342);
   U1884 : HS65_LH_OAI22X6 port map( A => n2698, B => n317, C => n314, D => 
                           n128, Z => n2234);
   U1885 : HS65_LH_OAI22X6 port map( A => n2700, B => n317, C => n313, D => 
                           n127, Z => n2235);
   U1886 : HS65_LH_OAI22X6 port map( A => n2702, B => n317, C => n314, D => 
                           n126, Z => n2236);
   U1887 : HS65_LH_OAI22X6 port map( A => n2704, B => n317, C => n313, D => 
                           n125, Z => n2237);
   U1888 : HS65_LH_OAI22X6 port map( A => n2706, B => n317, C => n314, D => 
                           n124, Z => n2238);
   U1889 : HS65_LH_OAI22X6 port map( A => n2708, B => n317, C => n313, D => 
                           n123, Z => n2239);
   U1890 : HS65_LH_OAI22X6 port map( A => n2710, B => n317, C => n314, D => 
                           n122, Z => n2240);
   U1891 : HS65_LH_OAI22X6 port map( A => n2712, B => n317, C => n314, D => 
                           n121, Z => n2241);
   U1892 : HS65_LH_OAI22X6 port map( A => n2714, B => n317, C => n314, D => 
                           n120, Z => n2242);
   U1893 : HS65_LH_OAI22X6 port map( A => n2716, B => n317, C => n314, D => 
                           n119, Z => n2243);
   U1894 : HS65_LH_OAI22X6 port map( A => n2718, B => n317, C => n314, D => 
                           n118, Z => n2244);
   U1895 : HS65_LH_OAI22X6 port map( A => n2720, B => n317, C => n314, D => 
                           n117, Z => n2245);
   U1896 : HS65_LH_OAI22X6 port map( A => n2722, B => n317, C => n314, D => 
                           n116, Z => n2246);
   U1897 : HS65_LH_OAI22X6 port map( A => n2698, B => n312, C => n309, D => n96
                           , Z => n2266);
   U1898 : HS65_LH_OAI22X6 port map( A => n2700, B => n312, C => n308, D => n95
                           , Z => n2267);
   U1899 : HS65_LH_OAI22X6 port map( A => n2702, B => n312, C => n309, D => n94
                           , Z => n2268);
   U1900 : HS65_LH_OAI22X6 port map( A => n2704, B => n312, C => n308, D => n93
                           , Z => n2269);
   U1901 : HS65_LH_OAI22X6 port map( A => n2706, B => n312, C => n309, D => n92
                           , Z => n2270);
   U1902 : HS65_LH_OAI22X6 port map( A => n2708, B => n312, C => n308, D => n91
                           , Z => n2271);
   U1903 : HS65_LH_OAI22X6 port map( A => n2710, B => n312, C => n309, D => n90
                           , Z => n2272);
   U1904 : HS65_LH_OAI22X6 port map( A => n2712, B => n312, C => n309, D => n89
                           , Z => n2273);
   U1905 : HS65_LH_OAI22X6 port map( A => n2714, B => n312, C => n309, D => n88
                           , Z => n2274);
   U1906 : HS65_LH_OAI22X6 port map( A => n2716, B => n312, C => n309, D => n87
                           , Z => n2275);
   U1907 : HS65_LH_OAI22X6 port map( A => n2718, B => n312, C => n309, D => n86
                           , Z => n2276);
   U1908 : HS65_LH_OAI22X6 port map( A => n2720, B => n312, C => n309, D => n85
                           , Z => n2277);
   U1909 : HS65_LH_OAI22X6 port map( A => n2722, B => n312, C => n309, D => n84
                           , Z => n2278);
   U1910 : HS65_LH_NAND3X5 port map( A => n2908, B => n2909, C => n2910, Z => 
                           n836);
   U1911 : HS65_LH_NAND2X7 port map( A => registers_1_0_port, B => n2670, Z => 
                           n2910);
   U1912 : HS65_LH_NAND2X7 port map( A => registers_3_0_port, B => n2664, Z => 
                           n2909);
   U1913 : HS65_LH_NAND2X7 port map( A => registers_2_0_port, B => n2667, Z => 
                           n2908);
   U1914 : HS65_LH_NAND3X5 port map( A => n2914, B => n2915, C => n2916, Z => 
                           n671);
   U1915 : HS65_LH_NAND2X7 port map( A => registers_1_1_port, B => n2670, Z => 
                           n2916);
   U1916 : HS65_LH_NAND2X7 port map( A => registers_3_1_port, B => n2664, Z => 
                           n2915);
   U1917 : HS65_LH_NAND2X7 port map( A => registers_2_1_port, B => n2667, Z => 
                           n2914);
   U1918 : HS65_LH_NAND3X5 port map( A => n2920, B => n2921, C => n2922, Z => 
                           n506);
   U1919 : HS65_LH_NAND2X7 port map( A => registers_1_2_port, B => n2670, Z => 
                           n2922);
   U1920 : HS65_LH_NAND2X7 port map( A => registers_3_2_port, B => n2664, Z => 
                           n2921);
   U1921 : HS65_LH_NAND2X7 port map( A => registers_2_2_port, B => n2667, Z => 
                           n2920);
   U1922 : HS65_LH_NAND3X5 port map( A => n2926, B => n2927, C => n2928, Z => 
                           n461);
   U1923 : HS65_LH_NAND2X7 port map( A => registers_1_3_port, B => n2670, Z => 
                           n2928);
   U1924 : HS65_LH_NAND2X7 port map( A => registers_3_3_port, B => n2664, Z => 
                           n2927);
   U1925 : HS65_LH_NAND2X7 port map( A => registers_2_3_port, B => n2667, Z => 
                           n2926);
   U1926 : HS65_LH_NAND3X5 port map( A => n2932, B => n2933, C => n2934, Z => 
                           n446);
   U1927 : HS65_LH_NAND2X7 port map( A => registers_1_4_port, B => n2670, Z => 
                           n2934);
   U1928 : HS65_LH_NAND2X7 port map( A => registers_3_4_port, B => n2664, Z => 
                           n2933);
   U1929 : HS65_LH_NAND2X7 port map( A => registers_2_4_port, B => n2667, Z => 
                           n2932);
   U1930 : HS65_LH_NAND3X5 port map( A => n2938, B => n2939, C => n2940, Z => 
                           n431);
   U1931 : HS65_LH_NAND2X7 port map( A => registers_1_5_port, B => n2670, Z => 
                           n2940);
   U1932 : HS65_LH_NAND2X7 port map( A => registers_3_5_port, B => n2664, Z => 
                           n2939);
   U1933 : HS65_LH_NAND2X7 port map( A => registers_2_5_port, B => n2667, Z => 
                           n2938);
   U1934 : HS65_LH_NAND3X5 port map( A => n2944, B => n2945, C => n2946, Z => 
                           n416);
   U1935 : HS65_LH_NAND2X7 port map( A => registers_1_6_port, B => n2670, Z => 
                           n2946);
   U1936 : HS65_LH_NAND2X7 port map( A => registers_3_6_port, B => n2664, Z => 
                           n2945);
   U1937 : HS65_LH_NAND2X7 port map( A => registers_2_6_port, B => n2667, Z => 
                           n2944);
   U1938 : HS65_LH_NAND3X5 port map( A => n2950, B => n2951, C => n2952, Z => 
                           n401);
   U1939 : HS65_LH_NAND2X7 port map( A => registers_1_7_port, B => n2670, Z => 
                           n2952);
   U1940 : HS65_LH_NAND2X7 port map( A => registers_3_7_port, B => n2664, Z => 
                           n2951);
   U1941 : HS65_LH_NAND2X7 port map( A => registers_2_7_port, B => n2667, Z => 
                           n2950);
   U1942 : HS65_LH_NAND3X5 port map( A => n2956, B => n2957, C => n2958, Z => 
                           n386);
   U1943 : HS65_LH_NAND2X7 port map( A => registers_1_8_port, B => n2670, Z => 
                           n2958);
   U1944 : HS65_LH_NAND2X7 port map( A => registers_3_8_port, B => n2664, Z => 
                           n2957);
   U1945 : HS65_LH_NAND2X7 port map( A => registers_2_8_port, B => n2667, Z => 
                           n2956);
   U1946 : HS65_LH_NAND3X5 port map( A => n2962, B => n2963, C => n2964, Z => 
                           n339);
   U1947 : HS65_LH_NAND2X7 port map( A => registers_1_9_port, B => n2670, Z => 
                           n2964);
   U1948 : HS65_LH_NAND2X7 port map( A => registers_3_9_port, B => n2664, Z => 
                           n2963);
   U1949 : HS65_LH_NAND2X7 port map( A => registers_2_9_port, B => n2667, Z => 
                           n2962);
   U1950 : HS65_LH_NAND3X5 port map( A => n2974, B => n2975, C => n2976, Z => 
                           n806);
   U1951 : HS65_LH_NAND2X7 port map( A => registers_1_11_port, B => n2670, Z =>
                           n2976);
   U1952 : HS65_LH_NAND2X7 port map( A => registers_3_11_port, B => n2664, Z =>
                           n2975);
   U1953 : HS65_LH_NAND2X7 port map( A => registers_2_11_port, B => n2667, Z =>
                           n2974);
   U1954 : HS65_LH_NAND3X5 port map( A => n2980, B => n2981, C => n2982, Z => 
                           n791);
   U1955 : HS65_LH_NAND2X7 port map( A => registers_1_12_port, B => n2671, Z =>
                           n2982);
   U1956 : HS65_LH_NAND2X7 port map( A => registers_3_12_port, B => n2665, Z =>
                           n2981);
   U1957 : HS65_LH_NAND2X7 port map( A => registers_2_12_port, B => n2668, Z =>
                           n2980);
   U1958 : HS65_LH_NAND3X5 port map( A => n2986, B => n2987, C => n2988, Z => 
                           n776);
   U1959 : HS65_LH_NAND2X7 port map( A => registers_1_13_port, B => n2671, Z =>
                           n2988);
   U1960 : HS65_LH_NAND2X7 port map( A => registers_3_13_port, B => n2665, Z =>
                           n2987);
   U1961 : HS65_LH_NAND2X7 port map( A => registers_2_13_port, B => n2668, Z =>
                           n2986);
   U1962 : HS65_LH_NAND3X5 port map( A => n2992, B => n2993, C => n2994, Z => 
                           n761);
   U1963 : HS65_LH_NAND2X7 port map( A => registers_1_14_port, B => n2671, Z =>
                           n2994);
   U1964 : HS65_LH_NAND2X7 port map( A => registers_3_14_port, B => n2665, Z =>
                           n2993);
   U1965 : HS65_LH_NAND2X7 port map( A => registers_2_14_port, B => n2668, Z =>
                           n2992);
   U1966 : HS65_LH_NAND3X5 port map( A => n2998, B => n2999, C => n3000, Z => 
                           n746);
   U1967 : HS65_LH_NAND2X7 port map( A => registers_1_15_port, B => n2671, Z =>
                           n3000);
   U1968 : HS65_LH_NAND2X7 port map( A => registers_3_15_port, B => n2665, Z =>
                           n2999);
   U1969 : HS65_LH_NAND2X7 port map( A => registers_2_15_port, B => n2668, Z =>
                           n2998);
   U1970 : HS65_LH_NAND3X5 port map( A => n3004, B => n3005, C => n3006, Z => 
                           n731);
   U1971 : HS65_LH_NAND2X7 port map( A => registers_1_16_port, B => n2671, Z =>
                           n3006);
   U1972 : HS65_LH_NAND2X7 port map( A => registers_3_16_port, B => n2665, Z =>
                           n3005);
   U1973 : HS65_LH_NAND2X7 port map( A => registers_2_16_port, B => n2668, Z =>
                           n3004);
   U1974 : HS65_LH_NAND3X5 port map( A => n3010, B => n3011, C => n3012, Z => 
                           n716);
   U1975 : HS65_LH_NAND2X7 port map( A => registers_1_17_port, B => n2671, Z =>
                           n3012);
   U1976 : HS65_LH_NAND2X7 port map( A => registers_3_17_port, B => n2665, Z =>
                           n3011);
   U1977 : HS65_LH_NAND2X7 port map( A => registers_2_17_port, B => n2668, Z =>
                           n3010);
   U1978 : HS65_LH_NAND3X5 port map( A => n3016, B => n3017, C => n3018, Z => 
                           n701);
   U1979 : HS65_LH_NAND2X7 port map( A => registers_1_18_port, B => n2671, Z =>
                           n3018);
   U1980 : HS65_LH_NAND2X7 port map( A => registers_3_18_port, B => n2665, Z =>
                           n3017);
   U1981 : HS65_LH_NAND2X7 port map( A => registers_2_18_port, B => n2668, Z =>
                           n3016);
   U1982 : HS65_LH_NAND3X5 port map( A => n3022, B => n3023, C => n3024, Z => 
                           n686);
   U1983 : HS65_LH_NAND2X7 port map( A => registers_1_19_port, B => n2671, Z =>
                           n3024);
   U1984 : HS65_LH_NAND2X7 port map( A => registers_3_19_port, B => n2665, Z =>
                           n3023);
   U1985 : HS65_LH_NAND2X7 port map( A => registers_2_19_port, B => n2668, Z =>
                           n3022);
   U1986 : HS65_LH_NAND3X5 port map( A => n3028, B => n3029, C => n3030, Z => 
                           n656);
   U1987 : HS65_LH_NAND2X7 port map( A => registers_1_20_port, B => n2671, Z =>
                           n3030);
   U1988 : HS65_LH_NAND2X7 port map( A => registers_3_20_port, B => n2665, Z =>
                           n3029);
   U1989 : HS65_LH_NAND2X7 port map( A => registers_2_20_port, B => n2668, Z =>
                           n3028);
   U1990 : HS65_LH_NAND3X5 port map( A => n3034, B => n3035, C => n3036, Z => 
                           n641);
   U1991 : HS65_LH_NAND2X7 port map( A => registers_1_21_port, B => n2671, Z =>
                           n3036);
   U1992 : HS65_LH_NAND2X7 port map( A => registers_3_21_port, B => n2665, Z =>
                           n3035);
   U1993 : HS65_LH_NAND2X7 port map( A => registers_2_21_port, B => n2668, Z =>
                           n3034);
   U1994 : HS65_LH_NAND3X5 port map( A => n3040, B => n3041, C => n3042, Z => 
                           n626);
   U1995 : HS65_LH_NAND2X7 port map( A => registers_1_22_port, B => n2671, Z =>
                           n3042);
   U1996 : HS65_LH_NAND2X7 port map( A => registers_3_22_port, B => n2665, Z =>
                           n3041);
   U1997 : HS65_LH_NAND2X7 port map( A => registers_2_22_port, B => n2668, Z =>
                           n3040);
   U1998 : HS65_LH_NAND3X5 port map( A => n3046, B => n3047, C => n3048, Z => 
                           n611);
   U1999 : HS65_LH_NAND2X7 port map( A => registers_1_23_port, B => n2671, Z =>
                           n3048);
   U2000 : HS65_LH_NAND2X7 port map( A => registers_3_23_port, B => n2665, Z =>
                           n3047);
   U2001 : HS65_LH_NAND2X7 port map( A => registers_2_23_port, B => n2668, Z =>
                           n3046);
   U2002 : HS65_LH_NAND3X5 port map( A => n3052, B => n3053, C => n3054, Z => 
                           n596);
   U2003 : HS65_LH_NAND2X7 port map( A => registers_1_24_port, B => n2672, Z =>
                           n3054);
   U2004 : HS65_LH_NAND2X7 port map( A => registers_3_24_port, B => n2666, Z =>
                           n3053);
   U2005 : HS65_LH_NAND2X7 port map( A => registers_2_24_port, B => n2669, Z =>
                           n3052);
   U2006 : HS65_LH_NAND3X5 port map( A => n3058, B => n3059, C => n3060, Z => 
                           n581);
   U2007 : HS65_LH_NAND2X7 port map( A => registers_1_25_port, B => n2672, Z =>
                           n3060);
   U2008 : HS65_LH_NAND2X7 port map( A => registers_3_25_port, B => n2666, Z =>
                           n3059);
   U2009 : HS65_LH_NAND2X7 port map( A => registers_2_25_port, B => n2669, Z =>
                           n3058);
   U2010 : HS65_LH_NAND3X5 port map( A => n3064, B => n3065, C => n3066, Z => 
                           n566);
   U2011 : HS65_LH_NAND2X7 port map( A => registers_1_26_port, B => n2672, Z =>
                           n3066);
   U2012 : HS65_LH_NAND2X7 port map( A => registers_3_26_port, B => n2666, Z =>
                           n3065);
   U2013 : HS65_LH_NAND2X7 port map( A => registers_2_26_port, B => n2669, Z =>
                           n3064);
   U2014 : HS65_LH_NAND3X5 port map( A => n3070, B => n3071, C => n3072, Z => 
                           n551);
   U2015 : HS65_LH_NAND2X7 port map( A => registers_1_27_port, B => n2672, Z =>
                           n3072);
   U2016 : HS65_LH_NAND2X7 port map( A => registers_3_27_port, B => n2666, Z =>
                           n3071);
   U2017 : HS65_LH_NAND2X7 port map( A => registers_2_27_port, B => n2669, Z =>
                           n3070);
   U2018 : HS65_LH_NAND3X5 port map( A => n3076, B => n3077, C => n3078, Z => 
                           n536);
   U2019 : HS65_LH_NAND2X7 port map( A => registers_1_28_port, B => n2672, Z =>
                           n3078);
   U2020 : HS65_LH_NAND2X7 port map( A => registers_3_28_port, B => n2666, Z =>
                           n3077);
   U2021 : HS65_LH_NAND2X7 port map( A => registers_2_28_port, B => n2669, Z =>
                           n3076);
   U2022 : HS65_LH_NAND3X5 port map( A => n3082, B => n3083, C => n3084, Z => 
                           n521);
   U2023 : HS65_LH_NAND2X7 port map( A => registers_1_29_port, B => n2672, Z =>
                           n3084);
   U2024 : HS65_LH_NAND2X7 port map( A => registers_3_29_port, B => n2666, Z =>
                           n3083);
   U2025 : HS65_LH_NAND2X7 port map( A => registers_2_29_port, B => n2669, Z =>
                           n3082);
   U2026 : HS65_LH_NAND3X5 port map( A => n3088, B => n3089, C => n3090, Z => 
                           n491);
   U2027 : HS65_LH_NAND2X7 port map( A => registers_1_30_port, B => n2672, Z =>
                           n3090);
   U2028 : HS65_LH_NAND2X7 port map( A => registers_3_30_port, B => n2666, Z =>
                           n3089);
   U2029 : HS65_LH_NAND2X7 port map( A => registers_2_30_port, B => n2669, Z =>
                           n3088);
   U2030 : HS65_LH_NAND3X5 port map( A => n3094, B => n3095, C => n3096, Z => 
                           n476);
   U2031 : HS65_LH_NAND2X7 port map( A => registers_1_31_port, B => n2672, Z =>
                           n3096);
   U2032 : HS65_LH_NAND2X7 port map( A => registers_3_31_port, B => n2666, Z =>
                           n3095);
   U2033 : HS65_LH_NAND2X7 port map( A => registers_2_31_port, B => n2669, Z =>
                           n3094);
   U2034 : HS65_LH_NAND3X5 port map( A => n2911, B => n2912, C => n2913, Z => 
                           n1364);
   U2035 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_0_port, Z => 
                           n2913);
   U2036 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_0_port, Z => 
                           n2912);
   U2037 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_0_port, Z => 
                           n2911);
   U2038 : HS65_LH_NAND3X5 port map( A => n2917, B => n2918, C => n2919, Z => 
                           n1199);
   U2039 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_1_port, Z => 
                           n2919);
   U2040 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_1_port, Z => 
                           n2918);
   U2041 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_1_port, Z => 
                           n2917);
   U2042 : HS65_LH_NAND3X5 port map( A => n2923, B => n2924, C => n2925, Z => 
                           n1034);
   U2043 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_2_port, Z => 
                           n2925);
   U2044 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_2_port, Z => 
                           n2924);
   U2045 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_2_port, Z => 
                           n2923);
   U2046 : HS65_LH_NAND3X5 port map( A => n2929, B => n2930, C => n2931, Z => 
                           n989);
   U2047 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_3_port, Z => 
                           n2931);
   U2048 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_3_port, Z => 
                           n2930);
   U2049 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_3_port, Z => 
                           n2929);
   U2050 : HS65_LH_NAND3X5 port map( A => n2935, B => n2936, C => n2937, Z => 
                           n974);
   U2051 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_4_port, Z => 
                           n2937);
   U2052 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_4_port, Z => 
                           n2936);
   U2053 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_4_port, Z => 
                           n2935);
   U2054 : HS65_LH_NAND3X5 port map( A => n2941, B => n2942, C => n2943, Z => 
                           n959);
   U2055 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_5_port, Z => 
                           n2943);
   U2056 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_5_port, Z => 
                           n2942);
   U2057 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_5_port, Z => 
                           n2941);
   U2058 : HS65_LH_NAND3X5 port map( A => n2947, B => n2948, C => n2949, Z => 
                           n944);
   U2059 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_6_port, Z => 
                           n2949);
   U2060 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_6_port, Z => 
                           n2948);
   U2061 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_6_port, Z => 
                           n2947);
   U2062 : HS65_LH_NAND3X5 port map( A => n2953, B => n2954, C => n2955, Z => 
                           n929);
   U2063 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_7_port, Z => 
                           n2955);
   U2064 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_7_port, Z => 
                           n2954);
   U2065 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_7_port, Z => 
                           n2953);
   U2066 : HS65_LH_NAND3X5 port map( A => n2959, B => n2960, C => n2961, Z => 
                           n914);
   U2067 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_8_port, Z => 
                           n2961);
   U2068 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_8_port, Z => 
                           n2960);
   U2069 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_8_port, Z => 
                           n2959);
   U2070 : HS65_LH_NAND3X5 port map( A => n2965, B => n2966, C => n2967, Z => 
                           n867);
   U2071 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_9_port, Z => 
                           n2967);
   U2072 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_9_port, Z => 
                           n2966);
   U2073 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_9_port, Z => 
                           n2965);
   U2074 : HS65_LH_NAND3X5 port map( A => n2971, B => n2972, C => n2973, Z => 
                           n1349);
   U2075 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_10_port, Z =>
                           n2973);
   U2076 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_10_port, Z =>
                           n2972);
   U2077 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_10_port, Z =>
                           n2971);
   U2078 : HS65_LH_NAND3X5 port map( A => n2977, B => n2978, C => n2979, Z => 
                           n1334);
   U2079 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_11_port, Z =>
                           n2979);
   U2080 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_11_port, Z =>
                           n2978);
   U2081 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_11_port, Z =>
                           n2977);
   U2082 : HS65_LH_NAND3X5 port map( A => n2983, B => n2984, C => n2985, Z => 
                           n1319);
   U2083 : HS65_LH_NAND2X7 port map( A => n2577, B => registers_1_12_port, Z =>
                           n2985);
   U2084 : HS65_LH_NAND2X7 port map( A => n2571, B => registers_3_12_port, Z =>
                           n2984);
   U2085 : HS65_LH_NAND2X7 port map( A => n2574, B => registers_2_12_port, Z =>
                           n2983);
   U2086 : HS65_LH_NAND3X5 port map( A => n2989, B => n2990, C => n2991, Z => 
                           n1304);
   U2087 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_13_port, Z =>
                           n2991);
   U2088 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_13_port, Z =>
                           n2990);
   U2089 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_13_port, Z =>
                           n2989);
   U2090 : HS65_LH_NAND3X5 port map( A => n2995, B => n2996, C => n2997, Z => 
                           n1289);
   U2091 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_14_port, Z =>
                           n2997);
   U2092 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_14_port, Z =>
                           n2996);
   U2093 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_14_port, Z =>
                           n2995);
   U2094 : HS65_LH_NAND3X5 port map( A => n3001, B => n3002, C => n3003, Z => 
                           n1274);
   U2095 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_15_port, Z =>
                           n3003);
   U2096 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_15_port, Z =>
                           n3002);
   U2097 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_15_port, Z =>
                           n3001);
   U2098 : HS65_LH_NAND3X5 port map( A => n3007, B => n3008, C => n3009, Z => 
                           n1259);
   U2099 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_16_port, Z =>
                           n3009);
   U2100 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_16_port, Z =>
                           n3008);
   U2101 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_16_port, Z =>
                           n3007);
   U2102 : HS65_LH_NAND3X5 port map( A => n3013, B => n3014, C => n3015, Z => 
                           n1244);
   U2103 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_17_port, Z =>
                           n3015);
   U2104 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_17_port, Z =>
                           n3014);
   U2105 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_17_port, Z =>
                           n3013);
   U2106 : HS65_LH_NAND3X5 port map( A => n3019, B => n3020, C => n3021, Z => 
                           n1229);
   U2107 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_18_port, Z =>
                           n3021);
   U2108 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_18_port, Z =>
                           n3020);
   U2109 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_18_port, Z =>
                           n3019);
   U2110 : HS65_LH_NAND3X5 port map( A => n3025, B => n3026, C => n3027, Z => 
                           n1214);
   U2111 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_19_port, Z =>
                           n3027);
   U2112 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_19_port, Z =>
                           n3026);
   U2113 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_19_port, Z =>
                           n3025);
   U2114 : HS65_LH_NAND3X5 port map( A => n3031, B => n3032, C => n3033, Z => 
                           n1184);
   U2115 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_20_port, Z =>
                           n3033);
   U2116 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_20_port, Z =>
                           n3032);
   U2117 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_20_port, Z =>
                           n3031);
   U2118 : HS65_LH_NAND3X5 port map( A => n3037, B => n3038, C => n3039, Z => 
                           n1169);
   U2119 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_21_port, Z =>
                           n3039);
   U2120 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_21_port, Z =>
                           n3038);
   U2121 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_21_port, Z =>
                           n3037);
   U2122 : HS65_LH_NAND3X5 port map( A => n3043, B => n3044, C => n3045, Z => 
                           n1154);
   U2123 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_22_port, Z =>
                           n3045);
   U2124 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_22_port, Z =>
                           n3044);
   U2125 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_22_port, Z =>
                           n3043);
   U2126 : HS65_LH_NAND3X5 port map( A => n3049, B => n3050, C => n3051, Z => 
                           n1139);
   U2127 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_23_port, Z =>
                           n3051);
   U2128 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_23_port, Z =>
                           n3050);
   U2129 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_23_port, Z =>
                           n3049);
   U2130 : HS65_LH_NAND3X5 port map( A => n3055, B => n3056, C => n3057, Z => 
                           n1124);
   U2131 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_24_port, Z =>
                           n3057);
   U2132 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_24_port, Z =>
                           n3056);
   U2133 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_24_port, Z =>
                           n3055);
   U2134 : HS65_LH_NAND3X5 port map( A => n3061, B => n3062, C => n3063, Z => 
                           n1109);
   U2135 : HS65_LH_NAND2X7 port map( A => n2578, B => registers_1_25_port, Z =>
                           n3063);
   U2136 : HS65_LH_NAND2X7 port map( A => n2572, B => registers_3_25_port, Z =>
                           n3062);
   U2137 : HS65_LH_NAND2X7 port map( A => n2575, B => registers_2_25_port, Z =>
                           n3061);
   U2138 : HS65_LH_NAND3X5 port map( A => n3067, B => n3068, C => n3069, Z => 
                           n1094);
   U2139 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_26_port, Z =>
                           n3069);
   U2140 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_26_port, Z =>
                           n3068);
   U2141 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_26_port, Z =>
                           n3067);
   U2142 : HS65_LH_NAND3X5 port map( A => n3073, B => n3074, C => n3075, Z => 
                           n1079);
   U2143 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_27_port, Z =>
                           n3075);
   U2144 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_27_port, Z =>
                           n3074);
   U2145 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_27_port, Z =>
                           n3073);
   U2146 : HS65_LH_NAND3X5 port map( A => n3079, B => n3080, C => n3081, Z => 
                           n1064);
   U2147 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_28_port, Z =>
                           n3081);
   U2148 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_28_port, Z =>
                           n3080);
   U2149 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_28_port, Z =>
                           n3079);
   U2150 : HS65_LH_NAND3X5 port map( A => n3085, B => n3086, C => n3087, Z => 
                           n1049);
   U2151 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_29_port, Z =>
                           n3087);
   U2152 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_29_port, Z =>
                           n3086);
   U2153 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_29_port, Z =>
                           n3085);
   U2154 : HS65_LH_NAND3X5 port map( A => n3091, B => n3092, C => n3093, Z => 
                           n1019);
   U2155 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_30_port, Z =>
                           n3093);
   U2156 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_30_port, Z =>
                           n3092);
   U2157 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_30_port, Z =>
                           n3091);
   U2158 : HS65_LH_NAND3X5 port map( A => n3097, B => n3098, C => n3099, Z => 
                           n1004);
   U2159 : HS65_LH_NAND2X7 port map( A => n2579, B => registers_1_31_port, Z =>
                           n3099);
   U2160 : HS65_LH_NAND2X7 port map( A => n2573, B => registers_3_31_port, Z =>
                           n3098);
   U2161 : HS65_LH_NAND2X7 port map( A => n2576, B => registers_2_31_port, Z =>
                           n3097);
   U2162 : HS65_LH_NAND2X7 port map( A => registers_2_10_port, B => n2667, Z =>
                           n2968);
   U2163 : HS65_LH_NAND2X7 port map( A => registers_3_10_port, B => n2664, Z =>
                           n2969);
   U2164 : HS65_LH_NAND2X7 port map( A => registers_1_10_port, B => n2670, Z =>
                           n2970);
   U2165 : HS65_LH_AO22X9 port map( A => n2697, B => n2510, C => n2507, D => 
                           registers_1_0_port, Z => n1434);
   U2166 : HS65_LH_AO22X9 port map( A => n2699, B => n2510, C => n2506, D => 
                           registers_1_1_port, Z => n1435);
   U2167 : HS65_LH_AO22X9 port map( A => n2701, B => n2510, C => n2507, D => 
                           registers_1_2_port, Z => n1436);
   U2168 : HS65_LH_AO22X9 port map( A => n2703, B => n2510, C => n2506, D => 
                           registers_1_3_port, Z => n1437);
   U2169 : HS65_LH_AO22X9 port map( A => n2705, B => n2510, C => n2507, D => 
                           registers_1_4_port, Z => n1438);
   U2170 : HS65_LH_AO22X9 port map( A => n2707, B => n2510, C => n2506, D => 
                           registers_1_5_port, Z => n1439);
   U2171 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2510, C => n2507, 
                           D => registers_1_6_port, Z => n1440);
   U2172 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2510, C => n2507,
                           D => registers_1_7_port, Z => n1441);
   U2173 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2510, C => n2507,
                           D => registers_1_8_port, Z => n1442);
   U2174 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2510, C => n2507,
                           D => registers_1_9_port, Z => n1443);
   U2175 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2510, C => n2507,
                           D => registers_1_10_port, Z => n1444);
   U2176 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2509, C => n2507,
                           D => registers_1_11_port, Z => n1445);
   U2177 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2509, C => n2507,
                           D => registers_1_12_port, Z => n1446);
   U2178 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2509, C => n2507,
                           D => registers_1_13_port, Z => n1447);
   U2179 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2509, C => n2507,
                           D => registers_1_14_port, Z => n1448);
   U2180 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2509, C => n2507,
                           D => registers_1_15_port, Z => n1449);
   U2181 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2509, C => n2507,
                           D => registers_1_16_port, Z => n1450);
   U2182 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2509, C => n2507,
                           D => registers_1_17_port, Z => n1451);
   U2183 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2509, C => n2507,
                           D => registers_1_18_port, Z => n1452);
   U2184 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2509, C => n2506,
                           D => registers_1_19_port, Z => n1453);
   U2185 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2509, C => n2506,
                           D => registers_1_20_port, Z => n1454);
   U2186 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2509, C => n2506,
                           D => registers_1_21_port, Z => n1455);
   U2187 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2509, C => n2506,
                           D => registers_1_22_port, Z => n1456);
   U2188 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2509, C => n2506,
                           D => registers_1_23_port, Z => n1457);
   U2189 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2509, C => n2506,
                           D => registers_1_24_port, Z => n1458);
   U2190 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2509, C => n2506,
                           D => registers_1_25_port, Z => n1459);
   U2191 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2509, C => n2506,
                           D => registers_1_26_port, Z => n1460);
   U2192 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2509, C => n2506,
                           D => registers_1_27_port, Z => n1461);
   U2193 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2509, C => n2506,
                           D => registers_1_28_port, Z => n1462);
   U2194 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2509, C => n2506,
                           D => registers_1_29_port, Z => n1463);
   U2195 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2509, C => n2506,
                           D => registers_1_30_port, Z => n1464);
   U2196 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2508, C => n2506,
                           D => registers_1_31_port, Z => n1465);
   U2197 : HS65_LH_AO22X9 port map( A => n2697, B => n2505, C => n2502, D => 
                           registers_2_0_port, Z => n1466);
   U2198 : HS65_LH_AO22X9 port map( A => n2699, B => n2505, C => n2501, D => 
                           registers_2_1_port, Z => n1467);
   U2199 : HS65_LH_AO22X9 port map( A => n2701, B => n2505, C => n2502, D => 
                           registers_2_2_port, Z => n1468);
   U2200 : HS65_LH_AO22X9 port map( A => n2703, B => n2505, C => n2501, D => 
                           registers_2_3_port, Z => n1469);
   U2201 : HS65_LH_AO22X9 port map( A => n2705, B => n2505, C => n2502, D => 
                           registers_2_4_port, Z => n1470);
   U2202 : HS65_LH_AO22X9 port map( A => n2707, B => n2505, C => n2501, D => 
                           registers_2_5_port, Z => n1471);
   U2203 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2505, C => n2502, 
                           D => registers_2_6_port, Z => n1472);
   U2204 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2505, C => n2502,
                           D => registers_2_7_port, Z => n1473);
   U2205 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2505, C => n2502,
                           D => registers_2_8_port, Z => n1474);
   U2206 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2505, C => n2502,
                           D => registers_2_9_port, Z => n1475);
   U2207 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2505, C => n2502,
                           D => registers_2_10_port, Z => n1476);
   U2208 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2504, C => n2502,
                           D => registers_2_11_port, Z => n1477);
   U2209 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2504, C => n2502,
                           D => registers_2_12_port, Z => n1478);
   U2210 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2504, C => n2502,
                           D => registers_2_13_port, Z => n1479);
   U2211 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2504, C => n2502,
                           D => registers_2_14_port, Z => n1480);
   U2212 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2504, C => n2502,
                           D => registers_2_15_port, Z => n1481);
   U2213 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2504, C => n2502,
                           D => registers_2_16_port, Z => n1482);
   U2214 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2504, C => n2502,
                           D => registers_2_17_port, Z => n1483);
   U2215 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2504, C => n2502,
                           D => registers_2_18_port, Z => n1484);
   U2216 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2504, C => n2501,
                           D => registers_2_19_port, Z => n1485);
   U2217 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2504, C => n2501,
                           D => registers_2_20_port, Z => n1486);
   U2218 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2504, C => n2501,
                           D => registers_2_21_port, Z => n1487);
   U2219 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2504, C => n2501,
                           D => registers_2_22_port, Z => n1488);
   U2220 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2504, C => n2501,
                           D => registers_2_23_port, Z => n1489);
   U2221 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2504, C => n2501,
                           D => registers_2_24_port, Z => n1490);
   U2222 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2504, C => n2501,
                           D => registers_2_25_port, Z => n1491);
   U2223 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2504, C => n2501,
                           D => registers_2_26_port, Z => n1492);
   U2224 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2504, C => n2501,
                           D => registers_2_27_port, Z => n1493);
   U2225 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2504, C => n2501,
                           D => registers_2_28_port, Z => n1494);
   U2226 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2504, C => n2501,
                           D => registers_2_29_port, Z => n1495);
   U2227 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2504, C => n2501,
                           D => registers_2_30_port, Z => n1496);
   U2228 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2503, C => n2501,
                           D => registers_2_31_port, Z => n1497);
   U2229 : HS65_LH_AO22X9 port map( A => n2697, B => n2500, C => n2497, D => 
                           registers_3_0_port, Z => n1498);
   U2230 : HS65_LH_AO22X9 port map( A => n2699, B => n2500, C => n2496, D => 
                           registers_3_1_port, Z => n1499);
   U2231 : HS65_LH_AO22X9 port map( A => n2701, B => n2500, C => n2497, D => 
                           registers_3_2_port, Z => n1500);
   U2232 : HS65_LH_AO22X9 port map( A => n2703, B => n2500, C => n2496, D => 
                           registers_3_3_port, Z => n1501);
   U2233 : HS65_LH_AO22X9 port map( A => n2705, B => n2500, C => n2497, D => 
                           registers_3_4_port, Z => n1502);
   U2234 : HS65_LH_AO22X9 port map( A => n2707, B => n2500, C => n2496, D => 
                           registers_3_5_port, Z => n1503);
   U2235 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2500, C => n2497, 
                           D => registers_3_6_port, Z => n1504);
   U2236 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2500, C => n2497,
                           D => registers_3_7_port, Z => n1505);
   U2237 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2500, C => n2497,
                           D => registers_3_8_port, Z => n1506);
   U2238 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2500, C => n2497,
                           D => registers_3_9_port, Z => n1507);
   U2239 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2500, C => n2497,
                           D => registers_3_10_port, Z => n1508);
   U2240 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2499, C => n2497,
                           D => registers_3_11_port, Z => n1509);
   U2241 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2499, C => n2497,
                           D => registers_3_12_port, Z => n1510);
   U2242 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2499, C => n2497,
                           D => registers_3_13_port, Z => n1511);
   U2243 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2499, C => n2497,
                           D => registers_3_14_port, Z => n1512);
   U2244 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2499, C => n2497,
                           D => registers_3_15_port, Z => n1513);
   U2245 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2499, C => n2497,
                           D => registers_3_16_port, Z => n1514);
   U2246 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2499, C => n2497,
                           D => registers_3_17_port, Z => n1515);
   U2247 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2499, C => n2497,
                           D => registers_3_18_port, Z => n1516);
   U2248 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2499, C => n2496,
                           D => registers_3_19_port, Z => n1517);
   U2249 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2499, C => n2496,
                           D => registers_3_20_port, Z => n1518);
   U2250 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2499, C => n2496,
                           D => registers_3_21_port, Z => n1519);
   U2251 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2499, C => n2496,
                           D => registers_3_22_port, Z => n1520);
   U2252 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2499, C => n2496,
                           D => registers_3_23_port, Z => n1521);
   U2253 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2499, C => n2496,
                           D => registers_3_24_port, Z => n1522);
   U2254 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2499, C => n2496,
                           D => registers_3_25_port, Z => n1523);
   U2255 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2499, C => n2496,
                           D => registers_3_26_port, Z => n1524);
   U2256 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2499, C => n2496,
                           D => registers_3_27_port, Z => n1525);
   U2257 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2499, C => n2496,
                           D => registers_3_28_port, Z => n1526);
   U2258 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2499, C => n2496,
                           D => registers_3_29_port, Z => n1527);
   U2259 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2499, C => n2496,
                           D => registers_3_30_port, Z => n1528);
   U2260 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2498, C => n2496,
                           D => registers_3_31_port, Z => n1529);
   U2261 : HS65_LH_AO22X9 port map( A => n2697, B => n2460, C => n2457, D => 
                           registers_11_0_port, Z => n1754);
   U2262 : HS65_LH_AO22X9 port map( A => n2699, B => n2460, C => n2456, D => 
                           registers_11_1_port, Z => n1755);
   U2263 : HS65_LH_AO22X9 port map( A => n2701, B => n2460, C => n2457, D => 
                           registers_11_2_port, Z => n1756);
   U2264 : HS65_LH_AO22X9 port map( A => n2703, B => n2460, C => n2456, D => 
                           registers_11_3_port, Z => n1757);
   U2265 : HS65_LH_AO22X9 port map( A => n2705, B => n2460, C => n2457, D => 
                           registers_11_4_port, Z => n1758);
   U2266 : HS65_LH_AO22X9 port map( A => n2707, B => n2460, C => n2456, D => 
                           registers_11_5_port, Z => n1759);
   U2267 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2460, C => n2457, 
                           D => registers_11_6_port, Z => n1760);
   U2268 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2460, C => n2457,
                           D => registers_11_7_port, Z => n1761);
   U2269 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2460, C => n2457,
                           D => registers_11_8_port, Z => n1762);
   U2270 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2460, C => n2457,
                           D => registers_11_9_port, Z => n1763);
   U2271 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2460, C => n2457,
                           D => registers_11_10_port, Z => n1764);
   U2272 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2459, C => n2457,
                           D => registers_11_11_port, Z => n1765);
   U2273 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2459, C => n2457,
                           D => registers_11_12_port, Z => n1766);
   U2274 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2459, C => n2457,
                           D => registers_11_13_port, Z => n1767);
   U2275 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2459, C => n2457,
                           D => registers_11_14_port, Z => n1768);
   U2276 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2459, C => n2457,
                           D => registers_11_15_port, Z => n1769);
   U2277 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2459, C => n2457,
                           D => registers_11_16_port, Z => n1770);
   U2278 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2459, C => n2457,
                           D => registers_11_17_port, Z => n1771);
   U2279 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2459, C => n2457,
                           D => registers_11_18_port, Z => n1772);
   U2280 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2459, C => n2456,
                           D => registers_11_19_port, Z => n1773);
   U2281 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2459, C => n2456,
                           D => registers_11_20_port, Z => n1774);
   U2282 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2459, C => n2456,
                           D => registers_11_21_port, Z => n1775);
   U2283 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2459, C => n2456,
                           D => registers_11_22_port, Z => n1776);
   U2284 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2459, C => n2456,
                           D => registers_11_23_port, Z => n1777);
   U2285 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2459, C => n2456,
                           D => registers_11_24_port, Z => n1778);
   U2286 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2459, C => n2456,
                           D => registers_11_25_port, Z => n1779);
   U2287 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2459, C => n2456,
                           D => registers_11_26_port, Z => n1780);
   U2288 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2459, C => n2456,
                           D => registers_11_27_port, Z => n1781);
   U2289 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2459, C => n2456,
                           D => registers_11_28_port, Z => n1782);
   U2290 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2459, C => n2456,
                           D => registers_11_29_port, Z => n1783);
   U2291 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2459, C => n2456,
                           D => registers_11_30_port, Z => n1784);
   U2292 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2458, C => n2456,
                           D => registers_11_31_port, Z => n1785);
   U2293 : HS65_LH_AO22X9 port map( A => n2697, B => n2450, C => n2447, D => 
                           registers_13_0_port, Z => n1818);
   U2294 : HS65_LH_AO22X9 port map( A => n2699, B => n2450, C => n2446, D => 
                           registers_13_1_port, Z => n1819);
   U2295 : HS65_LH_AO22X9 port map( A => n2701, B => n2450, C => n2447, D => 
                           registers_13_2_port, Z => n1820);
   U2296 : HS65_LH_AO22X9 port map( A => n2703, B => n2450, C => n2446, D => 
                           registers_13_3_port, Z => n1821);
   U2297 : HS65_LH_AO22X9 port map( A => n2705, B => n2450, C => n2447, D => 
                           registers_13_4_port, Z => n1822);
   U2298 : HS65_LH_AO22X9 port map( A => n2707, B => n2450, C => n2446, D => 
                           registers_13_5_port, Z => n1823);
   U2299 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2450, C => n2447, 
                           D => registers_13_6_port, Z => n1824);
   U2300 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2450, C => n2447,
                           D => registers_13_7_port, Z => n1825);
   U2301 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2450, C => n2447,
                           D => registers_13_8_port, Z => n1826);
   U2302 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2450, C => n2447,
                           D => registers_13_9_port, Z => n1827);
   U2303 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2450, C => n2447,
                           D => registers_13_10_port, Z => n1828);
   U2304 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2449, C => n2447,
                           D => registers_13_11_port, Z => n1829);
   U2305 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2449, C => n2447,
                           D => registers_13_12_port, Z => n1830);
   U2306 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2449, C => n2447,
                           D => registers_13_13_port, Z => n1831);
   U2307 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2449, C => n2447,
                           D => registers_13_14_port, Z => n1832);
   U2308 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2449, C => n2447,
                           D => registers_13_15_port, Z => n1833);
   U2309 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2449, C => n2447,
                           D => registers_13_16_port, Z => n1834);
   U2310 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2449, C => n2447,
                           D => registers_13_17_port, Z => n1835);
   U2311 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2449, C => n2447,
                           D => registers_13_18_port, Z => n1836);
   U2312 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2449, C => n2446,
                           D => registers_13_19_port, Z => n1837);
   U2313 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2449, C => n2446,
                           D => registers_13_20_port, Z => n1838);
   U2314 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2449, C => n2446,
                           D => registers_13_21_port, Z => n1839);
   U2315 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2449, C => n2446,
                           D => registers_13_22_port, Z => n1840);
   U2316 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2449, C => n2446,
                           D => registers_13_23_port, Z => n1841);
   U2317 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2449, C => n2446,
                           D => registers_13_24_port, Z => n1842);
   U2318 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2449, C => n2446,
                           D => registers_13_25_port, Z => n1843);
   U2319 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2449, C => n2446,
                           D => registers_13_26_port, Z => n1844);
   U2320 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2449, C => n2446,
                           D => registers_13_27_port, Z => n1845);
   U2321 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2449, C => n2446,
                           D => registers_13_28_port, Z => n1846);
   U2322 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2449, C => n2446,
                           D => registers_13_29_port, Z => n1847);
   U2323 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2449, C => n2446,
                           D => registers_13_30_port, Z => n1848);
   U2324 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2448, C => n2446,
                           D => registers_13_31_port, Z => n1849);
   U2325 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n322, C => n319, D 
                           => registers_25_0_port, Z => n2202);
   U2326 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n322, C => n318, D 
                           => registers_25_1_port, Z => n2203);
   U2327 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n322, C => n319, D 
                           => registers_25_2_port, Z => n2204);
   U2328 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n322, C => n318, D 
                           => registers_25_3_port, Z => n2205);
   U2329 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n322, C => n319, D 
                           => registers_25_4_port, Z => n2206);
   U2330 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n322, C => n318, D 
                           => registers_25_5_port, Z => n2207);
   U2331 : HS65_LH_AO22X9 port map( A => n2709, B => n322, C => n319, D => 
                           registers_25_6_port, Z => n2208);
   U2332 : HS65_LH_AO22X9 port map( A => n2711, B => n322, C => n319, D => 
                           registers_25_7_port, Z => n2209);
   U2333 : HS65_LH_AO22X9 port map( A => n2713, B => n322, C => n319, D => 
                           registers_25_8_port, Z => n2210);
   U2334 : HS65_LH_AO22X9 port map( A => n2715, B => n322, C => n319, D => 
                           registers_25_9_port, Z => n2211);
   U2335 : HS65_LH_AO22X9 port map( A => n2717, B => n322, C => n319, D => 
                           registers_25_10_port, Z => n2212);
   U2336 : HS65_LH_AO22X9 port map( A => n2719, B => n321, C => n319, D => 
                           registers_25_11_port, Z => n2213);
   U2337 : HS65_LH_AO22X9 port map( A => n2721, B => n321, C => n319, D => 
                           registers_25_12_port, Z => n2214);
   U2338 : HS65_LH_AO22X9 port map( A => n2723, B => n321, C => n319, D => 
                           registers_25_13_port, Z => n2215);
   U2339 : HS65_LH_AO22X9 port map( A => n2725, B => n321, C => n319, D => 
                           registers_25_14_port, Z => n2216);
   U2340 : HS65_LH_AO22X9 port map( A => n2727, B => n321, C => n319, D => 
                           registers_25_15_port, Z => n2217);
   U2341 : HS65_LH_AO22X9 port map( A => n2729, B => n321, C => n319, D => 
                           registers_25_16_port, Z => n2218);
   U2342 : HS65_LH_AO22X9 port map( A => n2731, B => n321, C => n319, D => 
                           registers_25_17_port, Z => n2219);
   U2343 : HS65_LH_AO22X9 port map( A => n2733, B => n321, C => n319, D => 
                           registers_25_18_port, Z => n2220);
   U2344 : HS65_LH_AO22X9 port map( A => n2735, B => n321, C => n318, D => 
                           registers_25_19_port, Z => n2221);
   U2345 : HS65_LH_AO22X9 port map( A => n2737, B => n321, C => n318, D => 
                           registers_25_20_port, Z => n2222);
   U2346 : HS65_LH_AO22X9 port map( A => n2739, B => n321, C => n318, D => 
                           registers_25_21_port, Z => n2223);
   U2347 : HS65_LH_AO22X9 port map( A => n2741, B => n321, C => n318, D => 
                           registers_25_22_port, Z => n2224);
   U2348 : HS65_LH_AO22X9 port map( A => n2743, B => n321, C => n318, D => 
                           registers_25_23_port, Z => n2225);
   U2349 : HS65_LH_AO22X9 port map( A => n2745, B => n321, C => n318, D => 
                           registers_25_24_port, Z => n2226);
   U2350 : HS65_LH_AO22X9 port map( A => n2747, B => n321, C => n318, D => 
                           registers_25_25_port, Z => n2227);
   U2351 : HS65_LH_AO22X9 port map( A => n2749, B => n321, C => n318, D => 
                           registers_25_26_port, Z => n2228);
   U2352 : HS65_LH_AO22X9 port map( A => n2751, B => n321, C => n318, D => 
                           registers_25_27_port, Z => n2229);
   U2353 : HS65_LH_AO22X9 port map( A => n2753, B => n321, C => n318, D => 
                           registers_25_28_port, Z => n2230);
   U2354 : HS65_LH_AO22X9 port map( A => n2755, B => n321, C => n318, D => 
                           registers_25_29_port, Z => n2231);
   U2355 : HS65_LH_AO22X9 port map( A => n2757, B => n321, C => n318, D => 
                           registers_25_30_port, Z => n2232);
   U2356 : HS65_LH_AO22X9 port map( A => n2759, B => n320, C => n318, D => 
                           registers_25_31_port, Z => n2233);
   U2357 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n292, C => n289, D 
                           => registers_31_0_port, Z => n2394);
   U2358 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n292, C => n288, D 
                           => registers_31_1_port, Z => n2395);
   U2359 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n292, C => n289, D 
                           => registers_31_2_port, Z => n2396);
   U2360 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n292, C => n288, D 
                           => registers_31_3_port, Z => n2397);
   U2361 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n292, C => n289, D 
                           => registers_31_4_port, Z => n2398);
   U2362 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n292, C => n288, D 
                           => registers_31_5_port, Z => n2399);
   U2363 : HS65_LH_AO22X9 port map( A => n2709, B => n292, C => n289, D => 
                           registers_31_6_port, Z => n2400);
   U2364 : HS65_LH_AO22X9 port map( A => n2711, B => n292, C => n289, D => 
                           registers_31_7_port, Z => n2401);
   U2365 : HS65_LH_AO22X9 port map( A => n2713, B => n292, C => n289, D => 
                           registers_31_8_port, Z => n2402);
   U2366 : HS65_LH_AO22X9 port map( A => n2715, B => n292, C => n289, D => 
                           registers_31_9_port, Z => n2403);
   U2367 : HS65_LH_AO22X9 port map( A => n2717, B => n292, C => n289, D => 
                           registers_31_10_port, Z => n2404);
   U2368 : HS65_LH_AO22X9 port map( A => n2719, B => n291, C => n289, D => 
                           registers_31_11_port, Z => n2405);
   U2369 : HS65_LH_AO22X9 port map( A => n2721, B => n291, C => n289, D => 
                           registers_31_12_port, Z => n2406);
   U2370 : HS65_LH_AO22X9 port map( A => n2723, B => n291, C => n289, D => 
                           registers_31_13_port, Z => n2407);
   U2371 : HS65_LH_AO22X9 port map( A => n2725, B => n291, C => n289, D => 
                           registers_31_14_port, Z => n2408);
   U2372 : HS65_LH_AO22X9 port map( A => n2727, B => n291, C => n289, D => 
                           registers_31_15_port, Z => n2409);
   U2373 : HS65_LH_AO22X9 port map( A => n2729, B => n291, C => n289, D => 
                           registers_31_16_port, Z => n2410);
   U2374 : HS65_LH_AO22X9 port map( A => n2731, B => n291, C => n289, D => 
                           registers_31_17_port, Z => n2411);
   U2375 : HS65_LH_AO22X9 port map( A => n2733, B => n291, C => n289, D => 
                           registers_31_18_port, Z => n2412);
   U2376 : HS65_LH_AO22X9 port map( A => n2735, B => n291, C => n288, D => 
                           registers_31_19_port, Z => n2413);
   U2377 : HS65_LH_AO22X9 port map( A => n2737, B => n291, C => n288, D => 
                           registers_31_20_port, Z => n2414);
   U2378 : HS65_LH_AO22X9 port map( A => n2739, B => n291, C => n288, D => 
                           registers_31_21_port, Z => n2415);
   U2379 : HS65_LH_AO22X9 port map( A => n2741, B => n291, C => n288, D => 
                           registers_31_22_port, Z => n2416);
   U2380 : HS65_LH_AO22X9 port map( A => n2743, B => n291, C => n288, D => 
                           registers_31_23_port, Z => n2417);
   U2381 : HS65_LH_AO22X9 port map( A => n2745, B => n291, C => n288, D => 
                           registers_31_24_port, Z => n2418);
   U2382 : HS65_LH_AO22X9 port map( A => n2747, B => n291, C => n288, D => 
                           registers_31_25_port, Z => n2419);
   U2383 : HS65_LH_AO22X9 port map( A => n2749, B => n291, C => n288, D => 
                           registers_31_26_port, Z => n2420);
   U2384 : HS65_LH_AO22X9 port map( A => n2751, B => n291, C => n288, D => 
                           registers_31_27_port, Z => n2421);
   U2385 : HS65_LH_AO22X9 port map( A => n2753, B => n291, C => n288, D => 
                           registers_31_28_port, Z => n2422);
   U2386 : HS65_LH_AO22X9 port map( A => n2755, B => n291, C => n288, D => 
                           registers_31_29_port, Z => n2423);
   U2387 : HS65_LH_AO22X9 port map( A => n2757, B => n291, C => n288, D => 
                           registers_31_30_port, Z => n2424);
   U2388 : HS65_LH_AO22X9 port map( A => n2759, B => n290, C => n288, D => 
                           registers_31_31_port, Z => n2425);
   U2389 : HS65_LH_AO22X9 port map( A => n2697, B => n2465, C => n2462, D => 
                           registers_10_0_port, Z => n1722);
   U2390 : HS65_LH_AO22X9 port map( A => n2699, B => n2465, C => n2461, D => 
                           registers_10_1_port, Z => n1723);
   U2391 : HS65_LH_AO22X9 port map( A => n2701, B => n2465, C => n2462, D => 
                           registers_10_2_port, Z => n1724);
   U2392 : HS65_LH_AO22X9 port map( A => n2703, B => n2465, C => n2461, D => 
                           registers_10_3_port, Z => n1725);
   U2393 : HS65_LH_AO22X9 port map( A => n2705, B => n2465, C => n2462, D => 
                           registers_10_4_port, Z => n1726);
   U2394 : HS65_LH_AO22X9 port map( A => n2707, B => n2465, C => n2461, D => 
                           registers_10_5_port, Z => n1727);
   U2395 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2465, C => n2462, 
                           D => registers_10_6_port, Z => n1728);
   U2396 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2465, C => n2462,
                           D => registers_10_7_port, Z => n1729);
   U2397 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2465, C => n2462,
                           D => registers_10_8_port, Z => n1730);
   U2398 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2465, C => n2462,
                           D => registers_10_9_port, Z => n1731);
   U2399 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2465, C => n2462,
                           D => registers_10_10_port, Z => n1732);
   U2400 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2464, C => n2462,
                           D => registers_10_11_port, Z => n1733);
   U2401 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2464, C => n2462,
                           D => registers_10_12_port, Z => n1734);
   U2402 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2464, C => n2462,
                           D => registers_10_13_port, Z => n1735);
   U2403 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2464, C => n2462,
                           D => registers_10_14_port, Z => n1736);
   U2404 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2464, C => n2462,
                           D => registers_10_15_port, Z => n1737);
   U2405 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2464, C => n2462,
                           D => registers_10_16_port, Z => n1738);
   U2406 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2464, C => n2462,
                           D => registers_10_17_port, Z => n1739);
   U2407 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2464, C => n2462,
                           D => registers_10_18_port, Z => n1740);
   U2408 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2464, C => n2461,
                           D => registers_10_19_port, Z => n1741);
   U2409 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2464, C => n2461,
                           D => registers_10_20_port, Z => n1742);
   U2410 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2464, C => n2461,
                           D => registers_10_21_port, Z => n1743);
   U2411 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2464, C => n2461,
                           D => registers_10_22_port, Z => n1744);
   U2412 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2464, C => n2461,
                           D => registers_10_23_port, Z => n1745);
   U2413 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2464, C => n2461,
                           D => registers_10_24_port, Z => n1746);
   U2414 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2464, C => n2461,
                           D => registers_10_25_port, Z => n1747);
   U2415 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2464, C => n2461,
                           D => registers_10_26_port, Z => n1748);
   U2416 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2464, C => n2461,
                           D => registers_10_27_port, Z => n1749);
   U2417 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2464, C => n2461,
                           D => registers_10_28_port, Z => n1750);
   U2418 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2464, C => n2461,
                           D => registers_10_29_port, Z => n1751);
   U2419 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2464, C => n2461,
                           D => registers_10_30_port, Z => n1752);
   U2420 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2463, C => n2461,
                           D => registers_10_31_port, Z => n1753);
   U2421 : HS65_LH_AO22X9 port map( A => n2697, B => n2455, C => n2452, D => 
                           registers_12_0_port, Z => n1786);
   U2422 : HS65_LH_AO22X9 port map( A => n2699, B => n2455, C => n2451, D => 
                           registers_12_1_port, Z => n1787);
   U2423 : HS65_LH_AO22X9 port map( A => n2701, B => n2455, C => n2452, D => 
                           registers_12_2_port, Z => n1788);
   U2424 : HS65_LH_AO22X9 port map( A => n2703, B => n2455, C => n2451, D => 
                           registers_12_3_port, Z => n1789);
   U2425 : HS65_LH_AO22X9 port map( A => n2705, B => n2455, C => n2452, D => 
                           registers_12_4_port, Z => n1790);
   U2426 : HS65_LH_AO22X9 port map( A => n2707, B => n2455, C => n2451, D => 
                           registers_12_5_port, Z => n1791);
   U2427 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2455, C => n2452, 
                           D => registers_12_6_port, Z => n1792);
   U2428 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2455, C => n2452,
                           D => registers_12_7_port, Z => n1793);
   U2429 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2455, C => n2452,
                           D => registers_12_8_port, Z => n1794);
   U2430 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2455, C => n2452,
                           D => registers_12_9_port, Z => n1795);
   U2431 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2455, C => n2452,
                           D => registers_12_10_port, Z => n1796);
   U2432 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2454, C => n2452,
                           D => registers_12_11_port, Z => n1797);
   U2433 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2454, C => n2452,
                           D => registers_12_12_port, Z => n1798);
   U2434 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2454, C => n2452,
                           D => registers_12_13_port, Z => n1799);
   U2435 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2454, C => n2452,
                           D => registers_12_14_port, Z => n1800);
   U2436 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2454, C => n2452,
                           D => registers_12_15_port, Z => n1801);
   U2437 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2454, C => n2452,
                           D => registers_12_16_port, Z => n1802);
   U2438 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2454, C => n2452,
                           D => registers_12_17_port, Z => n1803);
   U2439 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2454, C => n2452,
                           D => registers_12_18_port, Z => n1804);
   U2440 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2454, C => n2451,
                           D => registers_12_19_port, Z => n1805);
   U2441 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2454, C => n2451,
                           D => registers_12_20_port, Z => n1806);
   U2442 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2454, C => n2451,
                           D => registers_12_21_port, Z => n1807);
   U2443 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2454, C => n2451,
                           D => registers_12_22_port, Z => n1808);
   U2444 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2454, C => n2451,
                           D => registers_12_23_port, Z => n1809);
   U2445 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2454, C => n2451,
                           D => registers_12_24_port, Z => n1810);
   U2446 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2454, C => n2451,
                           D => registers_12_25_port, Z => n1811);
   U2447 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2454, C => n2451,
                           D => registers_12_26_port, Z => n1812);
   U2448 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2454, C => n2451,
                           D => registers_12_27_port, Z => n1813);
   U2449 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2454, C => n2451,
                           D => registers_12_28_port, Z => n1814);
   U2450 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2454, C => n2451,
                           D => registers_12_29_port, Z => n1815);
   U2451 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2454, C => n2451,
                           D => registers_12_30_port, Z => n1816);
   U2452 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2453, C => n2451,
                           D => registers_12_31_port, Z => n1817);
   U2453 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n326, C => n323, D 
                           => registers_24_0_port, Z => n2170);
   U2454 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n326, C => n323, D 
                           => registers_24_1_port, Z => n2171);
   U2455 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n326, C => n323, D 
                           => registers_24_2_port, Z => n2172);
   U2456 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n326, C => n323, D 
                           => registers_24_3_port, Z => n2173);
   U2457 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n326, C => n323, D 
                           => registers_24_4_port, Z => n2174);
   U2458 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n326, C => n323, D 
                           => registers_24_5_port, Z => n2175);
   U2459 : HS65_LH_AO22X9 port map( A => n2709, B => n326, C => n323, D => 
                           registers_24_6_port, Z => n2176);
   U2460 : HS65_LH_AO22X9 port map( A => n2711, B => n326, C => n323, D => 
                           registers_24_7_port, Z => n2177);
   U2461 : HS65_LH_AO22X9 port map( A => n2713, B => n326, C => n323, D => 
                           registers_24_8_port, Z => n2178);
   U2462 : HS65_LH_AO22X9 port map( A => n2715, B => n326, C => n323, D => 
                           registers_24_9_port, Z => n2179);
   U2463 : HS65_LH_AO22X9 port map( A => n2717, B => n326, C => n323, D => 
                           registers_24_10_port, Z => n2180);
   U2464 : HS65_LH_AO22X9 port map( A => n2719, B => n325, C => n323, D => 
                           registers_24_11_port, Z => n2181);
   U2465 : HS65_LH_AO22X9 port map( A => n2721, B => n325, C => n323, D => 
                           registers_24_12_port, Z => n2182);
   U2466 : HS65_LH_AO22X9 port map( A => n2723, B => n325, C => n323, D => 
                           registers_24_13_port, Z => n2183);
   U2467 : HS65_LH_AO22X9 port map( A => n2725, B => n325, C => n323, D => 
                           registers_24_14_port, Z => n2184);
   U2468 : HS65_LH_AO22X9 port map( A => n2727, B => n325, C => n323, D => 
                           registers_24_15_port, Z => n2185);
   U2469 : HS65_LH_AO22X9 port map( A => n2729, B => n325, C => n323, D => 
                           registers_24_16_port, Z => n2186);
   U2470 : HS65_LH_AO22X9 port map( A => n2731, B => n325, C => n323, D => 
                           registers_24_17_port, Z => n2187);
   U2471 : HS65_LH_AO22X9 port map( A => n2733, B => n325, C => n323, D => 
                           registers_24_18_port, Z => n2188);
   U2472 : HS65_LH_AO22X9 port map( A => n2735, B => n325, C => n323, D => 
                           registers_24_19_port, Z => n2189);
   U2473 : HS65_LH_AO22X9 port map( A => n2737, B => n325, C => n1425, D => 
                           registers_24_20_port, Z => n2190);
   U2474 : HS65_LH_AO22X9 port map( A => n2739, B => n325, C => n1425, D => 
                           registers_24_21_port, Z => n2191);
   U2475 : HS65_LH_AO22X9 port map( A => n2741, B => n325, C => n1425, D => 
                           registers_24_22_port, Z => n2192);
   U2476 : HS65_LH_AO22X9 port map( A => n2743, B => n325, C => n1425, D => 
                           registers_24_23_port, Z => n2193);
   U2477 : HS65_LH_AO22X9 port map( A => n2745, B => n325, C => n1425, D => 
                           registers_24_24_port, Z => n2194);
   U2478 : HS65_LH_AO22X9 port map( A => n2747, B => n325, C => n1425, D => 
                           registers_24_25_port, Z => n2195);
   U2479 : HS65_LH_AO22X9 port map( A => n2749, B => n325, C => n1425, D => 
                           registers_24_26_port, Z => n2196);
   U2480 : HS65_LH_AO22X9 port map( A => n2751, B => n325, C => n1425, D => 
                           registers_24_27_port, Z => n2197);
   U2481 : HS65_LH_AO22X9 port map( A => n2753, B => n325, C => n1425, D => 
                           registers_24_28_port, Z => n2198);
   U2482 : HS65_LH_AO22X9 port map( A => n2755, B => n325, C => n1425, D => 
                           registers_24_29_port, Z => n2199);
   U2483 : HS65_LH_AO22X9 port map( A => n2757, B => n325, C => n1425, D => 
                           registers_24_30_port, Z => n2200);
   U2484 : HS65_LH_AO22X9 port map( A => n2759, B => n324, C => n1425, D => 
                           registers_24_31_port, Z => n2201);
   U2485 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n297, C => n294, D 
                           => registers_30_0_port, Z => n2362);
   U2486 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n297, C => n293, D 
                           => registers_30_1_port, Z => n2363);
   U2487 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n297, C => n294, D 
                           => registers_30_2_port, Z => n2364);
   U2488 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n297, C => n293, D 
                           => registers_30_3_port, Z => n2365);
   U2489 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n297, C => n294, D 
                           => registers_30_4_port, Z => n2366);
   U2490 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n297, C => n293, D 
                           => registers_30_5_port, Z => n2367);
   U2491 : HS65_LH_AO22X9 port map( A => n2709, B => n297, C => n294, D => 
                           registers_30_6_port, Z => n2368);
   U2492 : HS65_LH_AO22X9 port map( A => n2711, B => n297, C => n294, D => 
                           registers_30_7_port, Z => n2369);
   U2493 : HS65_LH_AO22X9 port map( A => n2713, B => n297, C => n294, D => 
                           registers_30_8_port, Z => n2370);
   U2494 : HS65_LH_AO22X9 port map( A => n2715, B => n297, C => n294, D => 
                           registers_30_9_port, Z => n2371);
   U2495 : HS65_LH_AO22X9 port map( A => n2717, B => n297, C => n294, D => 
                           registers_30_10_port, Z => n2372);
   U2496 : HS65_LH_AO22X9 port map( A => n2719, B => n296, C => n294, D => 
                           registers_30_11_port, Z => n2373);
   U2497 : HS65_LH_AO22X9 port map( A => n2721, B => n296, C => n294, D => 
                           registers_30_12_port, Z => n2374);
   U2498 : HS65_LH_AO22X9 port map( A => n2723, B => n296, C => n294, D => 
                           registers_30_13_port, Z => n2375);
   U2499 : HS65_LH_AO22X9 port map( A => n2725, B => n296, C => n294, D => 
                           registers_30_14_port, Z => n2376);
   U2500 : HS65_LH_AO22X9 port map( A => n2727, B => n296, C => n294, D => 
                           registers_30_15_port, Z => n2377);
   U2501 : HS65_LH_AO22X9 port map( A => n2729, B => n296, C => n294, D => 
                           registers_30_16_port, Z => n2378);
   U2502 : HS65_LH_AO22X9 port map( A => n2731, B => n296, C => n294, D => 
                           registers_30_17_port, Z => n2379);
   U2503 : HS65_LH_AO22X9 port map( A => n2733, B => n296, C => n294, D => 
                           registers_30_18_port, Z => n2380);
   U2504 : HS65_LH_AO22X9 port map( A => n2735, B => n296, C => n293, D => 
                           registers_30_19_port, Z => n2381);
   U2505 : HS65_LH_AO22X9 port map( A => n2737, B => n296, C => n293, D => 
                           registers_30_20_port, Z => n2382);
   U2506 : HS65_LH_AO22X9 port map( A => n2739, B => n296, C => n293, D => 
                           registers_30_21_port, Z => n2383);
   U2507 : HS65_LH_AO22X9 port map( A => n2741, B => n296, C => n293, D => 
                           registers_30_22_port, Z => n2384);
   U2508 : HS65_LH_AO22X9 port map( A => n2743, B => n296, C => n293, D => 
                           registers_30_23_port, Z => n2385);
   U2509 : HS65_LH_AO22X9 port map( A => n2745, B => n296, C => n293, D => 
                           registers_30_24_port, Z => n2386);
   U2510 : HS65_LH_AO22X9 port map( A => n2747, B => n296, C => n293, D => 
                           registers_30_25_port, Z => n2387);
   U2511 : HS65_LH_AO22X9 port map( A => n2749, B => n296, C => n293, D => 
                           registers_30_26_port, Z => n2388);
   U2512 : HS65_LH_AO22X9 port map( A => n2751, B => n296, C => n293, D => 
                           registers_30_27_port, Z => n2389);
   U2513 : HS65_LH_AO22X9 port map( A => n2753, B => n296, C => n293, D => 
                           registers_30_28_port, Z => n2390);
   U2514 : HS65_LH_AO22X9 port map( A => n2755, B => n296, C => n293, D => 
                           registers_30_29_port, Z => n2391);
   U2515 : HS65_LH_AO22X9 port map( A => n2757, B => n296, C => n293, D => 
                           registers_30_30_port, Z => n2392);
   U2516 : HS65_LH_AO22X9 port map( A => n2759, B => n295, C => n293, D => 
                           registers_30_31_port, Z => n2393);
   U2517 : HS65_LH_AO22X9 port map( A => n2697, B => n2480, C => n2477, D => 
                           registers_7_0_port, Z => n1626);
   U2518 : HS65_LH_AO22X9 port map( A => n2699, B => n2480, C => n2476, D => 
                           registers_7_1_port, Z => n1627);
   U2519 : HS65_LH_AO22X9 port map( A => n2701, B => n2480, C => n2477, D => 
                           registers_7_2_port, Z => n1628);
   U2520 : HS65_LH_AO22X9 port map( A => n2703, B => n2480, C => n2476, D => 
                           registers_7_3_port, Z => n1629);
   U2521 : HS65_LH_AO22X9 port map( A => n2705, B => n2480, C => n2477, D => 
                           registers_7_4_port, Z => n1630);
   U2522 : HS65_LH_AO22X9 port map( A => n2707, B => n2480, C => n2476, D => 
                           registers_7_5_port, Z => n1631);
   U2523 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2480, C => n2477, 
                           D => registers_7_6_port, Z => n1632);
   U2524 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2480, C => n2477,
                           D => registers_7_7_port, Z => n1633);
   U2525 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2480, C => n2477,
                           D => registers_7_8_port, Z => n1634);
   U2526 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2480, C => n2477,
                           D => registers_7_9_port, Z => n1635);
   U2527 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2480, C => n2477,
                           D => registers_7_10_port, Z => n1636);
   U2528 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2479, C => n2477,
                           D => registers_7_11_port, Z => n1637);
   U2529 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2479, C => n2477,
                           D => registers_7_12_port, Z => n1638);
   U2530 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2479, C => n2477,
                           D => registers_7_13_port, Z => n1639);
   U2531 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2479, C => n2477,
                           D => registers_7_14_port, Z => n1640);
   U2532 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2479, C => n2477,
                           D => registers_7_15_port, Z => n1641);
   U2533 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2479, C => n2477,
                           D => registers_7_16_port, Z => n1642);
   U2534 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2479, C => n2477,
                           D => registers_7_17_port, Z => n1643);
   U2535 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2479, C => n2477,
                           D => registers_7_18_port, Z => n1644);
   U2536 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2479, C => n2476,
                           D => registers_7_19_port, Z => n1645);
   U2537 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2479, C => n2476,
                           D => registers_7_20_port, Z => n1646);
   U2538 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2479, C => n2476,
                           D => registers_7_21_port, Z => n1647);
   U2539 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2479, C => n2476,
                           D => registers_7_22_port, Z => n1648);
   U2540 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2479, C => n2476,
                           D => registers_7_23_port, Z => n1649);
   U2541 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2479, C => n2476,
                           D => registers_7_24_port, Z => n1650);
   U2542 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2479, C => n2476,
                           D => registers_7_25_port, Z => n1651);
   U2543 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2479, C => n2476,
                           D => registers_7_26_port, Z => n1652);
   U2544 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2479, C => n2476,
                           D => registers_7_27_port, Z => n1653);
   U2545 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2479, C => n2476,
                           D => registers_7_28_port, Z => n1654);
   U2546 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2479, C => n2476,
                           D => registers_7_29_port, Z => n1655);
   U2547 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2479, C => n2476,
                           D => registers_7_30_port, Z => n1656);
   U2548 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2478, C => n2476,
                           D => registers_7_31_port, Z => n1657);
   U2549 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n1422, C => n1419, 
                           D => registers_19_0_port, Z => n2010);
   U2550 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n1422, C => n1418, 
                           D => registers_19_1_port, Z => n2011);
   U2551 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n1422, C => n1419, 
                           D => registers_19_2_port, Z => n2012);
   U2552 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n1422, C => n1418, 
                           D => registers_19_3_port, Z => n2013);
   U2553 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n1422, C => n1419, 
                           D => registers_19_4_port, Z => n2014);
   U2554 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n1422, C => n1418, 
                           D => registers_19_5_port, Z => n2015);
   U2555 : HS65_LH_AO22X9 port map( A => n2709, B => n1422, C => n1419, D => 
                           registers_19_6_port, Z => n2016);
   U2556 : HS65_LH_AO22X9 port map( A => n2711, B => n1422, C => n1419, D => 
                           registers_19_7_port, Z => n2017);
   U2557 : HS65_LH_AO22X9 port map( A => n2713, B => n1422, C => n1419, D => 
                           registers_19_8_port, Z => n2018);
   U2558 : HS65_LH_AO22X9 port map( A => n2715, B => n1422, C => n1419, D => 
                           registers_19_9_port, Z => n2019);
   U2559 : HS65_LH_AO22X9 port map( A => n2717, B => n1422, C => n1419, D => 
                           registers_19_10_port, Z => n2020);
   U2560 : HS65_LH_AO22X9 port map( A => n2719, B => n1421, C => n1419, D => 
                           registers_19_11_port, Z => n2021);
   U2561 : HS65_LH_AO22X9 port map( A => n2721, B => n1421, C => n1419, D => 
                           registers_19_12_port, Z => n2022);
   U2562 : HS65_LH_AO22X9 port map( A => n2723, B => n1421, C => n1419, D => 
                           registers_19_13_port, Z => n2023);
   U2563 : HS65_LH_AO22X9 port map( A => n2725, B => n1421, C => n1419, D => 
                           registers_19_14_port, Z => n2024);
   U2564 : HS65_LH_AO22X9 port map( A => n2727, B => n1421, C => n1419, D => 
                           registers_19_15_port, Z => n2025);
   U2565 : HS65_LH_AO22X9 port map( A => n2729, B => n1421, C => n1419, D => 
                           registers_19_16_port, Z => n2026);
   U2566 : HS65_LH_AO22X9 port map( A => n2731, B => n1421, C => n1419, D => 
                           registers_19_17_port, Z => n2027);
   U2567 : HS65_LH_AO22X9 port map( A => n2733, B => n1421, C => n1419, D => 
                           registers_19_18_port, Z => n2028);
   U2568 : HS65_LH_AO22X9 port map( A => n2735, B => n1421, C => n1418, D => 
                           registers_19_19_port, Z => n2029);
   U2569 : HS65_LH_AO22X9 port map( A => n2737, B => n1421, C => n1418, D => 
                           registers_19_20_port, Z => n2030);
   U2570 : HS65_LH_AO22X9 port map( A => n2739, B => n1421, C => n1418, D => 
                           registers_19_21_port, Z => n2031);
   U2571 : HS65_LH_AO22X9 port map( A => n2741, B => n1421, C => n1418, D => 
                           registers_19_22_port, Z => n2032);
   U2572 : HS65_LH_AO22X9 port map( A => n2743, B => n1421, C => n1418, D => 
                           registers_19_23_port, Z => n2033);
   U2573 : HS65_LH_AO22X9 port map( A => n2745, B => n1421, C => n1418, D => 
                           registers_19_24_port, Z => n2034);
   U2574 : HS65_LH_AO22X9 port map( A => n2747, B => n1421, C => n1418, D => 
                           registers_19_25_port, Z => n2035);
   U2575 : HS65_LH_AO22X9 port map( A => n2749, B => n1421, C => n1418, D => 
                           registers_19_26_port, Z => n2036);
   U2576 : HS65_LH_AO22X9 port map( A => n2751, B => n1421, C => n1418, D => 
                           registers_19_27_port, Z => n2037);
   U2577 : HS65_LH_AO22X9 port map( A => n2753, B => n1421, C => n1418, D => 
                           registers_19_28_port, Z => n2038);
   U2578 : HS65_LH_AO22X9 port map( A => n2755, B => n1421, C => n1418, D => 
                           registers_19_29_port, Z => n2039);
   U2579 : HS65_LH_AO22X9 port map( A => n2757, B => n1421, C => n1418, D => 
                           registers_19_30_port, Z => n2040);
   U2580 : HS65_LH_AO22X9 port map( A => n2759, B => n1420, C => n1418, D => 
                           registers_19_31_port, Z => n2041);
   U2581 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n332, C => n329, D 
                           => registers_23_0_port, Z => n2138);
   U2582 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n332, C => n328, D 
                           => registers_23_1_port, Z => n2139);
   U2583 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n332, C => n329, D 
                           => registers_23_2_port, Z => n2140);
   U2584 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n332, C => n328, D 
                           => registers_23_3_port, Z => n2141);
   U2585 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n332, C => n329, D 
                           => registers_23_4_port, Z => n2142);
   U2586 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n332, C => n328, D 
                           => registers_23_5_port, Z => n2143);
   U2587 : HS65_LH_AO22X9 port map( A => n2709, B => n332, C => n329, D => 
                           registers_23_6_port, Z => n2144);
   U2588 : HS65_LH_AO22X9 port map( A => n2711, B => n332, C => n329, D => 
                           registers_23_7_port, Z => n2145);
   U2589 : HS65_LH_AO22X9 port map( A => n2713, B => n332, C => n329, D => 
                           registers_23_8_port, Z => n2146);
   U2590 : HS65_LH_AO22X9 port map( A => n2715, B => n332, C => n329, D => 
                           registers_23_9_port, Z => n2147);
   U2591 : HS65_LH_AO22X9 port map( A => n2717, B => n332, C => n329, D => 
                           registers_23_10_port, Z => n2148);
   U2592 : HS65_LH_AO22X9 port map( A => n2719, B => n331, C => n329, D => 
                           registers_23_11_port, Z => n2149);
   U2593 : HS65_LH_AO22X9 port map( A => n2721, B => n331, C => n329, D => 
                           registers_23_12_port, Z => n2150);
   U2594 : HS65_LH_AO22X9 port map( A => n2723, B => n331, C => n329, D => 
                           registers_23_13_port, Z => n2151);
   U2595 : HS65_LH_AO22X9 port map( A => n2725, B => n331, C => n329, D => 
                           registers_23_14_port, Z => n2152);
   U2596 : HS65_LH_AO22X9 port map( A => n2727, B => n331, C => n329, D => 
                           registers_23_15_port, Z => n2153);
   U2597 : HS65_LH_AO22X9 port map( A => n2729, B => n331, C => n329, D => 
                           registers_23_16_port, Z => n2154);
   U2598 : HS65_LH_AO22X9 port map( A => n2731, B => n331, C => n329, D => 
                           registers_23_17_port, Z => n2155);
   U2599 : HS65_LH_AO22X9 port map( A => n2733, B => n331, C => n329, D => 
                           registers_23_18_port, Z => n2156);
   U2600 : HS65_LH_AO22X9 port map( A => n2735, B => n331, C => n328, D => 
                           registers_23_19_port, Z => n2157);
   U2601 : HS65_LH_AO22X9 port map( A => n2737, B => n331, C => n328, D => 
                           registers_23_20_port, Z => n2158);
   U2602 : HS65_LH_AO22X9 port map( A => n2739, B => n331, C => n328, D => 
                           registers_23_21_port, Z => n2159);
   U2603 : HS65_LH_AO22X9 port map( A => n2741, B => n331, C => n328, D => 
                           registers_23_22_port, Z => n2160);
   U2604 : HS65_LH_AO22X9 port map( A => n2743, B => n331, C => n328, D => 
                           registers_23_23_port, Z => n2161);
   U2605 : HS65_LH_AO22X9 port map( A => n2745, B => n331, C => n328, D => 
                           registers_23_24_port, Z => n2162);
   U2606 : HS65_LH_AO22X9 port map( A => n2747, B => n331, C => n328, D => 
                           registers_23_25_port, Z => n2163);
   U2607 : HS65_LH_AO22X9 port map( A => n2749, B => n331, C => n328, D => 
                           registers_23_26_port, Z => n2164);
   U2608 : HS65_LH_AO22X9 port map( A => n2751, B => n331, C => n328, D => 
                           registers_23_27_port, Z => n2165);
   U2609 : HS65_LH_AO22X9 port map( A => n2753, B => n331, C => n328, D => 
                           registers_23_28_port, Z => n2166);
   U2610 : HS65_LH_AO22X9 port map( A => n2755, B => n331, C => n328, D => 
                           registers_23_29_port, Z => n2167);
   U2611 : HS65_LH_AO22X9 port map( A => n2757, B => n331, C => n328, D => 
                           registers_23_30_port, Z => n2168);
   U2612 : HS65_LH_AO22X9 port map( A => n2759, B => n330, C => n328, D => 
                           registers_23_31_port, Z => n2169);
   U2613 : HS65_LH_AO22X9 port map( A => n2697, B => n2490, C => n2487, D => 
                           registers_5_0_port, Z => n1562);
   U2614 : HS65_LH_AO22X9 port map( A => n2699, B => n2490, C => n2486, D => 
                           registers_5_1_port, Z => n1563);
   U2615 : HS65_LH_AO22X9 port map( A => n2701, B => n2490, C => n2487, D => 
                           registers_5_2_port, Z => n1564);
   U2616 : HS65_LH_AO22X9 port map( A => n2703, B => n2490, C => n2486, D => 
                           registers_5_3_port, Z => n1565);
   U2617 : HS65_LH_AO22X9 port map( A => n2705, B => n2490, C => n2487, D => 
                           registers_5_4_port, Z => n1566);
   U2618 : HS65_LH_AO22X9 port map( A => n2707, B => n2490, C => n2486, D => 
                           registers_5_5_port, Z => n1567);
   U2619 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2490, C => n2487, 
                           D => registers_5_6_port, Z => n1568);
   U2620 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2490, C => n2487,
                           D => registers_5_7_port, Z => n1569);
   U2621 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2490, C => n2487,
                           D => registers_5_8_port, Z => n1570);
   U2622 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2490, C => n2487,
                           D => registers_5_9_port, Z => n1571);
   U2623 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2490, C => n2487,
                           D => registers_5_10_port, Z => n1572);
   U2624 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2489, C => n2487,
                           D => registers_5_11_port, Z => n1573);
   U2625 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2489, C => n2487,
                           D => registers_5_12_port, Z => n1574);
   U2626 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2489, C => n2487,
                           D => registers_5_13_port, Z => n1575);
   U2627 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2489, C => n2487,
                           D => registers_5_14_port, Z => n1576);
   U2628 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2489, C => n2487,
                           D => registers_5_15_port, Z => n1577);
   U2629 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2489, C => n2487,
                           D => registers_5_16_port, Z => n1578);
   U2630 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2489, C => n2487,
                           D => registers_5_17_port, Z => n1579);
   U2631 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2489, C => n2487,
                           D => registers_5_18_port, Z => n1580);
   U2632 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2489, C => n2486,
                           D => registers_5_19_port, Z => n1581);
   U2633 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2489, C => n2486,
                           D => registers_5_20_port, Z => n1582);
   U2634 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2489, C => n2486,
                           D => registers_5_21_port, Z => n1583);
   U2635 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2489, C => n2486,
                           D => registers_5_22_port, Z => n1584);
   U2636 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2489, C => n2486,
                           D => registers_5_23_port, Z => n1585);
   U2637 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2489, C => n2486,
                           D => registers_5_24_port, Z => n1586);
   U2638 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2489, C => n2486,
                           D => registers_5_25_port, Z => n1587);
   U2639 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2489, C => n2486,
                           D => registers_5_26_port, Z => n1588);
   U2640 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2489, C => n2486,
                           D => registers_5_27_port, Z => n1589);
   U2641 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2489, C => n2486,
                           D => registers_5_28_port, Z => n1590);
   U2642 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2489, C => n2486,
                           D => registers_5_29_port, Z => n1591);
   U2643 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2489, C => n2486,
                           D => registers_5_30_port, Z => n1592);
   U2644 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2488, C => n2486,
                           D => registers_5_31_port, Z => n1593);
   U2645 : HS65_LH_AO22X9 port map( A => n2697, B => n2485, C => n2482, D => 
                           registers_6_0_port, Z => n1594);
   U2646 : HS65_LH_AO22X9 port map( A => n2699, B => n2485, C => n2481, D => 
                           registers_6_1_port, Z => n1595);
   U2647 : HS65_LH_AO22X9 port map( A => n2701, B => n2485, C => n2482, D => 
                           registers_6_2_port, Z => n1596);
   U2648 : HS65_LH_AO22X9 port map( A => n2703, B => n2485, C => n2481, D => 
                           registers_6_3_port, Z => n1597);
   U2649 : HS65_LH_AO22X9 port map( A => n2705, B => n2485, C => n2482, D => 
                           registers_6_4_port, Z => n1598);
   U2650 : HS65_LH_AO22X9 port map( A => n2707, B => n2485, C => n2481, D => 
                           registers_6_5_port, Z => n1599);
   U2651 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2485, C => n2482, 
                           D => registers_6_6_port, Z => n1600);
   U2652 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2485, C => n2482,
                           D => registers_6_7_port, Z => n1601);
   U2653 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2485, C => n2482,
                           D => registers_6_8_port, Z => n1602);
   U2654 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2485, C => n2482,
                           D => registers_6_9_port, Z => n1603);
   U2655 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2485, C => n2482,
                           D => registers_6_10_port, Z => n1604);
   U2656 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2484, C => n2482,
                           D => registers_6_11_port, Z => n1605);
   U2657 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2484, C => n2482,
                           D => registers_6_12_port, Z => n1606);
   U2658 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2484, C => n2482,
                           D => registers_6_13_port, Z => n1607);
   U2659 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2484, C => n2482,
                           D => registers_6_14_port, Z => n1608);
   U2660 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2484, C => n2482,
                           D => registers_6_15_port, Z => n1609);
   U2661 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2484, C => n2482,
                           D => registers_6_16_port, Z => n1610);
   U2662 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2484, C => n2482,
                           D => registers_6_17_port, Z => n1611);
   U2663 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2484, C => n2482,
                           D => registers_6_18_port, Z => n1612);
   U2664 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2484, C => n2481,
                           D => registers_6_19_port, Z => n1613);
   U2665 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2484, C => n2481,
                           D => registers_6_20_port, Z => n1614);
   U2666 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2484, C => n2481,
                           D => registers_6_21_port, Z => n1615);
   U2667 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2484, C => n2481,
                           D => registers_6_22_port, Z => n1616);
   U2668 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2484, C => n2481,
                           D => registers_6_23_port, Z => n1617);
   U2669 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2484, C => n2481,
                           D => registers_6_24_port, Z => n1618);
   U2670 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2484, C => n2481,
                           D => registers_6_25_port, Z => n1619);
   U2671 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2484, C => n2481,
                           D => registers_6_26_port, Z => n1620);
   U2672 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2484, C => n2481,
                           D => registers_6_27_port, Z => n1621);
   U2673 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2484, C => n2481,
                           D => registers_6_28_port, Z => n1622);
   U2674 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2484, C => n2481,
                           D => registers_6_29_port, Z => n1623);
   U2675 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2484, C => n2481,
                           D => registers_6_30_port, Z => n1624);
   U2676 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2483, C => n2481,
                           D => registers_6_31_port, Z => n1625);
   U2677 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n2430, C => n2427, 
                           D => registers_17_0_port, Z => n1946);
   U2678 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n2430, C => n2426, 
                           D => registers_17_1_port, Z => n1947);
   U2679 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n2430, C => n2427, 
                           D => registers_17_2_port, Z => n1948);
   U2680 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n2430, C => n2426, 
                           D => registers_17_3_port, Z => n1949);
   U2681 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n2430, C => n2427, 
                           D => registers_17_4_port, Z => n1950);
   U2682 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n2430, C => n2426, 
                           D => registers_17_5_port, Z => n1951);
   U2683 : HS65_LH_AO22X9 port map( A => n2709, B => n2430, C => n2427, D => 
                           registers_17_6_port, Z => n1952);
   U2684 : HS65_LH_AO22X9 port map( A => n2711, B => n2430, C => n2427, D => 
                           registers_17_7_port, Z => n1953);
   U2685 : HS65_LH_AO22X9 port map( A => n2713, B => n2430, C => n2427, D => 
                           registers_17_8_port, Z => n1954);
   U2686 : HS65_LH_AO22X9 port map( A => n2715, B => n2430, C => n2427, D => 
                           registers_17_9_port, Z => n1955);
   U2687 : HS65_LH_AO22X9 port map( A => n2717, B => n2430, C => n2427, D => 
                           registers_17_10_port, Z => n1956);
   U2688 : HS65_LH_AO22X9 port map( A => n2719, B => n2429, C => n2427, D => 
                           registers_17_11_port, Z => n1957);
   U2689 : HS65_LH_AO22X9 port map( A => n2721, B => n2429, C => n2427, D => 
                           registers_17_12_port, Z => n1958);
   U2690 : HS65_LH_AO22X9 port map( A => n2723, B => n2429, C => n2427, D => 
                           registers_17_13_port, Z => n1959);
   U2691 : HS65_LH_AO22X9 port map( A => n2725, B => n2429, C => n2427, D => 
                           registers_17_14_port, Z => n1960);
   U2692 : HS65_LH_AO22X9 port map( A => n2727, B => n2429, C => n2427, D => 
                           registers_17_15_port, Z => n1961);
   U2693 : HS65_LH_AO22X9 port map( A => n2729, B => n2429, C => n2427, D => 
                           registers_17_16_port, Z => n1962);
   U2694 : HS65_LH_AO22X9 port map( A => n2731, B => n2429, C => n2427, D => 
                           registers_17_17_port, Z => n1963);
   U2695 : HS65_LH_AO22X9 port map( A => n2733, B => n2429, C => n2427, D => 
                           registers_17_18_port, Z => n1964);
   U2696 : HS65_LH_AO22X9 port map( A => n2735, B => n2429, C => n2426, D => 
                           registers_17_19_port, Z => n1965);
   U2697 : HS65_LH_AO22X9 port map( A => n2737, B => n2429, C => n2426, D => 
                           registers_17_20_port, Z => n1966);
   U2698 : HS65_LH_AO22X9 port map( A => n2739, B => n2429, C => n2426, D => 
                           registers_17_21_port, Z => n1967);
   U2699 : HS65_LH_AO22X9 port map( A => n2741, B => n2429, C => n2426, D => 
                           registers_17_22_port, Z => n1968);
   U2700 : HS65_LH_AO22X9 port map( A => n2743, B => n2429, C => n2426, D => 
                           registers_17_23_port, Z => n1969);
   U2701 : HS65_LH_AO22X9 port map( A => n2745, B => n2429, C => n2426, D => 
                           registers_17_24_port, Z => n1970);
   U2702 : HS65_LH_AO22X9 port map( A => n2747, B => n2429, C => n2426, D => 
                           registers_17_25_port, Z => n1971);
   U2703 : HS65_LH_AO22X9 port map( A => n2749, B => n2429, C => n2426, D => 
                           registers_17_26_port, Z => n1972);
   U2704 : HS65_LH_AO22X9 port map( A => n2751, B => n2429, C => n2426, D => 
                           registers_17_27_port, Z => n1973);
   U2705 : HS65_LH_AO22X9 port map( A => n2753, B => n2429, C => n2426, D => 
                           registers_17_28_port, Z => n1974);
   U2706 : HS65_LH_AO22X9 port map( A => n2755, B => n2429, C => n2426, D => 
                           registers_17_29_port, Z => n1975);
   U2707 : HS65_LH_AO22X9 port map( A => n2757, B => n2429, C => n2426, D => 
                           registers_17_30_port, Z => n1976);
   U2708 : HS65_LH_AO22X9 port map( A => n2759, B => n2428, C => n2426, D => 
                           registers_17_31_port, Z => n1977);
   U2709 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n1433, C => n1424, 
                           D => registers_18_0_port, Z => n1978);
   U2710 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n1433, C => n1423, 
                           D => registers_18_1_port, Z => n1979);
   U2711 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n1433, C => n1424, 
                           D => registers_18_2_port, Z => n1980);
   U2712 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n1433, C => n1423, 
                           D => registers_18_3_port, Z => n1981);
   U2713 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n1433, C => n1424, 
                           D => registers_18_4_port, Z => n1982);
   U2714 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n1433, C => n1423, 
                           D => registers_18_5_port, Z => n1983);
   U2715 : HS65_LH_AO22X9 port map( A => n2709, B => n1433, C => n1424, D => 
                           registers_18_6_port, Z => n1984);
   U2716 : HS65_LH_AO22X9 port map( A => n2711, B => n1433, C => n1424, D => 
                           registers_18_7_port, Z => n1985);
   U2717 : HS65_LH_AO22X9 port map( A => n2713, B => n1433, C => n1424, D => 
                           registers_18_8_port, Z => n1986);
   U2718 : HS65_LH_AO22X9 port map( A => n2715, B => n1433, C => n1424, D => 
                           registers_18_9_port, Z => n1987);
   U2719 : HS65_LH_AO22X9 port map( A => n2717, B => n1433, C => n1424, D => 
                           registers_18_10_port, Z => n1988);
   U2720 : HS65_LH_AO22X9 port map( A => n2719, B => n1432, C => n1424, D => 
                           registers_18_11_port, Z => n1989);
   U2721 : HS65_LH_AO22X9 port map( A => n2721, B => n1432, C => n1424, D => 
                           registers_18_12_port, Z => n1990);
   U2722 : HS65_LH_AO22X9 port map( A => n2723, B => n1432, C => n1424, D => 
                           registers_18_13_port, Z => n1991);
   U2723 : HS65_LH_AO22X9 port map( A => n2725, B => n1432, C => n1424, D => 
                           registers_18_14_port, Z => n1992);
   U2724 : HS65_LH_AO22X9 port map( A => n2727, B => n1432, C => n1424, D => 
                           registers_18_15_port, Z => n1993);
   U2725 : HS65_LH_AO22X9 port map( A => n2729, B => n1432, C => n1424, D => 
                           registers_18_16_port, Z => n1994);
   U2726 : HS65_LH_AO22X9 port map( A => n2731, B => n1432, C => n1424, D => 
                           registers_18_17_port, Z => n1995);
   U2727 : HS65_LH_AO22X9 port map( A => n2733, B => n1432, C => n1424, D => 
                           registers_18_18_port, Z => n1996);
   U2728 : HS65_LH_AO22X9 port map( A => n2735, B => n1432, C => n1423, D => 
                           registers_18_19_port, Z => n1997);
   U2729 : HS65_LH_AO22X9 port map( A => n2737, B => n1432, C => n1423, D => 
                           registers_18_20_port, Z => n1998);
   U2730 : HS65_LH_AO22X9 port map( A => n2739, B => n1432, C => n1423, D => 
                           registers_18_21_port, Z => n1999);
   U2731 : HS65_LH_AO22X9 port map( A => n2741, B => n1432, C => n1423, D => 
                           registers_18_22_port, Z => n2000);
   U2732 : HS65_LH_AO22X9 port map( A => n2743, B => n1432, C => n1423, D => 
                           registers_18_23_port, Z => n2001);
   U2733 : HS65_LH_AO22X9 port map( A => n2745, B => n1432, C => n1423, D => 
                           registers_18_24_port, Z => n2002);
   U2734 : HS65_LH_AO22X9 port map( A => n2747, B => n1432, C => n1423, D => 
                           registers_18_25_port, Z => n2003);
   U2735 : HS65_LH_AO22X9 port map( A => n2749, B => n1432, C => n1423, D => 
                           registers_18_26_port, Z => n2004);
   U2736 : HS65_LH_AO22X9 port map( A => n2751, B => n1432, C => n1423, D => 
                           registers_18_27_port, Z => n2005);
   U2737 : HS65_LH_AO22X9 port map( A => n2753, B => n1432, C => n1423, D => 
                           registers_18_28_port, Z => n2006);
   U2738 : HS65_LH_AO22X9 port map( A => n2755, B => n1432, C => n1423, D => 
                           registers_18_29_port, Z => n2007);
   U2739 : HS65_LH_AO22X9 port map( A => n2757, B => n1432, C => n1423, D => 
                           registers_18_30_port, Z => n2008);
   U2740 : HS65_LH_AO22X9 port map( A => n2759, B => n1427, C => n1423, D => 
                           registers_18_31_port, Z => n2009);
   U2741 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n1403, C => n1397, 
                           D => registers_21_0_port, Z => n2074);
   U2742 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n1403, C => n1395, 
                           D => registers_21_1_port, Z => n2075);
   U2743 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n1403, C => n1397, 
                           D => registers_21_2_port, Z => n2076);
   U2744 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n1403, C => n1395, 
                           D => registers_21_3_port, Z => n2077);
   U2745 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n1403, C => n1397, 
                           D => registers_21_4_port, Z => n2078);
   U2746 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n1403, C => n1395, 
                           D => registers_21_5_port, Z => n2079);
   U2747 : HS65_LH_AO22X9 port map( A => n2709, B => n1403, C => n1397, D => 
                           registers_21_6_port, Z => n2080);
   U2748 : HS65_LH_AO22X9 port map( A => n2711, B => n1403, C => n1397, D => 
                           registers_21_7_port, Z => n2081);
   U2749 : HS65_LH_AO22X9 port map( A => n2713, B => n1403, C => n1397, D => 
                           registers_21_8_port, Z => n2082);
   U2750 : HS65_LH_AO22X9 port map( A => n2715, B => n1403, C => n1397, D => 
                           registers_21_9_port, Z => n2083);
   U2751 : HS65_LH_AO22X9 port map( A => n2717, B => n1403, C => n1397, D => 
                           registers_21_10_port, Z => n2084);
   U2752 : HS65_LH_AO22X9 port map( A => n2719, B => n1401, C => n1397, D => 
                           registers_21_11_port, Z => n2085);
   U2753 : HS65_LH_AO22X9 port map( A => n2721, B => n1401, C => n1397, D => 
                           registers_21_12_port, Z => n2086);
   U2754 : HS65_LH_AO22X9 port map( A => n2723, B => n1401, C => n1397, D => 
                           registers_21_13_port, Z => n2087);
   U2755 : HS65_LH_AO22X9 port map( A => n2725, B => n1401, C => n1397, D => 
                           registers_21_14_port, Z => n2088);
   U2756 : HS65_LH_AO22X9 port map( A => n2727, B => n1401, C => n1397, D => 
                           registers_21_15_port, Z => n2089);
   U2757 : HS65_LH_AO22X9 port map( A => n2729, B => n1401, C => n1397, D => 
                           registers_21_16_port, Z => n2090);
   U2758 : HS65_LH_AO22X9 port map( A => n2731, B => n1401, C => n1397, D => 
                           registers_21_17_port, Z => n2091);
   U2759 : HS65_LH_AO22X9 port map( A => n2733, B => n1401, C => n1397, D => 
                           registers_21_18_port, Z => n2092);
   U2760 : HS65_LH_AO22X9 port map( A => n2735, B => n1401, C => n1395, D => 
                           registers_21_19_port, Z => n2093);
   U2761 : HS65_LH_AO22X9 port map( A => n2737, B => n1401, C => n1395, D => 
                           registers_21_20_port, Z => n2094);
   U2762 : HS65_LH_AO22X9 port map( A => n2739, B => n1401, C => n1395, D => 
                           registers_21_21_port, Z => n2095);
   U2763 : HS65_LH_AO22X9 port map( A => n2741, B => n1401, C => n1395, D => 
                           registers_21_22_port, Z => n2096);
   U2764 : HS65_LH_AO22X9 port map( A => n2743, B => n1401, C => n1395, D => 
                           registers_21_23_port, Z => n2097);
   U2765 : HS65_LH_AO22X9 port map( A => n2745, B => n1401, C => n1395, D => 
                           registers_21_24_port, Z => n2098);
   U2766 : HS65_LH_AO22X9 port map( A => n2747, B => n1401, C => n1395, D => 
                           registers_21_25_port, Z => n2099);
   U2767 : HS65_LH_AO22X9 port map( A => n2749, B => n1401, C => n1395, D => 
                           registers_21_26_port, Z => n2100);
   U2768 : HS65_LH_AO22X9 port map( A => n2751, B => n1401, C => n1395, D => 
                           registers_21_27_port, Z => n2101);
   U2769 : HS65_LH_AO22X9 port map( A => n2753, B => n1401, C => n1395, D => 
                           registers_21_28_port, Z => n2102);
   U2770 : HS65_LH_AO22X9 port map( A => n2755, B => n1401, C => n1395, D => 
                           registers_21_29_port, Z => n2103);
   U2771 : HS65_LH_AO22X9 port map( A => n2757, B => n1401, C => n1395, D => 
                           registers_21_30_port, Z => n2104);
   U2772 : HS65_LH_AO22X9 port map( A => n2759, B => n1399, C => n1395, D => 
                           registers_21_31_port, Z => n2105);
   U2773 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n1392, C => n334, D
                           => registers_22_0_port, Z => n2106);
   U2774 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n1392, C => n333, D
                           => registers_22_1_port, Z => n2107);
   U2775 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n1392, C => n334, D
                           => registers_22_2_port, Z => n2108);
   U2776 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n1392, C => n333, D
                           => registers_22_3_port, Z => n2109);
   U2777 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n1392, C => n334, D
                           => registers_22_4_port, Z => n2110);
   U2778 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n1392, C => n333, D
                           => registers_22_5_port, Z => n2111);
   U2779 : HS65_LH_AO22X9 port map( A => n2709, B => n1392, C => n334, D => 
                           registers_22_6_port, Z => n2112);
   U2780 : HS65_LH_AO22X9 port map( A => n2711, B => n1392, C => n334, D => 
                           registers_22_7_port, Z => n2113);
   U2781 : HS65_LH_AO22X9 port map( A => n2713, B => n1392, C => n334, D => 
                           registers_22_8_port, Z => n2114);
   U2782 : HS65_LH_AO22X9 port map( A => n2715, B => n1392, C => n334, D => 
                           registers_22_9_port, Z => n2115);
   U2783 : HS65_LH_AO22X9 port map( A => n2717, B => n1392, C => n334, D => 
                           registers_22_10_port, Z => n2116);
   U2784 : HS65_LH_AO22X9 port map( A => n2719, B => n880, C => n334, D => 
                           registers_22_11_port, Z => n2117);
   U2785 : HS65_LH_AO22X9 port map( A => n2721, B => n880, C => n334, D => 
                           registers_22_12_port, Z => n2118);
   U2786 : HS65_LH_AO22X9 port map( A => n2723, B => n880, C => n334, D => 
                           registers_22_13_port, Z => n2119);
   U2787 : HS65_LH_AO22X9 port map( A => n2725, B => n880, C => n334, D => 
                           registers_22_14_port, Z => n2120);
   U2788 : HS65_LH_AO22X9 port map( A => n2727, B => n880, C => n334, D => 
                           registers_22_15_port, Z => n2121);
   U2789 : HS65_LH_AO22X9 port map( A => n2729, B => n880, C => n334, D => 
                           registers_22_16_port, Z => n2122);
   U2790 : HS65_LH_AO22X9 port map( A => n2731, B => n880, C => n334, D => 
                           registers_22_17_port, Z => n2123);
   U2791 : HS65_LH_AO22X9 port map( A => n2733, B => n880, C => n334, D => 
                           registers_22_18_port, Z => n2124);
   U2792 : HS65_LH_AO22X9 port map( A => n2735, B => n880, C => n333, D => 
                           registers_22_19_port, Z => n2125);
   U2793 : HS65_LH_AO22X9 port map( A => n2737, B => n880, C => n333, D => 
                           registers_22_20_port, Z => n2126);
   U2794 : HS65_LH_AO22X9 port map( A => n2739, B => n880, C => n333, D => 
                           registers_22_21_port, Z => n2127);
   U2795 : HS65_LH_AO22X9 port map( A => n2741, B => n880, C => n333, D => 
                           registers_22_22_port, Z => n2128);
   U2796 : HS65_LH_AO22X9 port map( A => n2743, B => n880, C => n333, D => 
                           registers_22_23_port, Z => n2129);
   U2797 : HS65_LH_AO22X9 port map( A => n2745, B => n880, C => n333, D => 
                           registers_22_24_port, Z => n2130);
   U2798 : HS65_LH_AO22X9 port map( A => n2747, B => n880, C => n333, D => 
                           registers_22_25_port, Z => n2131);
   U2799 : HS65_LH_AO22X9 port map( A => n2749, B => n880, C => n333, D => 
                           registers_22_26_port, Z => n2132);
   U2800 : HS65_LH_AO22X9 port map( A => n2751, B => n880, C => n333, D => 
                           registers_22_27_port, Z => n2133);
   U2801 : HS65_LH_AO22X9 port map( A => n2753, B => n880, C => n333, D => 
                           registers_22_28_port, Z => n2134);
   U2802 : HS65_LH_AO22X9 port map( A => n2755, B => n880, C => n333, D => 
                           registers_22_29_port, Z => n2135);
   U2803 : HS65_LH_AO22X9 port map( A => n2757, B => n880, C => n333, D => 
                           registers_22_30_port, Z => n2136);
   U2804 : HS65_LH_AO22X9 port map( A => n2759, B => n352, C => n333, D => 
                           registers_22_31_port, Z => n2137);
   U2805 : HS65_LH_AO22X9 port map( A => n2697, B => n2495, C => n2492, D => 
                           registers_4_0_port, Z => n1530);
   U2806 : HS65_LH_AO22X9 port map( A => n2699, B => n2495, C => n2491, D => 
                           registers_4_1_port, Z => n1531);
   U2807 : HS65_LH_AO22X9 port map( A => n2701, B => n2495, C => n2492, D => 
                           registers_4_2_port, Z => n1532);
   U2808 : HS65_LH_AO22X9 port map( A => n2703, B => n2495, C => n2491, D => 
                           registers_4_3_port, Z => n1533);
   U2809 : HS65_LH_AO22X9 port map( A => n2705, B => n2495, C => n2492, D => 
                           registers_4_4_port, Z => n1534);
   U2810 : HS65_LH_AO22X9 port map( A => n2707, B => n2495, C => n2491, D => 
                           registers_4_5_port, Z => n1535);
   U2811 : HS65_LH_AO22X9 port map( A => regfile_i(9), B => n2495, C => n2492, 
                           D => registers_4_6_port, Z => n1536);
   U2812 : HS65_LH_AO22X9 port map( A => regfile_i(10), B => n2495, C => n2492,
                           D => registers_4_7_port, Z => n1537);
   U2813 : HS65_LH_AO22X9 port map( A => regfile_i(11), B => n2495, C => n2492,
                           D => registers_4_8_port, Z => n1538);
   U2814 : HS65_LH_AO22X9 port map( A => regfile_i(12), B => n2495, C => n2492,
                           D => registers_4_9_port, Z => n1539);
   U2815 : HS65_LH_AO22X9 port map( A => regfile_i(13), B => n2495, C => n2492,
                           D => registers_4_10_port, Z => n1540);
   U2816 : HS65_LH_AO22X9 port map( A => regfile_i(14), B => n2494, C => n2492,
                           D => registers_4_11_port, Z => n1541);
   U2817 : HS65_LH_AO22X9 port map( A => regfile_i(15), B => n2494, C => n2492,
                           D => registers_4_12_port, Z => n1542);
   U2818 : HS65_LH_AO22X9 port map( A => regfile_i(16), B => n2494, C => n2492,
                           D => registers_4_13_port, Z => n1543);
   U2819 : HS65_LH_AO22X9 port map( A => regfile_i(17), B => n2494, C => n2492,
                           D => registers_4_14_port, Z => n1544);
   U2820 : HS65_LH_AO22X9 port map( A => regfile_i(18), B => n2494, C => n2492,
                           D => registers_4_15_port, Z => n1545);
   U2821 : HS65_LH_AO22X9 port map( A => regfile_i(19), B => n2494, C => n2492,
                           D => registers_4_16_port, Z => n1546);
   U2822 : HS65_LH_AO22X9 port map( A => regfile_i(20), B => n2494, C => n2492,
                           D => registers_4_17_port, Z => n1547);
   U2823 : HS65_LH_AO22X9 port map( A => regfile_i(21), B => n2494, C => n2492,
                           D => registers_4_18_port, Z => n1548);
   U2824 : HS65_LH_AO22X9 port map( A => regfile_i(22), B => n2494, C => n2491,
                           D => registers_4_19_port, Z => n1549);
   U2825 : HS65_LH_AO22X9 port map( A => regfile_i(23), B => n2494, C => n2491,
                           D => registers_4_20_port, Z => n1550);
   U2826 : HS65_LH_AO22X9 port map( A => regfile_i(24), B => n2494, C => n2491,
                           D => registers_4_21_port, Z => n1551);
   U2827 : HS65_LH_AO22X9 port map( A => regfile_i(25), B => n2494, C => n2491,
                           D => registers_4_22_port, Z => n1552);
   U2828 : HS65_LH_AO22X9 port map( A => regfile_i(26), B => n2494, C => n2491,
                           D => registers_4_23_port, Z => n1553);
   U2829 : HS65_LH_AO22X9 port map( A => regfile_i(27), B => n2494, C => n2491,
                           D => registers_4_24_port, Z => n1554);
   U2830 : HS65_LH_AO22X9 port map( A => regfile_i(28), B => n2494, C => n2491,
                           D => registers_4_25_port, Z => n1555);
   U2831 : HS65_LH_AO22X9 port map( A => regfile_i(29), B => n2494, C => n2491,
                           D => registers_4_26_port, Z => n1556);
   U2832 : HS65_LH_AO22X9 port map( A => regfile_i(30), B => n2494, C => n2491,
                           D => registers_4_27_port, Z => n1557);
   U2833 : HS65_LH_AO22X9 port map( A => regfile_i(31), B => n2494, C => n2491,
                           D => registers_4_28_port, Z => n1558);
   U2834 : HS65_LH_AO22X9 port map( A => regfile_i(32), B => n2494, C => n2491,
                           D => registers_4_29_port, Z => n1559);
   U2835 : HS65_LH_AO22X9 port map( A => regfile_i(33), B => n2494, C => n2491,
                           D => registers_4_30_port, Z => n1560);
   U2836 : HS65_LH_AO22X9 port map( A => regfile_i(34), B => n2493, C => n2491,
                           D => registers_4_31_port, Z => n1561);
   U2837 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n2434, C => n2431, 
                           D => registers_16_0_port, Z => n1914);
   U2838 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n2434, C => n2431, 
                           D => registers_16_1_port, Z => n1915);
   U2839 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n2434, C => n2431, 
                           D => registers_16_2_port, Z => n1916);
   U2840 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n2434, C => n2431, 
                           D => registers_16_3_port, Z => n1917);
   U2841 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n2434, C => n2431, 
                           D => registers_16_4_port, Z => n1918);
   U2842 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n2434, C => n2431, 
                           D => registers_16_5_port, Z => n1919);
   U2843 : HS65_LH_AO22X9 port map( A => n2709, B => n2434, C => n2431, D => 
                           registers_16_6_port, Z => n1920);
   U2844 : HS65_LH_AO22X9 port map( A => n2711, B => n2434, C => n2431, D => 
                           registers_16_7_port, Z => n1921);
   U2845 : HS65_LH_AO22X9 port map( A => n2713, B => n2434, C => n2431, D => 
                           registers_16_8_port, Z => n1922);
   U2846 : HS65_LH_AO22X9 port map( A => n2715, B => n2434, C => n2431, D => 
                           registers_16_9_port, Z => n1923);
   U2847 : HS65_LH_AO22X9 port map( A => n2717, B => n2434, C => n2431, D => 
                           registers_16_10_port, Z => n1924);
   U2848 : HS65_LH_AO22X9 port map( A => n2719, B => n2433, C => n2431, D => 
                           registers_16_11_port, Z => n1925);
   U2849 : HS65_LH_AO22X9 port map( A => n2721, B => n2433, C => n2431, D => 
                           registers_16_12_port, Z => n1926);
   U2850 : HS65_LH_AO22X9 port map( A => n2723, B => n2433, C => n2431, D => 
                           registers_16_13_port, Z => n1927);
   U2851 : HS65_LH_AO22X9 port map( A => n2725, B => n2433, C => n2431, D => 
                           registers_16_14_port, Z => n1928);
   U2852 : HS65_LH_AO22X9 port map( A => n2727, B => n2433, C => n2431, D => 
                           registers_16_15_port, Z => n1929);
   U2853 : HS65_LH_AO22X9 port map( A => n2729, B => n2433, C => n2431, D => 
                           registers_16_16_port, Z => n1930);
   U2854 : HS65_LH_AO22X9 port map( A => n2731, B => n2433, C => n2431, D => 
                           registers_16_17_port, Z => n1931);
   U2855 : HS65_LH_AO22X9 port map( A => n2733, B => n2433, C => n2431, D => 
                           registers_16_18_port, Z => n1932);
   U2856 : HS65_LH_AO22X9 port map( A => n2735, B => n2433, C => n2431, D => 
                           registers_16_19_port, Z => n1933);
   U2857 : HS65_LH_AO22X9 port map( A => n2737, B => n2433, C => n1416, D => 
                           registers_16_20_port, Z => n1934);
   U2858 : HS65_LH_AO22X9 port map( A => n2739, B => n2433, C => n1416, D => 
                           registers_16_21_port, Z => n1935);
   U2859 : HS65_LH_AO22X9 port map( A => n2741, B => n2433, C => n1416, D => 
                           registers_16_22_port, Z => n1936);
   U2860 : HS65_LH_AO22X9 port map( A => n2743, B => n2433, C => n1416, D => 
                           registers_16_23_port, Z => n1937);
   U2861 : HS65_LH_AO22X9 port map( A => n2745, B => n2433, C => n1416, D => 
                           registers_16_24_port, Z => n1938);
   U2862 : HS65_LH_AO22X9 port map( A => n2747, B => n2433, C => n1416, D => 
                           registers_16_25_port, Z => n1939);
   U2863 : HS65_LH_AO22X9 port map( A => n2749, B => n2433, C => n1416, D => 
                           registers_16_26_port, Z => n1940);
   U2864 : HS65_LH_AO22X9 port map( A => n2751, B => n2433, C => n1416, D => 
                           registers_16_27_port, Z => n1941);
   U2865 : HS65_LH_AO22X9 port map( A => n2753, B => n2433, C => n1416, D => 
                           registers_16_28_port, Z => n1942);
   U2866 : HS65_LH_AO22X9 port map( A => n2755, B => n2433, C => n1416, D => 
                           registers_16_29_port, Z => n1943);
   U2867 : HS65_LH_AO22X9 port map( A => n2757, B => n2433, C => n1416, D => 
                           registers_16_30_port, Z => n1944);
   U2868 : HS65_LH_AO22X9 port map( A => n2759, B => n2432, C => n1416, D => 
                           registers_16_31_port, Z => n1945);
   U2869 : HS65_LH_AO22X9 port map( A => regfile_i(3), B => n1413, C => n1410, 
                           D => registers_20_0_port, Z => n2042);
   U2870 : HS65_LH_AO22X9 port map( A => regfile_i(4), B => n1413, C => n1405, 
                           D => registers_20_1_port, Z => n2043);
   U2871 : HS65_LH_AO22X9 port map( A => regfile_i(5), B => n1413, C => n1410, 
                           D => registers_20_2_port, Z => n2044);
   U2872 : HS65_LH_AO22X9 port map( A => regfile_i(6), B => n1413, C => n1405, 
                           D => registers_20_3_port, Z => n2045);
   U2873 : HS65_LH_AO22X9 port map( A => regfile_i(7), B => n1413, C => n1410, 
                           D => registers_20_4_port, Z => n2046);
   U2874 : HS65_LH_AO22X9 port map( A => regfile_i(8), B => n1413, C => n1405, 
                           D => registers_20_5_port, Z => n2047);
   U2875 : HS65_LH_AO22X9 port map( A => n2709, B => n1413, C => n1410, D => 
                           registers_20_6_port, Z => n2048);
   U2876 : HS65_LH_AO22X9 port map( A => n2711, B => n1413, C => n1410, D => 
                           registers_20_7_port, Z => n2049);
   U2877 : HS65_LH_AO22X9 port map( A => n2713, B => n1413, C => n1410, D => 
                           registers_20_8_port, Z => n2050);
   U2878 : HS65_LH_AO22X9 port map( A => n2715, B => n1413, C => n1410, D => 
                           registers_20_9_port, Z => n2051);
   U2879 : HS65_LH_AO22X9 port map( A => n2717, B => n1413, C => n1410, D => 
                           registers_20_10_port, Z => n2052);
   U2880 : HS65_LH_AO22X9 port map( A => n2719, B => n1412, C => n1410, D => 
                           registers_20_11_port, Z => n2053);
   U2881 : HS65_LH_AO22X9 port map( A => n2721, B => n1412, C => n1410, D => 
                           registers_20_12_port, Z => n2054);
   U2882 : HS65_LH_AO22X9 port map( A => n2723, B => n1412, C => n1410, D => 
                           registers_20_13_port, Z => n2055);
   U2883 : HS65_LH_AO22X9 port map( A => n2725, B => n1412, C => n1410, D => 
                           registers_20_14_port, Z => n2056);
   U2884 : HS65_LH_AO22X9 port map( A => n2727, B => n1412, C => n1410, D => 
                           registers_20_15_port, Z => n2057);
   U2885 : HS65_LH_AO22X9 port map( A => n2729, B => n1412, C => n1410, D => 
                           registers_20_16_port, Z => n2058);
   U2886 : HS65_LH_AO22X9 port map( A => n2731, B => n1412, C => n1410, D => 
                           registers_20_17_port, Z => n2059);
   U2887 : HS65_LH_AO22X9 port map( A => n2733, B => n1412, C => n1410, D => 
                           registers_20_18_port, Z => n2060);
   U2888 : HS65_LH_AO22X9 port map( A => n2735, B => n1412, C => n1405, D => 
                           registers_20_19_port, Z => n2061);
   U2889 : HS65_LH_AO22X9 port map( A => n2737, B => n1412, C => n1405, D => 
                           registers_20_20_port, Z => n2062);
   U2890 : HS65_LH_AO22X9 port map( A => n2739, B => n1412, C => n1405, D => 
                           registers_20_21_port, Z => n2063);
   U2891 : HS65_LH_AO22X9 port map( A => n2741, B => n1412, C => n1405, D => 
                           registers_20_22_port, Z => n2064);
   U2892 : HS65_LH_AO22X9 port map( A => n2743, B => n1412, C => n1405, D => 
                           registers_20_23_port, Z => n2065);
   U2893 : HS65_LH_AO22X9 port map( A => n2745, B => n1412, C => n1405, D => 
                           registers_20_24_port, Z => n2066);
   U2894 : HS65_LH_AO22X9 port map( A => n2747, B => n1412, C => n1405, D => 
                           registers_20_25_port, Z => n2067);
   U2895 : HS65_LH_AO22X9 port map( A => n2749, B => n1412, C => n1405, D => 
                           registers_20_26_port, Z => n2068);
   U2896 : HS65_LH_AO22X9 port map( A => n2751, B => n1412, C => n1405, D => 
                           registers_20_27_port, Z => n2069);
   U2897 : HS65_LH_AO22X9 port map( A => n2753, B => n1412, C => n1405, D => 
                           registers_20_28_port, Z => n2070);
   U2898 : HS65_LH_AO22X9 port map( A => n2755, B => n1412, C => n1405, D => 
                           registers_20_29_port, Z => n2071);
   U2899 : HS65_LH_AO22X9 port map( A => n2757, B => n1412, C => n1405, D => 
                           registers_20_30_port, Z => n2072);
   U2900 : HS65_LH_AO22X9 port map( A => n2759, B => n1411, C => n1405, D => 
                           registers_20_31_port, Z => n2073);
   U2901 : HS65_LH_NOR3X4 port map( A => regfile_i(35), B => regfile_i(37), C 
                           => n2896, Z => n1396);
   U2902 : HS65_LH_NOR3X4 port map( A => n2897, B => regfile_i(37), C => n2896,
                           Z => n1398);
   U2903 : HS65_LH_NOR3X4 port map( A => regfile_i(36), B => regfile_i(37), C 
                           => n2897, Z => n1393);
   U2904 : HS65_LH_IVX9 port map( A => regfile_i(35), Z => n2897);
   U2905 : HS65_LH_IVX9 port map( A => regfile_i(36), Z => n2896);
   U2906 : HS65_LH_IVX9 port map( A => regfile_i(38), Z => n2895);
   U2907 : HS65_LH_NOR3X4 port map( A => regfile_i(36), B => regfile_i(37), C 
                           => regfile_i(35), Z => n1391);
   U2908 : HS65_LH_AND3X9 port map( A => regfile_i(0), B => n2895, C => 
                           regfile_i(39), Z => n1417);
   U2909 : HS65_LH_AND3X9 port map( A => regfile_i(38), B => regfile_i(0), C =>
                           regfile_i(39), Z => n1426);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity pc is

   port( clk, rst_n, halt_i : in std_logic;  npc_i : in std_logic_vector (11 
         downto 0);  pc_o : out std_logic_vector (11 downto 0));

end pc;

architecture SYN_behavioral of pc is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPSQX9
      port( D, CP, SN : in std_logic;  Q : out std_logic);
   end component;
   
   signal pc_o_11_port, pc_o_10_port, pc_o_9_port, pc_o_8_port, pc_o_7_port, 
      pc_o_6_port, pc_o_5_port, pc_o_4_port, pc_o_3_port, pc_o_2_port, 
      pc_o_1_port, pc_o_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n1 : std_logic;

begin
   pc_o <= ( pc_o_11_port, pc_o_10_port, pc_o_9_port, pc_o_8_port, pc_o_7_port,
      pc_o_6_port, pc_o_5_port, pc_o_4_port, pc_o_3_port, pc_o_2_port, 
      pc_o_1_port, pc_o_0_port );
   
   pc_c_reg_11_inst : HS65_LH_DFPSQX9 port map( D => n13, CP => clk, SN => 
                           rst_n, Q => pc_o_11_port);
   pc_c_reg_10_inst : HS65_LH_DFPSQX9 port map( D => n12, CP => clk, SN => 
                           rst_n, Q => pc_o_10_port);
   pc_c_reg_9_inst : HS65_LH_DFPSQX9 port map( D => n11, CP => clk, SN => rst_n
                           , Q => pc_o_9_port);
   pc_c_reg_8_inst : HS65_LH_DFPSQX9 port map( D => n10, CP => clk, SN => rst_n
                           , Q => pc_o_8_port);
   pc_c_reg_7_inst : HS65_LH_DFPSQX9 port map( D => n9, CP => clk, SN => rst_n,
                           Q => pc_o_7_port);
   pc_c_reg_6_inst : HS65_LH_DFPSQX9 port map( D => n8, CP => clk, SN => rst_n,
                           Q => pc_o_6_port);
   pc_c_reg_5_inst : HS65_LH_DFPSQX9 port map( D => n7, CP => clk, SN => rst_n,
                           Q => pc_o_5_port);
   pc_c_reg_4_inst : HS65_LH_DFPSQX9 port map( D => n6, CP => clk, SN => rst_n,
                           Q => pc_o_4_port);
   pc_c_reg_3_inst : HS65_LH_DFPSQX9 port map( D => n5, CP => clk, SN => rst_n,
                           Q => pc_o_3_port);
   pc_c_reg_2_inst : HS65_LH_DFPSQX9 port map( D => n4, CP => clk, SN => rst_n,
                           Q => pc_o_2_port);
   pc_c_reg_1_inst : HS65_LH_DFPSQX9 port map( D => n3, CP => clk, SN => rst_n,
                           Q => pc_o_1_port);
   pc_c_reg_0_inst : HS65_LH_DFPSQX9 port map( D => n2, CP => clk, SN => rst_n,
                           Q => pc_o_0_port);
   U2 : HS65_LH_AO22X9 port map( A => pc_o_9_port, B => halt_i, C => npc_i(9), 
                           D => n1, Z => n11);
   U3 : HS65_LH_AO22X9 port map( A => pc_o_0_port, B => halt_i, C => npc_i(0), 
                           D => n1, Z => n2);
   U4 : HS65_LH_AO22X9 port map( A => pc_o_1_port, B => halt_i, C => npc_i(1), 
                           D => n1, Z => n3);
   U5 : HS65_LH_AO22X9 port map( A => pc_o_2_port, B => halt_i, C => npc_i(2), 
                           D => n1, Z => n4);
   U6 : HS65_LH_AO22X9 port map( A => pc_o_3_port, B => halt_i, C => npc_i(3), 
                           D => n1, Z => n5);
   U7 : HS65_LH_AO22X9 port map( A => pc_o_4_port, B => halt_i, C => npc_i(4), 
                           D => n1, Z => n6);
   U8 : HS65_LH_AO22X9 port map( A => pc_o_5_port, B => halt_i, C => npc_i(5), 
                           D => n1, Z => n7);
   U9 : HS65_LH_AO22X9 port map( A => pc_o_6_port, B => halt_i, C => npc_i(6), 
                           D => n1, Z => n8);
   U10 : HS65_LH_AO22X9 port map( A => pc_o_7_port, B => halt_i, C => npc_i(7),
                           D => n1, Z => n9);
   U11 : HS65_LH_AO22X9 port map( A => pc_o_8_port, B => halt_i, C => npc_i(8),
                           D => n1, Z => n10);
   U12 : HS65_LH_AO22X9 port map( A => pc_o_10_port, B => halt_i, C => 
                           npc_i(10), D => n1, Z => n12);
   U13 : HS65_LH_AO22X9 port map( A => pc_o_11_port, B => halt_i, C => 
                           npc_i(11), D => n1, Z => n13);
   U14 : HS65_LH_IVX9 port map( A => halt_i, Z => n1);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity mem_wb is

   port( clk, rst_n, halt_i : in std_logic;  MEM_WB_i : in std_logic_vector (38
         downto 0);  MEM_WB_o : out std_logic_vector (38 downto 0));

end mem_wb;

architecture SYN_Behavioral of mem_wb is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal MEM_WB_o_ALU_RES_31_port, MEM_WB_o_ALU_RES_30_port, 
      MEM_WB_o_ALU_RES_29_port, MEM_WB_o_ALU_RES_28_port, 
      MEM_WB_o_ALU_RES_27_port, MEM_WB_o_ALU_RES_26_port, 
      MEM_WB_o_ALU_RES_25_port, MEM_WB_o_ALU_RES_24_port, 
      MEM_WB_o_ALU_RES_23_port, MEM_WB_o_ALU_RES_22_port, 
      MEM_WB_o_ALU_RES_21_port, MEM_WB_o_ALU_RES_20_port, 
      MEM_WB_o_ALU_RES_19_port, MEM_WB_o_ALU_RES_18_port, 
      MEM_WB_o_ALU_RES_17_port, MEM_WB_o_ALU_RES_16_port, 
      MEM_WB_o_ALU_RES_15_port, MEM_WB_o_ALU_RES_14_port, 
      MEM_WB_o_ALU_RES_13_port, MEM_WB_o_ALU_RES_12_port, 
      MEM_WB_o_ALU_RES_11_port, MEM_WB_o_ALU_RES_10_port, 
      MEM_WB_o_ALU_RES_9_port, MEM_WB_o_ALU_RES_8_port, MEM_WB_o_ALU_RES_7_port
      , MEM_WB_o_ALU_RES_6_port, MEM_WB_o_ALU_RES_5_port, 
      MEM_WB_o_ALU_RES_4_port, MEM_WB_o_ALU_RES_3_port, MEM_WB_o_ALU_RES_2_port
      , MEM_WB_o_ALU_RES_1_port, MEM_WB_o_ALU_RES_0_port, 
      MEM_WB_o_WRITE_REG_4_port, MEM_WB_o_WRITE_REG_3_port, 
      MEM_WB_o_WRITE_REG_2_port, MEM_WB_o_WRITE_REG_1_port, 
      MEM_WB_o_WRITE_REG_0_port, MEM_WB_o_MEMTOREG_port, MEM_WB_o_REGWRITE_port
      , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n1, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52 : std_logic;

begin
   MEM_WB_o <= ( MEM_WB_o_ALU_RES_31_port, MEM_WB_o_ALU_RES_30_port, 
      MEM_WB_o_ALU_RES_29_port, MEM_WB_o_ALU_RES_28_port, 
      MEM_WB_o_ALU_RES_27_port, MEM_WB_o_ALU_RES_26_port, 
      MEM_WB_o_ALU_RES_25_port, MEM_WB_o_ALU_RES_24_port, 
      MEM_WB_o_ALU_RES_23_port, MEM_WB_o_ALU_RES_22_port, 
      MEM_WB_o_ALU_RES_21_port, MEM_WB_o_ALU_RES_20_port, 
      MEM_WB_o_ALU_RES_19_port, MEM_WB_o_ALU_RES_18_port, 
      MEM_WB_o_ALU_RES_17_port, MEM_WB_o_ALU_RES_16_port, 
      MEM_WB_o_ALU_RES_15_port, MEM_WB_o_ALU_RES_14_port, 
      MEM_WB_o_ALU_RES_13_port, MEM_WB_o_ALU_RES_12_port, 
      MEM_WB_o_ALU_RES_11_port, MEM_WB_o_ALU_RES_10_port, 
      MEM_WB_o_ALU_RES_9_port, MEM_WB_o_ALU_RES_8_port, MEM_WB_o_ALU_RES_7_port
      , MEM_WB_o_ALU_RES_6_port, MEM_WB_o_ALU_RES_5_port, 
      MEM_WB_o_ALU_RES_4_port, MEM_WB_o_ALU_RES_3_port, MEM_WB_o_ALU_RES_2_port
      , MEM_WB_o_ALU_RES_1_port, MEM_WB_o_ALU_RES_0_port, 
      MEM_WB_o_WRITE_REG_4_port, MEM_WB_o_WRITE_REG_3_port, 
      MEM_WB_o_WRITE_REG_2_port, MEM_WB_o_WRITE_REG_1_port, 
      MEM_WB_o_WRITE_REG_0_port, MEM_WB_o_MEMTOREG_port, MEM_WB_o_REGWRITE_port
      );
   
   mem_wb_c_reg_ALU_RES_31_inst : HS65_LH_DFPRQX9 port map( D => n40, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_31_port);
   mem_wb_c_reg_ALU_RES_30_inst : HS65_LH_DFPRQX9 port map( D => n39, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_30_port);
   mem_wb_c_reg_ALU_RES_29_inst : HS65_LH_DFPRQX9 port map( D => n38, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_29_port);
   mem_wb_c_reg_ALU_RES_28_inst : HS65_LH_DFPRQX9 port map( D => n37, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_28_port);
   mem_wb_c_reg_ALU_RES_27_inst : HS65_LH_DFPRQX9 port map( D => n36, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_27_port);
   mem_wb_c_reg_ALU_RES_26_inst : HS65_LH_DFPRQX9 port map( D => n35, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_26_port);
   mem_wb_c_reg_ALU_RES_25_inst : HS65_LH_DFPRQX9 port map( D => n34, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_25_port);
   mem_wb_c_reg_ALU_RES_24_inst : HS65_LH_DFPRQX9 port map( D => n33, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_24_port);
   mem_wb_c_reg_ALU_RES_23_inst : HS65_LH_DFPRQX9 port map( D => n32, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_23_port);
   mem_wb_c_reg_ALU_RES_22_inst : HS65_LH_DFPRQX9 port map( D => n31, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_22_port);
   mem_wb_c_reg_ALU_RES_21_inst : HS65_LH_DFPRQX9 port map( D => n30, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_21_port);
   mem_wb_c_reg_ALU_RES_20_inst : HS65_LH_DFPRQX9 port map( D => n29, CP => clk
                           , RN => n48, Q => MEM_WB_o_ALU_RES_20_port);
   mem_wb_c_reg_ALU_RES_19_inst : HS65_LH_DFPRQX9 port map( D => n28, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_19_port);
   mem_wb_c_reg_ALU_RES_18_inst : HS65_LH_DFPRQX9 port map( D => n27, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_18_port);
   mem_wb_c_reg_ALU_RES_17_inst : HS65_LH_DFPRQX9 port map( D => n26, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_17_port);
   mem_wb_c_reg_ALU_RES_16_inst : HS65_LH_DFPRQX9 port map( D => n25, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_16_port);
   mem_wb_c_reg_ALU_RES_15_inst : HS65_LH_DFPRQX9 port map( D => n24, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_15_port);
   mem_wb_c_reg_ALU_RES_14_inst : HS65_LH_DFPRQX9 port map( D => n23, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_14_port);
   mem_wb_c_reg_ALU_RES_13_inst : HS65_LH_DFPRQX9 port map( D => n22, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_13_port);
   mem_wb_c_reg_ALU_RES_12_inst : HS65_LH_DFPRQX9 port map( D => n21, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_12_port);
   mem_wb_c_reg_ALU_RES_11_inst : HS65_LH_DFPRQX9 port map( D => n20, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_11_port);
   mem_wb_c_reg_ALU_RES_10_inst : HS65_LH_DFPRQX9 port map( D => n19, CP => clk
                           , RN => n49, Q => MEM_WB_o_ALU_RES_10_port);
   mem_wb_c_reg_ALU_RES_9_inst : HS65_LH_DFPRQX9 port map( D => n18, CP => clk,
                           RN => n49, Q => MEM_WB_o_ALU_RES_9_port);
   mem_wb_c_reg_ALU_RES_8_inst : HS65_LH_DFPRQX9 port map( D => n17, CP => clk,
                           RN => n49, Q => MEM_WB_o_ALU_RES_8_port);
   mem_wb_c_reg_ALU_RES_7_inst : HS65_LH_DFPRQX9 port map( D => n16, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_7_port);
   mem_wb_c_reg_ALU_RES_6_inst : HS65_LH_DFPRQX9 port map( D => n15, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_6_port);
   mem_wb_c_reg_ALU_RES_5_inst : HS65_LH_DFPRQX9 port map( D => n14, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_5_port);
   mem_wb_c_reg_ALU_RES_4_inst : HS65_LH_DFPRQX9 port map( D => n13, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_4_port);
   mem_wb_c_reg_ALU_RES_3_inst : HS65_LH_DFPRQX9 port map( D => n12, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_3_port);
   mem_wb_c_reg_ALU_RES_2_inst : HS65_LH_DFPRQX9 port map( D => n11, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_2_port);
   mem_wb_c_reg_ALU_RES_1_inst : HS65_LH_DFPRQX9 port map( D => n10, CP => clk,
                           RN => n50, Q => MEM_WB_o_ALU_RES_1_port);
   mem_wb_c_reg_ALU_RES_0_inst : HS65_LH_DFPRQX9 port map( D => n9, CP => clk, 
                           RN => n50, Q => MEM_WB_o_ALU_RES_0_port);
   mem_wb_c_reg_WRITE_REG_4_inst : HS65_LH_DFPRQX9 port map( D => n8, CP => clk
                           , RN => n50, Q => MEM_WB_o_WRITE_REG_4_port);
   mem_wb_c_reg_WRITE_REG_3_inst : HS65_LH_DFPRQX9 port map( D => n7, CP => clk
                           , RN => n50, Q => MEM_WB_o_WRITE_REG_3_port);
   mem_wb_c_reg_WRITE_REG_2_inst : HS65_LH_DFPRQX9 port map( D => n6, CP => clk
                           , RN => n50, Q => MEM_WB_o_WRITE_REG_2_port);
   mem_wb_c_reg_WRITE_REG_1_inst : HS65_LH_DFPRQX9 port map( D => n5, CP => clk
                           , RN => n50, Q => MEM_WB_o_WRITE_REG_1_port);
   mem_wb_c_reg_WRITE_REG_0_inst : HS65_LH_DFPRQX9 port map( D => n4, CP => clk
                           , RN => n51, Q => MEM_WB_o_WRITE_REG_0_port);
   mem_wb_c_reg_MEMTOREG_inst : HS65_LH_DFPRQX9 port map( D => n3, CP => clk, 
                           RN => n51, Q => MEM_WB_o_MEMTOREG_port);
   mem_wb_c_reg_REGWRITE_inst : HS65_LH_DFPRQX9 port map( D => n2, CP => clk, 
                           RN => n51, Q => MEM_WB_o_REGWRITE_port);
   U2 : HS65_LH_BFX9 port map( A => n47, Z => n50);
   U3 : HS65_LH_BFX9 port map( A => n46, Z => n49);
   U4 : HS65_LH_BFX9 port map( A => n46, Z => n48);
   U5 : HS65_LH_BFX9 port map( A => n47, Z => n51);
   U6 : HS65_LH_BFX9 port map( A => rst_n, Z => n47);
   U7 : HS65_LH_BFX9 port map( A => rst_n, Z => n46);
   U8 : HS65_LH_BFX9 port map( A => n1, Z => n42);
   U9 : HS65_LH_BFX9 port map( A => n1, Z => n43);
   U10 : HS65_LH_BFX9 port map( A => n41, Z => n44);
   U11 : HS65_LH_BFX9 port map( A => n41, Z => n45);
   U12 : HS65_LH_BFX9 port map( A => n52, Z => n1);
   U13 : HS65_LH_BFX9 port map( A => n52, Z => n41);
   U14 : HS65_LH_AO22X9 port map( A => MEM_WB_o_WRITE_REG_2_port, B => halt_i, 
                           C => MEM_WB_i(4), D => n42, Z => n6);
   U15 : HS65_LH_AO22X9 port map( A => MEM_WB_o_WRITE_REG_4_port, B => halt_i, 
                           C => MEM_WB_i(6), D => n42, Z => n8);
   U16 : HS65_LH_AO22X9 port map( A => MEM_WB_o_WRITE_REG_0_port, B => halt_i, 
                           C => MEM_WB_i(2), D => n42, Z => n4);
   U17 : HS65_LH_AO22X9 port map( A => MEM_WB_o_WRITE_REG_3_port, B => halt_i, 
                           C => MEM_WB_i(5), D => n42, Z => n7);
   U18 : HS65_LH_AO22X9 port map( A => MEM_WB_o_WRITE_REG_1_port, B => halt_i, 
                           C => MEM_WB_i(3), D => n42, Z => n5);
   U19 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_0_port, B => halt_i, C 
                           => MEM_WB_i(7), D => n42, Z => n9);
   U20 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_1_port, B => halt_i, C 
                           => MEM_WB_i(8), D => n42, Z => n10);
   U21 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_2_port, B => halt_i, C 
                           => MEM_WB_i(9), D => n42, Z => n11);
   U22 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_3_port, B => halt_i, C 
                           => MEM_WB_i(10), D => n42, Z => n12);
   U23 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_4_port, B => halt_i, C 
                           => MEM_WB_i(11), D => n42, Z => n13);
   U24 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_5_port, B => halt_i, C 
                           => MEM_WB_i(12), D => n43, Z => n14);
   U25 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_6_port, B => halt_i, C 
                           => MEM_WB_i(13), D => n43, Z => n15);
   U26 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_7_port, B => halt_i, C 
                           => MEM_WB_i(14), D => n43, Z => n16);
   U27 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_8_port, B => halt_i, C 
                           => MEM_WB_i(15), D => n43, Z => n17);
   U28 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_9_port, B => halt_i, C 
                           => MEM_WB_i(16), D => n43, Z => n18);
   U29 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_10_port, B => halt_i, C
                           => MEM_WB_i(17), D => n43, Z => n19);
   U30 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_11_port, B => halt_i, C
                           => MEM_WB_i(18), D => n43, Z => n20);
   U31 : HS65_LH_AO22X9 port map( A => halt_i, B => MEM_WB_o_REGWRITE_port, C 
                           => MEM_WB_i(0), D => n42, Z => n2);
   U32 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_12_port, B => halt_i, C
                           => MEM_WB_i(19), D => n43, Z => n21);
   U33 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_13_port, B => halt_i, C
                           => MEM_WB_i(20), D => n43, Z => n22);
   U34 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_14_port, B => halt_i, C
                           => MEM_WB_i(21), D => n43, Z => n23);
   U35 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_15_port, B => halt_i, C
                           => MEM_WB_i(22), D => n43, Z => n24);
   U36 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_16_port, B => halt_i, C
                           => MEM_WB_i(23), D => n43, Z => n25);
   U37 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_17_port, B => halt_i, C
                           => MEM_WB_i(24), D => n44, Z => n26);
   U38 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_18_port, B => halt_i, C
                           => MEM_WB_i(25), D => n44, Z => n27);
   U39 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_19_port, B => halt_i, C
                           => MEM_WB_i(26), D => n44, Z => n28);
   U40 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_20_port, B => halt_i, C
                           => MEM_WB_i(27), D => n44, Z => n29);
   U41 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_21_port, B => halt_i, C
                           => MEM_WB_i(28), D => n44, Z => n30);
   U42 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_22_port, B => halt_i, C
                           => MEM_WB_i(29), D => n44, Z => n31);
   U43 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_23_port, B => halt_i, C
                           => MEM_WB_i(30), D => n44, Z => n32);
   U44 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_24_port, B => halt_i, C
                           => MEM_WB_i(31), D => n44, Z => n33);
   U45 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_25_port, B => halt_i, C
                           => MEM_WB_i(32), D => n44, Z => n34);
   U46 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_26_port, B => halt_i, C
                           => MEM_WB_i(33), D => n44, Z => n35);
   U47 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_27_port, B => halt_i, C
                           => MEM_WB_i(34), D => n44, Z => n36);
   U48 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_28_port, B => halt_i, C
                           => MEM_WB_i(35), D => n44, Z => n37);
   U49 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_29_port, B => halt_i, C
                           => MEM_WB_i(36), D => n45, Z => n38);
   U50 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_30_port, B => halt_i, C
                           => MEM_WB_i(37), D => n45, Z => n39);
   U51 : HS65_LH_AO22X9 port map( A => MEM_WB_o_ALU_RES_31_port, B => halt_i, C
                           => MEM_WB_i(38), D => n45, Z => n40);
   U52 : HS65_LH_AO22X9 port map( A => MEM_WB_o_MEMTOREG_port, B => halt_i, C 
                           => MEM_WB_i(1), D => n42, Z => n3);
   U53 : HS65_LH_IVX9 port map( A => halt_i, Z => n52);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity exe_mem is

   port( clk, rst_n, halt_i : in std_logic;  EXE_MEM_i : in std_logic_vector 
         (71 downto 0);  EXE_MEM_o : out std_logic_vector (71 downto 0));

end exe_mem;

architecture SYN_Behavioral of exe_mem is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPSQX9
      port( D, CP, SN : in std_logic;  Q : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal EXE_MEM_o_ALU_RES_31_port, EXE_MEM_o_ALU_RES_30_port, 
      EXE_MEM_o_ALU_RES_29_port, EXE_MEM_o_ALU_RES_28_port, 
      EXE_MEM_o_ALU_RES_27_port, EXE_MEM_o_ALU_RES_26_port, 
      EXE_MEM_o_ALU_RES_25_port, EXE_MEM_o_ALU_RES_24_port, 
      EXE_MEM_o_ALU_RES_23_port, EXE_MEM_o_ALU_RES_22_port, 
      EXE_MEM_o_ALU_RES_21_port, EXE_MEM_o_ALU_RES_20_port, 
      EXE_MEM_o_ALU_RES_19_port, EXE_MEM_o_ALU_RES_18_port, 
      EXE_MEM_o_ALU_RES_17_port, EXE_MEM_o_ALU_RES_16_port, 
      EXE_MEM_o_ALU_RES_15_port, EXE_MEM_o_ALU_RES_14_port, 
      EXE_MEM_o_ALU_RES_13_port, EXE_MEM_o_ALU_RES_12_port, 
      EXE_MEM_o_ALU_RES_11_port, EXE_MEM_o_ALU_RES_10_port, 
      EXE_MEM_o_ALU_RES_9_port, EXE_MEM_o_ALU_RES_8_port, 
      EXE_MEM_o_ALU_RES_7_port, EXE_MEM_o_ALU_RES_6_port, 
      EXE_MEM_o_ALU_RES_5_port, EXE_MEM_o_ALU_RES_4_port, 
      EXE_MEM_o_ALU_RES_3_port, EXE_MEM_o_ALU_RES_2_port, 
      EXE_MEM_o_ALU_RES_1_port, EXE_MEM_o_ALU_RES_0_port, 
      EXE_MEM_o_DMEM_DATA_31_port, EXE_MEM_o_DMEM_DATA_30_port, 
      EXE_MEM_o_DMEM_DATA_29_port, EXE_MEM_o_DMEM_DATA_28_port, 
      EXE_MEM_o_DMEM_DATA_27_port, EXE_MEM_o_DMEM_DATA_26_port, 
      EXE_MEM_o_DMEM_DATA_25_port, EXE_MEM_o_DMEM_DATA_24_port, 
      EXE_MEM_o_DMEM_DATA_23_port, EXE_MEM_o_DMEM_DATA_22_port, 
      EXE_MEM_o_DMEM_DATA_21_port, EXE_MEM_o_DMEM_DATA_20_port, 
      EXE_MEM_o_DMEM_DATA_19_port, EXE_MEM_o_DMEM_DATA_18_port, 
      EXE_MEM_o_DMEM_DATA_17_port, EXE_MEM_o_DMEM_DATA_16_port, 
      EXE_MEM_o_DMEM_DATA_15_port, EXE_MEM_o_DMEM_DATA_14_port, 
      EXE_MEM_o_DMEM_DATA_13_port, EXE_MEM_o_DMEM_DATA_12_port, 
      EXE_MEM_o_DMEM_DATA_11_port, EXE_MEM_o_DMEM_DATA_10_port, 
      EXE_MEM_o_DMEM_DATA_9_port, EXE_MEM_o_DMEM_DATA_8_port, 
      EXE_MEM_o_DMEM_DATA_7_port, EXE_MEM_o_DMEM_DATA_6_port, 
      EXE_MEM_o_DMEM_DATA_5_port, EXE_MEM_o_DMEM_DATA_4_port, 
      EXE_MEM_o_DMEM_DATA_3_port, EXE_MEM_o_DMEM_DATA_2_port, 
      EXE_MEM_o_DMEM_DATA_1_port, EXE_MEM_o_DMEM_DATA_0_port, 
      EXE_MEM_o_WRITE_REG_4_port, EXE_MEM_o_WRITE_REG_3_port, 
      EXE_MEM_o_WRITE_REG_2_port, EXE_MEM_o_WRITE_REG_1_port, 
      EXE_MEM_o_WRITE_REG_0_port, EXE_MEM_o_MEMTOREG_port, 
      EXE_MEM_o_REGWRITE_port, EXE_MEM_o_MEMWEN_N_port, n2, n3, n4, n5, n6, n7,
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n1, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89 : std_logic;

begin
   EXE_MEM_o <= ( EXE_MEM_o_ALU_RES_31_port, EXE_MEM_o_ALU_RES_30_port, 
      EXE_MEM_o_ALU_RES_29_port, EXE_MEM_o_ALU_RES_28_port, 
      EXE_MEM_o_ALU_RES_27_port, EXE_MEM_o_ALU_RES_26_port, 
      EXE_MEM_o_ALU_RES_25_port, EXE_MEM_o_ALU_RES_24_port, 
      EXE_MEM_o_ALU_RES_23_port, EXE_MEM_o_ALU_RES_22_port, 
      EXE_MEM_o_ALU_RES_21_port, EXE_MEM_o_ALU_RES_20_port, 
      EXE_MEM_o_ALU_RES_19_port, EXE_MEM_o_ALU_RES_18_port, 
      EXE_MEM_o_ALU_RES_17_port, EXE_MEM_o_ALU_RES_16_port, 
      EXE_MEM_o_ALU_RES_15_port, EXE_MEM_o_ALU_RES_14_port, 
      EXE_MEM_o_ALU_RES_13_port, EXE_MEM_o_ALU_RES_12_port, 
      EXE_MEM_o_ALU_RES_11_port, EXE_MEM_o_ALU_RES_10_port, 
      EXE_MEM_o_ALU_RES_9_port, EXE_MEM_o_ALU_RES_8_port, 
      EXE_MEM_o_ALU_RES_7_port, EXE_MEM_o_ALU_RES_6_port, 
      EXE_MEM_o_ALU_RES_5_port, EXE_MEM_o_ALU_RES_4_port, 
      EXE_MEM_o_ALU_RES_3_port, EXE_MEM_o_ALU_RES_2_port, 
      EXE_MEM_o_ALU_RES_1_port, EXE_MEM_o_ALU_RES_0_port, 
      EXE_MEM_o_DMEM_DATA_31_port, EXE_MEM_o_DMEM_DATA_30_port, 
      EXE_MEM_o_DMEM_DATA_29_port, EXE_MEM_o_DMEM_DATA_28_port, 
      EXE_MEM_o_DMEM_DATA_27_port, EXE_MEM_o_DMEM_DATA_26_port, 
      EXE_MEM_o_DMEM_DATA_25_port, EXE_MEM_o_DMEM_DATA_24_port, 
      EXE_MEM_o_DMEM_DATA_23_port, EXE_MEM_o_DMEM_DATA_22_port, 
      EXE_MEM_o_DMEM_DATA_21_port, EXE_MEM_o_DMEM_DATA_20_port, 
      EXE_MEM_o_DMEM_DATA_19_port, EXE_MEM_o_DMEM_DATA_18_port, 
      EXE_MEM_o_DMEM_DATA_17_port, EXE_MEM_o_DMEM_DATA_16_port, 
      EXE_MEM_o_DMEM_DATA_15_port, EXE_MEM_o_DMEM_DATA_14_port, 
      EXE_MEM_o_DMEM_DATA_13_port, EXE_MEM_o_DMEM_DATA_12_port, 
      EXE_MEM_o_DMEM_DATA_11_port, EXE_MEM_o_DMEM_DATA_10_port, 
      EXE_MEM_o_DMEM_DATA_9_port, EXE_MEM_o_DMEM_DATA_8_port, 
      EXE_MEM_o_DMEM_DATA_7_port, EXE_MEM_o_DMEM_DATA_6_port, 
      EXE_MEM_o_DMEM_DATA_5_port, EXE_MEM_o_DMEM_DATA_4_port, 
      EXE_MEM_o_DMEM_DATA_3_port, EXE_MEM_o_DMEM_DATA_2_port, 
      EXE_MEM_o_DMEM_DATA_1_port, EXE_MEM_o_DMEM_DATA_0_port, 
      EXE_MEM_o_WRITE_REG_4_port, EXE_MEM_o_WRITE_REG_3_port, 
      EXE_MEM_o_WRITE_REG_2_port, EXE_MEM_o_WRITE_REG_1_port, 
      EXE_MEM_o_WRITE_REG_0_port, EXE_MEM_o_MEMTOREG_port, 
      EXE_MEM_o_REGWRITE_port, EXE_MEM_o_MEMWEN_N_port );
   
   exe_mem_c_reg_ALU_RES_31_inst : HS65_LH_DFPRQX9 port map( D => n73, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_31_port);
   exe_mem_c_reg_ALU_RES_30_inst : HS65_LH_DFPRQX9 port map( D => n72, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_30_port);
   exe_mem_c_reg_ALU_RES_29_inst : HS65_LH_DFPRQX9 port map( D => n71, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_29_port);
   exe_mem_c_reg_ALU_RES_28_inst : HS65_LH_DFPRQX9 port map( D => n70, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_28_port);
   exe_mem_c_reg_ALU_RES_27_inst : HS65_LH_DFPRQX9 port map( D => n69, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_27_port);
   exe_mem_c_reg_ALU_RES_26_inst : HS65_LH_DFPRQX9 port map( D => n68, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_26_port);
   exe_mem_c_reg_ALU_RES_25_inst : HS65_LH_DFPRQX9 port map( D => n67, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_25_port);
   exe_mem_c_reg_ALU_RES_24_inst : HS65_LH_DFPRQX9 port map( D => n66, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_24_port);
   exe_mem_c_reg_ALU_RES_23_inst : HS65_LH_DFPRQX9 port map( D => n65, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_23_port);
   exe_mem_c_reg_ALU_RES_22_inst : HS65_LH_DFPRQX9 port map( D => n64, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_22_port);
   exe_mem_c_reg_ALU_RES_21_inst : HS65_LH_DFPRQX9 port map( D => n63, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_21_port);
   exe_mem_c_reg_ALU_RES_20_inst : HS65_LH_DFPRQX9 port map( D => n62, CP => 
                           clk, RN => n83, Q => EXE_MEM_o_ALU_RES_20_port);
   exe_mem_c_reg_ALU_RES_19_inst : HS65_LH_DFPRQX9 port map( D => n61, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_19_port);
   exe_mem_c_reg_ALU_RES_18_inst : HS65_LH_DFPRQX9 port map( D => n60, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_18_port);
   exe_mem_c_reg_ALU_RES_17_inst : HS65_LH_DFPRQX9 port map( D => n59, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_17_port);
   exe_mem_c_reg_ALU_RES_16_inst : HS65_LH_DFPRQX9 port map( D => n58, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_16_port);
   exe_mem_c_reg_ALU_RES_15_inst : HS65_LH_DFPRQX9 port map( D => n57, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_15_port);
   exe_mem_c_reg_ALU_RES_14_inst : HS65_LH_DFPRQX9 port map( D => n56, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_14_port);
   exe_mem_c_reg_ALU_RES_13_inst : HS65_LH_DFPRQX9 port map( D => n55, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_13_port);
   exe_mem_c_reg_ALU_RES_12_inst : HS65_LH_DFPRQX9 port map( D => n54, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_12_port);
   exe_mem_c_reg_ALU_RES_11_inst : HS65_LH_DFPRQX9 port map( D => n53, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_11_port);
   exe_mem_c_reg_ALU_RES_10_inst : HS65_LH_DFPRQX9 port map( D => n52, CP => 
                           clk, RN => n84, Q => EXE_MEM_o_ALU_RES_10_port);
   exe_mem_c_reg_ALU_RES_9_inst : HS65_LH_DFPRQX9 port map( D => n51, CP => clk
                           , RN => n84, Q => EXE_MEM_o_ALU_RES_9_port);
   exe_mem_c_reg_ALU_RES_8_inst : HS65_LH_DFPRQX9 port map( D => n50, CP => clk
                           , RN => n84, Q => EXE_MEM_o_ALU_RES_8_port);
   exe_mem_c_reg_ALU_RES_7_inst : HS65_LH_DFPRQX9 port map( D => n49, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_7_port);
   exe_mem_c_reg_ALU_RES_6_inst : HS65_LH_DFPRQX9 port map( D => n48, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_6_port);
   exe_mem_c_reg_ALU_RES_5_inst : HS65_LH_DFPRQX9 port map( D => n47, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_5_port);
   exe_mem_c_reg_ALU_RES_4_inst : HS65_LH_DFPRQX9 port map( D => n46, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_4_port);
   exe_mem_c_reg_ALU_RES_3_inst : HS65_LH_DFPRQX9 port map( D => n45, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_3_port);
   exe_mem_c_reg_ALU_RES_2_inst : HS65_LH_DFPRQX9 port map( D => n44, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_2_port);
   exe_mem_c_reg_ALU_RES_1_inst : HS65_LH_DFPRQX9 port map( D => n43, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_1_port);
   exe_mem_c_reg_ALU_RES_0_inst : HS65_LH_DFPRQX9 port map( D => n42, CP => clk
                           , RN => n85, Q => EXE_MEM_o_ALU_RES_0_port);
   exe_mem_c_reg_DMEM_DATA_31_inst : HS65_LH_DFPRQX9 port map( D => n41, CP => 
                           clk, RN => n85, Q => EXE_MEM_o_DMEM_DATA_31_port);
   exe_mem_c_reg_DMEM_DATA_30_inst : HS65_LH_DFPRQX9 port map( D => n40, CP => 
                           clk, RN => n85, Q => EXE_MEM_o_DMEM_DATA_30_port);
   exe_mem_c_reg_DMEM_DATA_29_inst : HS65_LH_DFPRQX9 port map( D => n39, CP => 
                           clk, RN => n85, Q => EXE_MEM_o_DMEM_DATA_29_port);
   exe_mem_c_reg_DMEM_DATA_28_inst : HS65_LH_DFPRQX9 port map( D => n38, CP => 
                           clk, RN => n85, Q => EXE_MEM_o_DMEM_DATA_28_port);
   exe_mem_c_reg_DMEM_DATA_27_inst : HS65_LH_DFPRQX9 port map( D => n37, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_27_port);
   exe_mem_c_reg_DMEM_DATA_26_inst : HS65_LH_DFPRQX9 port map( D => n36, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_26_port);
   exe_mem_c_reg_DMEM_DATA_25_inst : HS65_LH_DFPRQX9 port map( D => n35, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_25_port);
   exe_mem_c_reg_DMEM_DATA_24_inst : HS65_LH_DFPRQX9 port map( D => n34, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_24_port);
   exe_mem_c_reg_DMEM_DATA_23_inst : HS65_LH_DFPRQX9 port map( D => n33, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_23_port);
   exe_mem_c_reg_DMEM_DATA_22_inst : HS65_LH_DFPRQX9 port map( D => n32, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_22_port);
   exe_mem_c_reg_DMEM_DATA_21_inst : HS65_LH_DFPRQX9 port map( D => n31, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_21_port);
   exe_mem_c_reg_DMEM_DATA_20_inst : HS65_LH_DFPRQX9 port map( D => n30, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_20_port);
   exe_mem_c_reg_DMEM_DATA_19_inst : HS65_LH_DFPRQX9 port map( D => n29, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_19_port);
   exe_mem_c_reg_DMEM_DATA_18_inst : HS65_LH_DFPRQX9 port map( D => n28, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_18_port);
   exe_mem_c_reg_DMEM_DATA_17_inst : HS65_LH_DFPRQX9 port map( D => n27, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_17_port);
   exe_mem_c_reg_DMEM_DATA_16_inst : HS65_LH_DFPRQX9 port map( D => n26, CP => 
                           clk, RN => n86, Q => EXE_MEM_o_DMEM_DATA_16_port);
   exe_mem_c_reg_DMEM_DATA_15_inst : HS65_LH_DFPRQX9 port map( D => n25, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_15_port);
   exe_mem_c_reg_DMEM_DATA_14_inst : HS65_LH_DFPRQX9 port map( D => n24, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_14_port);
   exe_mem_c_reg_DMEM_DATA_13_inst : HS65_LH_DFPRQX9 port map( D => n23, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_13_port);
   exe_mem_c_reg_DMEM_DATA_12_inst : HS65_LH_DFPRQX9 port map( D => n22, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_12_port);
   exe_mem_c_reg_DMEM_DATA_11_inst : HS65_LH_DFPRQX9 port map( D => n21, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_11_port);
   exe_mem_c_reg_DMEM_DATA_10_inst : HS65_LH_DFPRQX9 port map( D => n20, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_10_port);
   exe_mem_c_reg_DMEM_DATA_9_inst : HS65_LH_DFPRQX9 port map( D => n19, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_9_port);
   exe_mem_c_reg_DMEM_DATA_8_inst : HS65_LH_DFPRQX9 port map( D => n18, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_8_port);
   exe_mem_c_reg_DMEM_DATA_7_inst : HS65_LH_DFPRQX9 port map( D => n17, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_7_port);
   exe_mem_c_reg_DMEM_DATA_6_inst : HS65_LH_DFPRQX9 port map( D => n16, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_6_port);
   exe_mem_c_reg_DMEM_DATA_5_inst : HS65_LH_DFPRQX9 port map( D => n15, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_5_port);
   exe_mem_c_reg_DMEM_DATA_4_inst : HS65_LH_DFPRQX9 port map( D => n14, CP => 
                           clk, RN => n87, Q => EXE_MEM_o_DMEM_DATA_4_port);
   exe_mem_c_reg_DMEM_DATA_3_inst : HS65_LH_DFPRQX9 port map( D => n13, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_DMEM_DATA_3_port);
   exe_mem_c_reg_DMEM_DATA_2_inst : HS65_LH_DFPRQX9 port map( D => n12, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_DMEM_DATA_2_port);
   exe_mem_c_reg_DMEM_DATA_1_inst : HS65_LH_DFPRQX9 port map( D => n11, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_DMEM_DATA_1_port);
   exe_mem_c_reg_DMEM_DATA_0_inst : HS65_LH_DFPRQX9 port map( D => n10, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_DMEM_DATA_0_port);
   exe_mem_c_reg_WRITE_REG_4_inst : HS65_LH_DFPRQX9 port map( D => n9, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_WRITE_REG_4_port);
   exe_mem_c_reg_WRITE_REG_3_inst : HS65_LH_DFPRQX9 port map( D => n8, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_WRITE_REG_3_port);
   exe_mem_c_reg_WRITE_REG_2_inst : HS65_LH_DFPRQX9 port map( D => n7, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_WRITE_REG_2_port);
   exe_mem_c_reg_WRITE_REG_1_inst : HS65_LH_DFPRQX9 port map( D => n6, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_WRITE_REG_1_port);
   exe_mem_c_reg_WRITE_REG_0_inst : HS65_LH_DFPRQX9 port map( D => n5, CP => 
                           clk, RN => n88, Q => EXE_MEM_o_WRITE_REG_0_port);
   exe_mem_c_reg_MEMTOREG_inst : HS65_LH_DFPRQX9 port map( D => n4, CP => clk, 
                           RN => n88, Q => EXE_MEM_o_MEMTOREG_port);
   exe_mem_c_reg_REGWRITE_inst : HS65_LH_DFPRQX9 port map( D => n3, CP => clk, 
                           RN => n88, Q => EXE_MEM_o_REGWRITE_port);
   exe_mem_c_reg_MEMWEN_N_inst : HS65_LH_DFPSQX9 port map( D => n2, CP => clk, 
                           SN => n88, Q => EXE_MEM_o_MEMWEN_N_port);
   U2 : HS65_LH_BFX9 port map( A => n82, Z => n87);
   U3 : HS65_LH_BFX9 port map( A => n82, Z => n86);
   U4 : HS65_LH_BFX9 port map( A => n81, Z => n85);
   U5 : HS65_LH_BFX9 port map( A => n81, Z => n84);
   U6 : HS65_LH_BFX9 port map( A => n81, Z => n83);
   U7 : HS65_LH_BFX9 port map( A => n82, Z => n88);
   U8 : HS65_LH_BFX9 port map( A => rst_n, Z => n82);
   U9 : HS65_LH_BFX9 port map( A => rst_n, Z => n81);
   U10 : HS65_LH_BFX9 port map( A => n1, Z => n75);
   U11 : HS65_LH_BFX9 port map( A => n1, Z => n76);
   U12 : HS65_LH_BFX9 port map( A => n1, Z => n77);
   U13 : HS65_LH_BFX9 port map( A => n74, Z => n78);
   U14 : HS65_LH_BFX9 port map( A => n74, Z => n79);
   U15 : HS65_LH_BFX9 port map( A => n74, Z => n80);
   U16 : HS65_LH_BFX9 port map( A => n89, Z => n1);
   U17 : HS65_LH_BFX9 port map( A => n89, Z => n74);
   U18 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_25_port, B => halt_i, 
                           C => EXE_MEM_i(65), D => n80, Z => n67);
   U19 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_26_port, B => halt_i, 
                           C => EXE_MEM_i(66), D => n80, Z => n68);
   U20 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_27_port, B => halt_i, 
                           C => EXE_MEM_i(67), D => n80, Z => n69);
   U21 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_29_port, B => halt_i, 
                           C => EXE_MEM_i(69), D => n80, Z => n71);
   U22 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_30_port, B => halt_i, 
                           C => EXE_MEM_i(70), D => n80, Z => n72);
   U23 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_28_port, B => halt_i, 
                           C => EXE_MEM_i(68), D => n80, Z => n70);
   U24 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_31_port, B => halt_i, 
                           C => EXE_MEM_i(71), D => n80, Z => n73);
   U25 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_21_port, B => halt_i, 
                           C => EXE_MEM_i(61), D => n80, Z => n63);
   U26 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_22_port, B => halt_i, 
                           C => EXE_MEM_i(62), D => n80, Z => n64);
   U27 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_23_port, B => halt_i, 
                           C => EXE_MEM_i(63), D => n80, Z => n65);
   U28 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_24_port, B => halt_i, 
                           C => EXE_MEM_i(64), D => n80, Z => n66);
   U29 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_17_port, B => halt_i, 
                           C => EXE_MEM_i(57), D => n79, Z => n59);
   U30 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_18_port, B => halt_i, 
                           C => EXE_MEM_i(58), D => n79, Z => n60);
   U31 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_19_port, B => halt_i, 
                           C => EXE_MEM_i(59), D => n79, Z => n61);
   U32 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_20_port, B => halt_i, 
                           C => EXE_MEM_i(60), D => n80, Z => n62);
   U33 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_0_port, B => halt_i, C
                           => EXE_MEM_i(40), D => n78, Z => n42);
   U34 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_16_port, B => halt_i, 
                           C => EXE_MEM_i(56), D => n79, Z => n58);
   U35 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_9_port, B => halt_i, C
                           => EXE_MEM_i(49), D => n79, Z => n51);
   U36 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_10_port, B => halt_i, 
                           C => EXE_MEM_i(50), D => n79, Z => n52);
   U37 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_11_port, B => halt_i, 
                           C => EXE_MEM_i(51), D => n79, Z => n53);
   U38 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_12_port, B => halt_i, 
                           C => EXE_MEM_i(52), D => n79, Z => n54);
   U39 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_13_port, B => halt_i, 
                           C => EXE_MEM_i(53), D => n79, Z => n55);
   U40 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_14_port, B => halt_i, 
                           C => EXE_MEM_i(54), D => n79, Z => n56);
   U41 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_15_port, B => halt_i, 
                           C => EXE_MEM_i(55), D => n79, Z => n57);
   U42 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_1_port, B => halt_i, C
                           => EXE_MEM_i(41), D => n78, Z => n43);
   U43 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_4_port, B => halt_i, C
                           => EXE_MEM_i(44), D => n78, Z => n46);
   U44 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_5_port, B => halt_i, C
                           => EXE_MEM_i(45), D => n78, Z => n47);
   U45 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_6_port, B => halt_i, C
                           => EXE_MEM_i(46), D => n78, Z => n48);
   U46 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_7_port, B => halt_i, C
                           => EXE_MEM_i(47), D => n78, Z => n49);
   U47 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_8_port, B => halt_i, C
                           => EXE_MEM_i(48), D => n79, Z => n50);
   U48 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_2_port, B => halt_i, C
                           => EXE_MEM_i(42), D => n78, Z => n44);
   U49 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_ALU_RES_3_port, B => halt_i, C
                           => EXE_MEM_i(43), D => n78, Z => n45);
   U50 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_9_port, B => halt_i,
                           C => EXE_MEM_i(17), D => n76, Z => n19);
   U51 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_12_port, B => halt_i
                           , C => EXE_MEM_i(20), D => n76, Z => n22);
   U52 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_13_port, B => halt_i
                           , C => EXE_MEM_i(21), D => n76, Z => n23);
   U53 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_14_port, B => halt_i
                           , C => EXE_MEM_i(22), D => n76, Z => n24);
   U54 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_15_port, B => halt_i
                           , C => EXE_MEM_i(23), D => n76, Z => n25);
   U55 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_16_port, B => halt_i
                           , C => EXE_MEM_i(24), D => n77, Z => n26);
   U56 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_17_port, B => halt_i
                           , C => EXE_MEM_i(25), D => n77, Z => n27);
   U57 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_18_port, B => halt_i
                           , C => EXE_MEM_i(26), D => n77, Z => n28);
   U58 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_19_port, B => halt_i
                           , C => EXE_MEM_i(27), D => n77, Z => n29);
   U59 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_20_port, B => halt_i
                           , C => EXE_MEM_i(28), D => n77, Z => n30);
   U60 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_21_port, B => halt_i
                           , C => EXE_MEM_i(29), D => n77, Z => n31);
   U61 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_22_port, B => halt_i
                           , C => EXE_MEM_i(30), D => n77, Z => n32);
   U62 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_23_port, B => halt_i
                           , C => EXE_MEM_i(31), D => n77, Z => n33);
   U63 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_24_port, B => halt_i
                           , C => EXE_MEM_i(32), D => n77, Z => n34);
   U64 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_25_port, B => halt_i
                           , C => EXE_MEM_i(33), D => n77, Z => n35);
   U65 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_26_port, B => halt_i
                           , C => EXE_MEM_i(34), D => n77, Z => n36);
   U66 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_27_port, B => halt_i
                           , C => EXE_MEM_i(35), D => n77, Z => n37);
   U67 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_28_port, B => halt_i
                           , C => EXE_MEM_i(36), D => n78, Z => n38);
   U68 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_29_port, B => halt_i
                           , C => EXE_MEM_i(37), D => n78, Z => n39);
   U69 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_30_port, B => halt_i
                           , C => EXE_MEM_i(38), D => n78, Z => n40);
   U70 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_31_port, B => halt_i
                           , C => EXE_MEM_i(39), D => n78, Z => n41);
   U71 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_0_port, B => halt_i,
                           C => EXE_MEM_i(8), D => n75, Z => n10);
   U72 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_1_port, B => halt_i,
                           C => EXE_MEM_i(9), D => n75, Z => n11);
   U73 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_2_port, B => halt_i,
                           C => EXE_MEM_i(10), D => n75, Z => n12);
   U74 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_3_port, B => halt_i,
                           C => EXE_MEM_i(11), D => n75, Z => n13);
   U75 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_4_port, B => halt_i,
                           C => EXE_MEM_i(12), D => n76, Z => n14);
   U76 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_5_port, B => halt_i,
                           C => EXE_MEM_i(13), D => n76, Z => n15);
   U77 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_6_port, B => halt_i,
                           C => EXE_MEM_i(14), D => n76, Z => n16);
   U78 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_7_port, B => halt_i,
                           C => EXE_MEM_i(15), D => n76, Z => n17);
   U79 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_8_port, B => halt_i,
                           C => EXE_MEM_i(16), D => n76, Z => n18);
   U80 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_10_port, B => halt_i
                           , C => EXE_MEM_i(18), D => n76, Z => n20);
   U81 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_DMEM_DATA_11_port, B => halt_i
                           , C => EXE_MEM_i(19), D => n76, Z => n21);
   U82 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_WRITE_REG_0_port, B => halt_i,
                           C => EXE_MEM_i(3), D => n75, Z => n5);
   U83 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_WRITE_REG_1_port, B => halt_i,
                           C => EXE_MEM_i(4), D => n75, Z => n6);
   U84 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_WRITE_REG_2_port, B => halt_i,
                           C => EXE_MEM_i(5), D => n75, Z => n7);
   U85 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_WRITE_REG_3_port, B => halt_i,
                           C => EXE_MEM_i(6), D => n75, Z => n8);
   U86 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_WRITE_REG_4_port, B => halt_i,
                           C => EXE_MEM_i(7), D => n75, Z => n9);
   U87 : HS65_LH_AO22X9 port map( A => halt_i, B => EXE_MEM_o_MEMWEN_N_port, C 
                           => EXE_MEM_i(0), D => n75, Z => n2);
   U88 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_REGWRITE_port, B => halt_i, C 
                           => EXE_MEM_i(1), D => n75, Z => n3);
   U89 : HS65_LH_AO22X9 port map( A => EXE_MEM_o_MEMTOREG_port, B => halt_i, C 
                           => EXE_MEM_i(2), D => n75, Z => n4);
   U90 : HS65_LH_IVX9 port map( A => halt_i, Z => n89);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity forwarding_unit is

   port( forwarding_unit_i : in std_logic_vector (31 downto 0);  
         forwarding_unit_o : out std_logic_vector (5 downto 0));

end forwarding_unit;

architecture SYN_behavioral of forwarding_unit is

   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OR3X9
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OA31X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   signal forwarding_unit_o_FORWARD_A_1_port, 
      forwarding_unit_o_FORWARD_A_0_port, forwarding_unit_o_FORWARD_B_1_port, 
      forwarding_unit_o_FORWARD_B_0_port, 
      forwarding_unit_o_REGFILE_FORWARD_A_port, 
      forwarding_unit_o_REGFILE_FORWARD_B_port, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n1 : std_logic;

begin
   forwarding_unit_o <= ( forwarding_unit_o_FORWARD_A_1_port, 
      forwarding_unit_o_FORWARD_A_0_port, forwarding_unit_o_FORWARD_B_1_port, 
      forwarding_unit_o_FORWARD_B_0_port, 
      forwarding_unit_o_REGFILE_FORWARD_A_port, 
      forwarding_unit_o_REGFILE_FORWARD_B_port );
   
   U2 : HS65_LH_NOR4ABX2 port map( A => n58, B => n59, C => n60, D => n61, Z =>
                           forwarding_unit_o_FORWARD_A_1_port);
   U3 : HS65_LH_NOR4ABX2 port map( A => n45, B => n46, C => n47, D => n48, Z =>
                           forwarding_unit_o_FORWARD_B_1_port);
   U4 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(7), B => 
                           forwarding_unit_i(27), Z => n60);
   U5 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(10), B => 
                           forwarding_unit_i(30), Z => n59);
   U6 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(8), B => 
                           forwarding_unit_i(28), Z => n58);
   U7 : HS65_LH_NOR4ABX2 port map( A => n51, B => n52, C => n53, D => n54, Z =>
                           forwarding_unit_o_FORWARD_A_0_port);
   U8 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(5), B => 
                           forwarding_unit_i(30), Z => n51);
   U9 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(2), B => 
                           forwarding_unit_i(27), Z => n54);
   U10 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(3), B => 
                           forwarding_unit_i(28), Z => n52);
   U11 : HS65_LH_OA31X9 port map( A => n57, B => forwarding_unit_i(3), C => 
                           forwarding_unit_i(2), D => forwarding_unit_i(0), Z 
                           => n27);
   U12 : HS65_LH_OR3X9 port map( A => forwarding_unit_i(6), B => 
                           forwarding_unit_i(5), C => forwarding_unit_i(4), Z 
                           => n57);
   U13 : HS65_LH_NAND4ABX3 port map( A => n62, B => n63, C => 
                           forwarding_unit_i(1), D => n1, Z => n61);
   U14 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(9), B => 
                           forwarding_unit_i(29), Z => n63);
   U15 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(11), B => 
                           forwarding_unit_i(31), Z => n62);
   U16 : HS65_LH_NAND4ABX3 port map( A => n55, B => 
                           forwarding_unit_o_FORWARD_A_1_port, C => n56, D => 
                           n27, Z => n53);
   U17 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(4), B => 
                           forwarding_unit_i(29), Z => n56);
   U18 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(6), B => 
                           forwarding_unit_i(31), Z => n55);
   U19 : HS65_LH_IVX9 port map( A => n64, Z => n1);
   U20 : HS65_LH_NOR3AX2 port map( A => n65, B => forwarding_unit_i(7), C => 
                           forwarding_unit_i(8), Z => n64);
   U21 : HS65_LH_NOR3X4 port map( A => forwarding_unit_i(9), B => 
                           forwarding_unit_i(11), C => forwarding_unit_i(10), Z
                           => n65);
   U22 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(10), B => 
                           forwarding_unit_i(25), Z => n47);
   U23 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(7), B => 
                           forwarding_unit_i(22), Z => n46);
   U24 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(8), B => 
                           forwarding_unit_i(23), Z => n45);
   U25 : HS65_LH_NOR4ABX2 port map( A => n39, B => n40, C => n41, D => n42, Z 
                           => forwarding_unit_o_FORWARD_B_0_port);
   U26 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(5), B => 
                           forwarding_unit_i(25), Z => n39);
   U27 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(2), B => 
                           forwarding_unit_i(22), Z => n42);
   U28 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(3), B => 
                           forwarding_unit_i(23), Z => n40);
   U29 : HS65_LH_NAND4ABX3 port map( A => n49, B => n50, C => 
                           forwarding_unit_i(1), D => n1, Z => n48);
   U30 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(9), B => 
                           forwarding_unit_i(24), Z => n50);
   U31 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(11), B => 
                           forwarding_unit_i(26), Z => n49);
   U32 : HS65_LH_NAND4ABX3 port map( A => n43, B => 
                           forwarding_unit_o_FORWARD_B_1_port, C => n44, D => 
                           n27, Z => n41);
   U33 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(4), B => 
                           forwarding_unit_i(24), Z => n44);
   U34 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(6), B => 
                           forwarding_unit_i(26), Z => n43);
   U35 : HS65_LH_NOR4ABX2 port map( A => n33, B => n27, C => n34, D => n35, Z 
                           => forwarding_unit_o_REGFILE_FORWARD_A_port);
   U36 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(6), B => 
                           forwarding_unit_i(21), Z => n35);
   U37 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(19), B => 
                           forwarding_unit_i(4), Z => n33);
   U38 : HS65_LH_NOR4ABX2 port map( A => n26, B => n27, C => n28, D => n29, Z 
                           => forwarding_unit_o_REGFILE_FORWARD_B_port);
   U39 : HS65_LHS_XOR2X6 port map( A => forwarding_unit_i(6), B => 
                           forwarding_unit_i(16), Z => n29);
   U40 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(15), B => 
                           forwarding_unit_i(5), Z => n26);
   U41 : HS65_LH_NAND3X5 port map( A => n30, B => n31, C => n32, Z => n28);
   U42 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(13), B => 
                           forwarding_unit_i(3), Z => n32);
   U43 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(14), B => 
                           forwarding_unit_i(4), Z => n31);
   U44 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(12), B => 
                           forwarding_unit_i(2), Z => n30);
   U45 : HS65_LH_NAND3X5 port map( A => n36, B => n37, C => n38, Z => n34);
   U46 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(18), B => 
                           forwarding_unit_i(3), Z => n38);
   U47 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(20), B => 
                           forwarding_unit_i(5), Z => n36);
   U48 : HS65_LHS_XNOR2X6 port map( A => forwarding_unit_i(17), B => 
                           forwarding_unit_i(2), Z => n37);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity exe_top is

   port( clk, rst_n : in std_logic;  exe_top_i : in std_logic_vector (134 
         downto 0);  exe_top_o : out std_logic_vector (81 downto 0));

end exe_top;

architecture SYN_Behavioral of exe_top is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO212X4
      port( A, B, C, D, E : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2AX3
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component exe_top_DW01_add_0
      port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (11 downto 0);  CO : out std_logic);
   end component;
   
   component alu_ctrl
      port( alu_ctrl_i : in std_logic_vector (9 downto 0);  alu_ctrl_o : out 
            std_logic_vector (6 downto 0));
   end component;
   
   component alu
      port( clk, rst_n : in std_logic;  alu_i : in std_logic_vector (73 downto 
            0);  alu_o : out std_logic_vector (32 downto 0));
   end component;
   
   signal op_aluCtrl_alu_4_port, op_aluCtrl_alu_3_port, op_aluCtrl_alu_2_port, 
      op_aluCtrl_alu_1_port, op_aluCtrl_alu_0_port, src_a_31_port, 
      src_a_30_port, src_a_29_port, src_a_28_port, src_a_27_port, src_a_26_port
      , src_a_25_port, src_a_24_port, src_a_23_port, src_a_22_port, 
      src_a_21_port, src_a_20_port, src_a_19_port, src_a_18_port, src_a_17_port
      , src_a_16_port, src_a_15_port, src_a_14_port, src_a_13_port, 
      src_a_12_port, src_a_11_port, src_a_10_port, src_a_9_port, src_a_8_port, 
      src_a_7_port, src_a_6_port, src_a_5_port, src_a_4_port, src_a_3_port, 
      src_a_2_port, src_a_1_port, src_a_0_port, src_b_31_port, src_b_30_port, 
      src_b_29_port, src_b_28_port, src_b_27_port, src_b_26_port, src_b_25_port
      , src_b_24_port, src_b_23_port, src_b_22_port, src_b_21_port, 
      src_b_20_port, src_b_19_port, src_b_18_port, src_b_17_port, src_b_16_port
      , src_b_15_port, src_b_14_port, src_b_13_port, src_b_12_port, 
      src_b_11_port, src_b_10_port, src_b_9_port, src_b_8_port, src_b_7_port, 
      src_b_6_port, src_b_5_port, src_b_4_port, src_b_3_port, src_b_2_port, 
      src_b_1_port, src_b_0_port, s_branch_src_1_port, s_branch_src_0_port, N22
      , N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, n3, n7, n8, n9, 
      n10, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n_1020 :
      std_logic;

begin
   
   n3 <= '0';
   alu_inst : alu port map( clk => clk, rst_n => n47, alu_i(73) => 
                           src_a_31_port, alu_i(72) => src_a_30_port, alu_i(71)
                           => src_a_29_port, alu_i(70) => src_a_28_port, 
                           alu_i(69) => src_a_27_port, alu_i(68) => 
                           src_a_26_port, alu_i(67) => src_a_25_port, alu_i(66)
                           => src_a_24_port, alu_i(65) => src_a_23_port, 
                           alu_i(64) => src_a_22_port, alu_i(63) => 
                           src_a_21_port, alu_i(62) => src_a_20_port, alu_i(61)
                           => src_a_19_port, alu_i(60) => src_a_18_port, 
                           alu_i(59) => src_a_17_port, alu_i(58) => 
                           src_a_16_port, alu_i(57) => src_a_15_port, alu_i(56)
                           => src_a_14_port, alu_i(55) => src_a_13_port, 
                           alu_i(54) => src_a_12_port, alu_i(53) => 
                           src_a_11_port, alu_i(52) => src_a_10_port, alu_i(51)
                           => src_a_9_port, alu_i(50) => src_a_8_port, 
                           alu_i(49) => src_a_7_port, alu_i(48) => src_a_6_port
                           , alu_i(47) => src_a_5_port, alu_i(46) => 
                           src_a_4_port, alu_i(45) => src_a_3_port, alu_i(44) 
                           => src_a_2_port, alu_i(43) => src_a_1_port, 
                           alu_i(42) => src_a_0_port, alu_i(41) => 
                           src_b_31_port, alu_i(40) => src_b_30_port, alu_i(39)
                           => src_b_29_port, alu_i(38) => src_b_28_port, 
                           alu_i(37) => src_b_27_port, alu_i(36) => 
                           src_b_26_port, alu_i(35) => src_b_25_port, alu_i(34)
                           => src_b_24_port, alu_i(33) => src_b_23_port, 
                           alu_i(32) => src_b_22_port, alu_i(31) => 
                           src_b_21_port, alu_i(30) => src_b_20_port, alu_i(29)
                           => src_b_19_port, alu_i(28) => src_b_18_port, 
                           alu_i(27) => src_b_17_port, alu_i(26) => 
                           src_b_16_port, alu_i(25) => src_b_15_port, alu_i(24)
                           => src_b_14_port, alu_i(23) => src_b_13_port, 
                           alu_i(22) => src_b_12_port, alu_i(21) => 
                           src_b_11_port, alu_i(20) => src_b_10_port, alu_i(19)
                           => src_b_9_port, alu_i(18) => src_b_8_port, 
                           alu_i(17) => src_b_7_port, alu_i(16) => src_b_6_port
                           , alu_i(15) => src_b_5_port, alu_i(14) => 
                           src_b_4_port, alu_i(13) => src_b_3_port, alu_i(12) 
                           => src_b_2_port, alu_i(11) => src_b_1_port, 
                           alu_i(10) => src_b_0_port, alu_i(9) => 
                           op_aluCtrl_alu_4_port, alu_i(8) => 
                           op_aluCtrl_alu_3_port, alu_i(7) => 
                           op_aluCtrl_alu_2_port, alu_i(6) => 
                           op_aluCtrl_alu_1_port, alu_i(5) => 
                           op_aluCtrl_alu_0_port, alu_i(4) => exe_top_i(134), 
                           alu_i(3) => exe_top_i(133), alu_i(2) => 
                           exe_top_i(132), alu_i(1) => exe_top_i(131), alu_i(0)
                           => exe_top_i(130), alu_o(32) => exe_top_o(81), 
                           alu_o(31) => exe_top_o(68), alu_o(30) => 
                           exe_top_o(67), alu_o(29) => exe_top_o(66), alu_o(28)
                           => exe_top_o(65), alu_o(27) => exe_top_o(64), 
                           alu_o(26) => exe_top_o(63), alu_o(25) => 
                           exe_top_o(62), alu_o(24) => exe_top_o(61), alu_o(23)
                           => exe_top_o(60), alu_o(22) => exe_top_o(59), 
                           alu_o(21) => exe_top_o(58), alu_o(20) => 
                           exe_top_o(57), alu_o(19) => exe_top_o(56), alu_o(18)
                           => exe_top_o(55), alu_o(17) => exe_top_o(54), 
                           alu_o(16) => exe_top_o(53), alu_o(15) => 
                           exe_top_o(52), alu_o(14) => exe_top_o(51), alu_o(13)
                           => exe_top_o(50), alu_o(12) => exe_top_o(49), 
                           alu_o(11) => exe_top_o(48), alu_o(10) => 
                           exe_top_o(47), alu_o(9) => exe_top_o(46), alu_o(8) 
                           => exe_top_o(45), alu_o(7) => exe_top_o(44), 
                           alu_o(6) => exe_top_o(43), alu_o(5) => exe_top_o(42)
                           , alu_o(4) => exe_top_o(41), alu_o(3) => 
                           exe_top_o(40), alu_o(2) => exe_top_o(39), alu_o(1) 
                           => exe_top_o(38), alu_o(0) => exe_top_o(37));
   alu_ctrl_inst : alu_ctrl port map( alu_ctrl_i(9) => exe_top_i(32), 
                           alu_ctrl_i(8) => exe_top_i(31), alu_ctrl_i(7) => 
                           exe_top_i(30), alu_ctrl_i(6) => exe_top_i(29), 
                           alu_ctrl_i(5) => exe_top_i(28), alu_ctrl_i(4) => 
                           exe_top_i(27), alu_ctrl_i(3) => exe_top_i(26), 
                           alu_ctrl_i(2) => exe_top_i(25), alu_ctrl_i(1) => 
                           exe_top_i(24), alu_ctrl_i(0) => exe_top_i(23), 
                           alu_ctrl_o(6) => op_aluCtrl_alu_4_port, 
                           alu_ctrl_o(5) => op_aluCtrl_alu_3_port, 
                           alu_ctrl_o(4) => op_aluCtrl_alu_2_port, 
                           alu_ctrl_o(3) => op_aluCtrl_alu_1_port, 
                           alu_ctrl_o(2) => op_aluCtrl_alu_0_port, 
                           alu_ctrl_o(1) => s_branch_src_1_port, alu_ctrl_o(0) 
                           => s_branch_src_0_port);
   add_53 : exe_top_DW01_add_0 port map( A(11) => exe_top_i(22), A(10) => 
                           exe_top_i(21), A(9) => exe_top_i(20), A(8) => 
                           exe_top_i(19), A(7) => exe_top_i(18), A(6) => 
                           exe_top_i(17), A(5) => exe_top_i(16), A(4) => 
                           exe_top_i(15), A(3) => exe_top_i(14), A(2) => 
                           exe_top_i(13), A(1) => exe_top_i(12), A(0) => 
                           exe_top_i(11), B(11) => exe_top_i(44), B(10) => 
                           exe_top_i(43), B(9) => exe_top_i(42), B(8) => 
                           exe_top_i(41), B(7) => exe_top_i(40), B(6) => 
                           exe_top_i(39), B(5) => exe_top_i(38), B(4) => 
                           exe_top_i(37), B(3) => exe_top_i(36), B(2) => 
                           exe_top_i(35), B(1) => exe_top_i(34), B(0) => 
                           exe_top_i(33), CI => n3, SUM(11) => N33, SUM(10) => 
                           N32, SUM(9) => N31, SUM(8) => N30, SUM(7) => N29, 
                           SUM(6) => N28, SUM(5) => N27, SUM(4) => N26, SUM(3) 
                           => N25, SUM(2) => N24, SUM(1) => N23, SUM(0) => N22,
                           CO => n_1020);
   U4 : HS65_LH_NOR2AX3 port map( A => exe_top_i(110), B => n38, Z => 
                           src_a_12_port);
   U5 : HS65_LH_NOR2AX3 port map( A => exe_top_i(111), B => n38, Z => 
                           src_a_13_port);
   U6 : HS65_LH_NOR2AX3 port map( A => exe_top_i(113), B => n38, Z => 
                           src_a_15_port);
   U7 : HS65_LH_NOR2AX3 port map( A => exe_top_i(120), B => n39, Z => 
                           src_a_22_port);
   U8 : HS65_LH_NOR2AX3 port map( A => exe_top_i(125), B => n39, Z => 
                           src_a_27_port);
   U9 : HS65_LH_NOR2AX3 port map( A => exe_top_i(126), B => n39, Z => 
                           src_a_28_port);
   U10 : HS65_LH_NOR2AX3 port map( A => exe_top_i(114), B => n38, Z => 
                           src_a_16_port);
   U11 : HS65_LH_NOR2AX3 port map( A => exe_top_i(116), B => n38, Z => 
                           src_a_18_port);
   U12 : HS65_LH_NOR2AX3 port map( A => exe_top_i(119), B => n38, Z => 
                           src_a_21_port);
   U13 : HS65_LH_NOR2AX3 port map( A => exe_top_i(122), B => n38, Z => 
                           src_a_24_port);
   U14 : HS65_LH_NOR2AX3 port map( A => exe_top_i(128), B => n38, Z => 
                           src_a_30_port);
   U15 : HS65_LH_NOR2AX3 port map( A => exe_top_i(129), B => n38, Z => 
                           src_a_31_port);
   U16 : HS65_LH_BFX9 port map( A => n48, Z => n39);
   U17 : HS65_LH_BFX9 port map( A => n48, Z => n38);
   U18 : HS65_LH_BFX9 port map( A => n48, Z => n40);
   U19 : HS65_LH_IVX9 port map( A => n7, Z => n48);
   U20 : HS65_LH_IVX9 port map( A => n44, Z => n42);
   U21 : HS65_LH_IVX9 port map( A => n44, Z => n43);
   U22 : HS65_LH_BFX9 port map( A => rst_n, Z => n47);
   U23 : HS65_LH_NAND3X5 port map( A => op_aluCtrl_alu_4_port, B => 
                           op_aluCtrl_alu_0_port, C => n8, Z => n7);
   U24 : HS65_LH_NOR3X4 port map( A => op_aluCtrl_alu_1_port, B => 
                           op_aluCtrl_alu_3_port, C => op_aluCtrl_alu_2_port, Z
                           => n8);
   U25 : HS65_LH_BFX9 port map( A => n41, Z => n44);
   U26 : HS65_LH_BFX9 port map( A => n41, Z => n45);
   U27 : HS65_LH_BFX9 port map( A => n41, Z => n46);
   U28 : HS65_LH_NOR2AX3 port map( A => s_branch_src_0_port, B => 
                           s_branch_src_1_port, Z => n9);
   U29 : HS65_LH_NOR2X6 port map( A => s_branch_src_0_port, B => 
                           s_branch_src_1_port, Z => n10);
   U30 : HS65_LH_AO22X9 port map( A => exe_top_i(100), B => n7, C => 
                           exe_top_i(13), D => n39, Z => src_a_2_port);
   U31 : HS65_LH_AO22X9 port map( A => exe_top_i(103), B => n7, C => 
                           exe_top_i(16), D => n39, Z => src_a_5_port);
   U32 : HS65_LH_AO22X9 port map( A => exe_top_i(106), B => n7, C => 
                           exe_top_i(19), D => n39, Z => src_a_8_port);
   U33 : HS65_LH_AO22X9 port map( A => exe_top_i(98), B => n7, C => 
                           exe_top_i(11), D => n40, Z => src_a_0_port);
   U34 : HS65_LH_AO22X9 port map( A => exe_top_i(102), B => n7, C => 
                           exe_top_i(15), D => n39, Z => src_a_4_port);
   U35 : HS65_LH_AO22X9 port map( A => exe_top_i(99), B => n7, C => 
                           exe_top_i(12), D => n40, Z => src_a_1_port);
   U36 : HS65_LH_AO22X9 port map( A => exe_top_i(101), B => n7, C => 
                           exe_top_i(14), D => n39, Z => src_a_3_port);
   U37 : HS65_LH_AO22X9 port map( A => exe_top_i(35), B => n46, C => 
                           exe_top_i(68), D => n43, Z => src_b_2_port);
   U38 : HS65_LH_AO22X9 port map( A => exe_top_i(33), B => n44, C => 
                           exe_top_i(66), D => n42, Z => src_b_0_port);
   U39 : HS65_LH_AO22X9 port map( A => exe_top_i(37), B => n46, C => 
                           exe_top_i(70), D => n43, Z => src_b_4_port);
   U40 : HS65_LH_AO22X9 port map( A => exe_top_i(109), B => n7, C => 
                           exe_top_i(22), D => n40, Z => src_a_11_port);
   U41 : HS65_LH_NOR2AX3 port map( A => exe_top_i(112), B => n38, Z => 
                           src_a_14_port);
   U42 : HS65_LH_NOR2AX3 port map( A => exe_top_i(115), B => n38, Z => 
                           src_a_17_port);
   U43 : HS65_LH_NOR2AX3 port map( A => exe_top_i(118), B => n39, Z => 
                           src_a_20_port);
   U44 : HS65_LH_AO22X9 port map( A => exe_top_i(108), B => n7, C => 
                           exe_top_i(21), D => n40, Z => src_a_10_port);
   U45 : HS65_LH_AO22X9 port map( A => exe_top_i(104), B => n7, C => 
                           exe_top_i(17), D => n39, Z => src_a_6_port);
   U46 : HS65_LH_AO22X9 port map( A => exe_top_i(105), B => n7, C => 
                           exe_top_i(18), D => n39, Z => src_a_7_port);
   U47 : HS65_LH_AO22X9 port map( A => exe_top_i(107), B => n7, C => 
                           exe_top_i(20), D => n39, Z => src_a_9_port);
   U48 : HS65_LH_AO22X9 port map( A => exe_top_i(40), B => n46, C => 
                           exe_top_i(73), D => n43, Z => src_b_7_port);
   U49 : HS65_LH_AO22X9 port map( A => exe_top_i(38), B => n46, C => 
                           exe_top_i(71), D => n43, Z => src_b_5_port);
   U50 : HS65_LH_AO22X9 port map( A => exe_top_i(34), B => n45, C => 
                           exe_top_i(67), D => n42, Z => src_b_1_port);
   U51 : HS65_LH_AO22X9 port map( A => exe_top_i(36), B => n46, C => 
                           exe_top_i(69), D => n43, Z => src_b_3_port);
   U52 : HS65_LH_AO22X9 port map( A => exe_top_i(39), B => n46, C => 
                           exe_top_i(72), D => n43, Z => src_b_6_port);
   U53 : HS65_LH_AO22X9 port map( A => exe_top_i(41), B => n46, C => 
                           exe_top_i(74), D => n43, Z => src_b_8_port);
   U54 : HS65_LH_AO22X9 port map( A => exe_top_i(44), B => n45, C => 
                           exe_top_i(77), D => n42, Z => src_b_11_port);
   U55 : HS65_LH_NOR2AX3 port map( A => exe_top_i(123), B => n39, Z => 
                           src_a_25_port);
   U56 : HS65_LH_NOR2AX3 port map( A => exe_top_i(117), B => n38, Z => 
                           src_a_19_port);
   U57 : HS65_LH_NOR2AX3 port map( A => exe_top_i(121), B => n38, Z => 
                           src_a_23_port);
   U58 : HS65_LH_NOR2AX3 port map( A => exe_top_i(124), B => n39, Z => 
                           src_a_26_port);
   U59 : HS65_LH_AO22X9 port map( A => exe_top_i(46), B => n45, C => 
                           exe_top_i(79), D => n42, Z => src_b_13_port);
   U60 : HS65_LH_AO22X9 port map( A => exe_top_i(45), B => n45, C => 
                           exe_top_i(78), D => n42, Z => src_b_12_port);
   U61 : HS65_LH_AO22X9 port map( A => exe_top_i(42), B => n46, C => 
                           exe_top_i(75), D => n43, Z => src_b_9_port);
   U62 : HS65_LH_AO22X9 port map( A => exe_top_i(47), B => n45, C => 
                           exe_top_i(80), D => n42, Z => src_b_14_port);
   U63 : HS65_LH_AO22X9 port map( A => exe_top_i(43), B => n45, C => 
                           exe_top_i(76), D => n42, Z => src_b_10_port);
   U64 : HS65_LH_NOR2AX3 port map( A => exe_top_i(127), B => n39, Z => 
                           src_a_29_port);
   U65 : HS65_LH_AO22X9 port map( A => exe_top_i(52), B => n45, C => 
                           exe_top_i(85), D => n42, Z => src_b_19_port);
   U66 : HS65_LH_AO22X9 port map( A => exe_top_i(48), B => n45, C => 
                           exe_top_i(81), D => n42, Z => src_b_15_port);
   U67 : HS65_LH_AO22X9 port map( A => exe_top_i(54), B => n45, C => 
                           exe_top_i(87), D => n43, Z => src_b_21_port);
   U68 : HS65_LH_AO22X9 port map( A => exe_top_i(50), B => n45, C => 
                           exe_top_i(83), D => n42, Z => src_b_17_port);
   U69 : HS65_LH_AO22X9 port map( A => exe_top_i(51), B => n45, C => 
                           exe_top_i(84), D => n42, Z => src_b_18_port);
   U70 : HS65_LH_AO22X9 port map( A => exe_top_i(53), B => n45, C => 
                           exe_top_i(86), D => n43, Z => src_b_20_port);
   U71 : HS65_LH_AO22X9 port map( A => exe_top_i(49), B => n45, C => 
                           exe_top_i(82), D => n42, Z => src_b_16_port);
   U72 : HS65_LH_BFX9 port map( A => exe_top_i(65), Z => n41);
   U73 : HS65_LH_AO22X9 port map( A => exe_top_i(56), B => n45, C => 
                           exe_top_i(89), D => n43, Z => src_b_23_port);
   U74 : HS65_LH_AO22X9 port map( A => exe_top_i(58), B => n45, C => 
                           exe_top_i(91), D => n43, Z => src_b_25_port);
   U75 : HS65_LH_AO22X9 port map( A => exe_top_i(55), B => n45, C => 
                           exe_top_i(88), D => n43, Z => src_b_22_port);
   U76 : HS65_LH_AO22X9 port map( A => exe_top_i(59), B => n45, C => 
                           exe_top_i(92), D => n43, Z => src_b_26_port);
   U77 : HS65_LH_AO22X9 port map( A => exe_top_i(57), B => n45, C => 
                           exe_top_i(90), D => n43, Z => src_b_24_port);
   U78 : HS65_LH_AO22X9 port map( A => exe_top_i(61), B => n45, C => 
                           exe_top_i(94), D => n43, Z => src_b_28_port);
   U79 : HS65_LH_AO22X9 port map( A => exe_top_i(60), B => n45, C => 
                           exe_top_i(93), D => n43, Z => src_b_27_port);
   U80 : HS65_LH_AO22X9 port map( A => exe_top_i(62), B => n46, C => 
                           exe_top_i(95), D => n43, Z => src_b_29_port);
   U81 : HS65_LH_AO22X9 port map( A => exe_top_i(63), B => n46, C => 
                           exe_top_i(96), D => n43, Z => src_b_30_port);
   U82 : HS65_LH_AO22X9 port map( A => exe_top_i(64), B => n46, C => 
                           exe_top_i(97), D => n43, Z => src_b_31_port);
   U83 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(107), C => N31, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(42), Z
                           => exe_top_o(78));
   U84 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(98), C => N22, D => 
                           n10, E => s_branch_src_1_port, F => exe_top_i(33), Z
                           => exe_top_o(69));
   U85 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(99), C => N23, D => 
                           n10, E => s_branch_src_1_port, F => exe_top_i(34), Z
                           => exe_top_o(70));
   U86 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(100), C => N24, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(35), Z
                           => exe_top_o(71));
   U87 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(101), C => N25, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(36), Z
                           => exe_top_o(72));
   U88 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(102), C => N26, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(37), Z
                           => exe_top_o(73));
   U89 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(103), C => N27, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(38), Z
                           => exe_top_o(74));
   U90 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(104), C => N28, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(39), Z
                           => exe_top_o(75));
   U91 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(105), C => N29, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(40), Z
                           => exe_top_o(76));
   U92 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(106), C => N30, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(41), Z
                           => exe_top_o(77));
   U93 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(108), C => N32, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(43), Z
                           => exe_top_o(79));
   U94 : HS65_LH_AO222X4 port map( A => n9, B => exe_top_i(109), C => N33, D =>
                           n10, E => s_branch_src_1_port, F => exe_top_i(44), Z
                           => exe_top_o(80));
   U95 : HS65_LH_BFX9 port map( A => exe_top_i(75), Z => exe_top_o(9));
   U96 : HS65_LH_BFX9 port map( A => exe_top_i(78), Z => exe_top_o(12));
   U97 : HS65_LH_BFX9 port map( A => exe_top_i(79), Z => exe_top_o(13));
   U98 : HS65_LH_BFX9 port map( A => exe_top_i(80), Z => exe_top_o(14));
   U99 : HS65_LH_BFX9 port map( A => exe_top_i(81), Z => exe_top_o(15));
   U100 : HS65_LH_BFX9 port map( A => exe_top_i(82), Z => exe_top_o(16));
   U101 : HS65_LH_BFX9 port map( A => exe_top_i(83), Z => exe_top_o(17));
   U102 : HS65_LH_BFX9 port map( A => exe_top_i(84), Z => exe_top_o(18));
   U103 : HS65_LH_BFX9 port map( A => exe_top_i(85), Z => exe_top_o(19));
   U104 : HS65_LH_BFX9 port map( A => exe_top_i(86), Z => exe_top_o(20));
   U105 : HS65_LH_BFX9 port map( A => exe_top_i(87), Z => exe_top_o(21));
   U106 : HS65_LH_BFX9 port map( A => exe_top_i(88), Z => exe_top_o(22));
   U107 : HS65_LH_BFX9 port map( A => exe_top_i(89), Z => exe_top_o(23));
   U108 : HS65_LH_BFX9 port map( A => exe_top_i(90), Z => exe_top_o(24));
   U109 : HS65_LH_BFX9 port map( A => exe_top_i(91), Z => exe_top_o(25));
   U110 : HS65_LH_BFX9 port map( A => exe_top_i(92), Z => exe_top_o(26));
   U111 : HS65_LH_BFX9 port map( A => exe_top_i(93), Z => exe_top_o(27));
   U112 : HS65_LH_BFX9 port map( A => exe_top_i(94), Z => exe_top_o(28));
   U113 : HS65_LH_BFX9 port map( A => exe_top_i(95), Z => exe_top_o(29));
   U114 : HS65_LH_BFX9 port map( A => exe_top_i(96), Z => exe_top_o(30));
   U115 : HS65_LH_BFX9 port map( A => exe_top_i(97), Z => exe_top_o(31));
   U116 : HS65_LH_BFX9 port map( A => exe_top_i(66), Z => exe_top_o(0));
   U117 : HS65_LH_BFX9 port map( A => exe_top_i(67), Z => exe_top_o(1));
   U118 : HS65_LH_BFX9 port map( A => exe_top_i(68), Z => exe_top_o(2));
   U119 : HS65_LH_BFX9 port map( A => exe_top_i(69), Z => exe_top_o(3));
   U120 : HS65_LH_BFX9 port map( A => exe_top_i(70), Z => exe_top_o(4));
   U121 : HS65_LH_BFX9 port map( A => exe_top_i(71), Z => exe_top_o(5));
   U122 : HS65_LH_BFX9 port map( A => exe_top_i(72), Z => exe_top_o(6));
   U123 : HS65_LH_BFX9 port map( A => exe_top_i(73), Z => exe_top_o(7));
   U124 : HS65_LH_BFX9 port map( A => exe_top_i(74), Z => exe_top_o(8));
   U125 : HS65_LH_BFX9 port map( A => exe_top_i(76), Z => exe_top_o(10));
   U126 : HS65_LH_BFX9 port map( A => exe_top_i(77), Z => exe_top_o(11));
   U127 : HS65_LH_AO212X4 port map( A => exe_top_i(0), B => exe_top_i(10), C =>
                           exe_top_i(5), D => n49, E => n40, Z => exe_top_o(32)
                           );
   U128 : HS65_LH_AO212X4 port map( A => exe_top_i(1), B => exe_top_i(10), C =>
                           exe_top_i(6), D => n49, E => n40, Z => exe_top_o(33)
                           );
   U129 : HS65_LH_AO212X4 port map( A => exe_top_i(2), B => exe_top_i(10), C =>
                           exe_top_i(7), D => n49, E => n40, Z => exe_top_o(34)
                           );
   U130 : HS65_LH_AO212X4 port map( A => exe_top_i(3), B => exe_top_i(10), C =>
                           exe_top_i(8), D => n49, E => n40, Z => exe_top_o(35)
                           );
   U131 : HS65_LH_AO212X4 port map( A => exe_top_i(10), B => exe_top_i(4), C =>
                           exe_top_i(9), D => n49, E => n40, Z => exe_top_o(36)
                           );
   U132 : HS65_LH_IVX9 port map( A => exe_top_i(10), Z => n49);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity id_exe is

   port( clk, rst_n, halt_i : in std_logic;  ID_EXE_i : in std_logic_vector 
         (142 downto 0);  ID_EXE_o : out std_logic_vector (142 downto 0));

end id_exe;

architecture SYN_Behavioral of id_exe is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   component HS65_LH_DFPSQX9
      port( D, CP, SN : in std_logic;  Q : out std_logic);
   end component;
   
   signal ID_EXE_o_REGA_31_port, ID_EXE_o_REGA_30_port, ID_EXE_o_REGA_29_port, 
      ID_EXE_o_REGA_28_port, ID_EXE_o_REGA_27_port, ID_EXE_o_REGA_26_port, 
      ID_EXE_o_REGA_25_port, ID_EXE_o_REGA_24_port, ID_EXE_o_REGA_23_port, 
      ID_EXE_o_REGA_22_port, ID_EXE_o_REGA_21_port, ID_EXE_o_REGA_20_port, 
      ID_EXE_o_REGA_19_port, ID_EXE_o_REGA_18_port, ID_EXE_o_REGA_17_port, 
      ID_EXE_o_REGA_16_port, ID_EXE_o_REGA_15_port, ID_EXE_o_REGA_14_port, 
      ID_EXE_o_REGA_13_port, ID_EXE_o_REGA_12_port, ID_EXE_o_REGA_11_port, 
      ID_EXE_o_REGA_10_port, ID_EXE_o_REGA_9_port, ID_EXE_o_REGA_8_port, 
      ID_EXE_o_REGA_7_port, ID_EXE_o_REGA_6_port, ID_EXE_o_REGA_5_port, 
      ID_EXE_o_REGA_4_port, ID_EXE_o_REGA_3_port, ID_EXE_o_REGA_2_port, 
      ID_EXE_o_REGA_1_port, ID_EXE_o_REGA_0_port, ID_EXE_o_REGB_31_port, 
      ID_EXE_o_REGB_30_port, ID_EXE_o_REGB_29_port, ID_EXE_o_REGB_28_port, 
      ID_EXE_o_REGB_27_port, ID_EXE_o_REGB_26_port, ID_EXE_o_REGB_25_port, 
      ID_EXE_o_REGB_24_port, ID_EXE_o_REGB_23_port, ID_EXE_o_REGB_22_port, 
      ID_EXE_o_REGB_21_port, ID_EXE_o_REGB_20_port, ID_EXE_o_REGB_19_port, 
      ID_EXE_o_REGB_18_port, ID_EXE_o_REGB_17_port, ID_EXE_o_REGB_16_port, 
      ID_EXE_o_REGB_15_port, ID_EXE_o_REGB_14_port, ID_EXE_o_REGB_13_port, 
      ID_EXE_o_REGB_12_port, ID_EXE_o_REGB_11_port, ID_EXE_o_REGB_10_port, 
      ID_EXE_o_REGB_9_port, ID_EXE_o_REGB_8_port, ID_EXE_o_REGB_7_port, 
      ID_EXE_o_REGB_6_port, ID_EXE_o_REGB_5_port, ID_EXE_o_REGB_4_port, 
      ID_EXE_o_REGB_3_port, ID_EXE_o_REGB_2_port, ID_EXE_o_REGB_1_port, 
      ID_EXE_o_REGB_0_port, ID_EXE_o_SHAMT_4_port, ID_EXE_o_SHAMT_3_port, 
      ID_EXE_o_SHAMT_2_port, ID_EXE_o_SHAMT_1_port, ID_EXE_o_SHAMT_0_port, 
      ID_EXE_o_FUNCT_5_port, ID_EXE_o_FUNCT_4_port, ID_EXE_o_FUNCT_3_port, 
      ID_EXE_o_FUNCT_2_port, ID_EXE_o_FUNCT_1_port, ID_EXE_o_FUNCT_0_port, 
      ID_EXE_o_SIGN_EXTEND_31_port, ID_EXE_o_SIGN_EXTEND_30_port, 
      ID_EXE_o_SIGN_EXTEND_29_port, ID_EXE_o_SIGN_EXTEND_28_port, 
      ID_EXE_o_SIGN_EXTEND_27_port, ID_EXE_o_SIGN_EXTEND_26_port, 
      ID_EXE_o_SIGN_EXTEND_25_port, ID_EXE_o_SIGN_EXTEND_24_port, 
      ID_EXE_o_SIGN_EXTEND_23_port, ID_EXE_o_SIGN_EXTEND_22_port, 
      ID_EXE_o_SIGN_EXTEND_21_port, ID_EXE_o_SIGN_EXTEND_20_port, 
      ID_EXE_o_SIGN_EXTEND_19_port, ID_EXE_o_SIGN_EXTEND_18_port, 
      ID_EXE_o_SIGN_EXTEND_17_port, ID_EXE_o_SIGN_EXTEND_16_port, 
      ID_EXE_o_SIGN_EXTEND_15_port, ID_EXE_o_SIGN_EXTEND_14_port, 
      ID_EXE_o_SIGN_EXTEND_13_port, ID_EXE_o_SIGN_EXTEND_12_port, 
      ID_EXE_o_SIGN_EXTEND_11_port, ID_EXE_o_SIGN_EXTEND_10_port, 
      ID_EXE_o_SIGN_EXTEND_9_port, ID_EXE_o_SIGN_EXTEND_8_port, 
      ID_EXE_o_SIGN_EXTEND_7_port, ID_EXE_o_SIGN_EXTEND_6_port, 
      ID_EXE_o_SIGN_EXTEND_5_port, ID_EXE_o_SIGN_EXTEND_4_port, 
      ID_EXE_o_SIGN_EXTEND_3_port, ID_EXE_o_SIGN_EXTEND_2_port, 
      ID_EXE_o_SIGN_EXTEND_1_port, ID_EXE_o_SIGN_EXTEND_0_port, 
      ID_EXE_o_PC_PLUS1_11_port, ID_EXE_o_PC_PLUS1_10_port, 
      ID_EXE_o_PC_PLUS1_9_port, ID_EXE_o_PC_PLUS1_8_port, 
      ID_EXE_o_PC_PLUS1_7_port, ID_EXE_o_PC_PLUS1_6_port, 
      ID_EXE_o_PC_PLUS1_5_port, ID_EXE_o_PC_PLUS1_4_port, 
      ID_EXE_o_PC_PLUS1_3_port, ID_EXE_o_PC_PLUS1_2_port, 
      ID_EXE_o_PC_PLUS1_1_port, ID_EXE_o_PC_PLUS1_0_port, ID_EXE_o_RS_4_port, 
      ID_EXE_o_RS_3_port, ID_EXE_o_RS_2_port, ID_EXE_o_RS_1_port, 
      ID_EXE_o_RS_0_port, ID_EXE_o_RT_4_port, ID_EXE_o_RT_3_port, 
      ID_EXE_o_RT_2_port, ID_EXE_o_RT_1_port, ID_EXE_o_RT_0_port, 
      ID_EXE_o_RD_4_port, ID_EXE_o_RD_3_port, ID_EXE_o_RD_2_port, 
      ID_EXE_o_RD_1_port, ID_EXE_o_RD_0_port, ID_EXE_o_ALUSRC_B_port, 
      ID_EXE_o_MEMTOREG_port, ID_EXE_o_REGWRITE_port, ID_EXE_o_MEMWEN_N_port, 
      ID_EXE_o_CALU_OP_3_port, ID_EXE_o_CALU_OP_2_port, ID_EXE_o_CALU_OP_1_port
      , ID_EXE_o_CALU_OP_0_port, ID_EXE_o_REGDST_port, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n1, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180 : std_logic;

begin
   ID_EXE_o <= ( ID_EXE_o_REGA_31_port, ID_EXE_o_REGA_30_port, 
      ID_EXE_o_REGA_29_port, ID_EXE_o_REGA_28_port, ID_EXE_o_REGA_27_port, 
      ID_EXE_o_REGA_26_port, ID_EXE_o_REGA_25_port, ID_EXE_o_REGA_24_port, 
      ID_EXE_o_REGA_23_port, ID_EXE_o_REGA_22_port, ID_EXE_o_REGA_21_port, 
      ID_EXE_o_REGA_20_port, ID_EXE_o_REGA_19_port, ID_EXE_o_REGA_18_port, 
      ID_EXE_o_REGA_17_port, ID_EXE_o_REGA_16_port, ID_EXE_o_REGA_15_port, 
      ID_EXE_o_REGA_14_port, ID_EXE_o_REGA_13_port, ID_EXE_o_REGA_12_port, 
      ID_EXE_o_REGA_11_port, ID_EXE_o_REGA_10_port, ID_EXE_o_REGA_9_port, 
      ID_EXE_o_REGA_8_port, ID_EXE_o_REGA_7_port, ID_EXE_o_REGA_6_port, 
      ID_EXE_o_REGA_5_port, ID_EXE_o_REGA_4_port, ID_EXE_o_REGA_3_port, 
      ID_EXE_o_REGA_2_port, ID_EXE_o_REGA_1_port, ID_EXE_o_REGA_0_port, 
      ID_EXE_o_REGB_31_port, ID_EXE_o_REGB_30_port, ID_EXE_o_REGB_29_port, 
      ID_EXE_o_REGB_28_port, ID_EXE_o_REGB_27_port, ID_EXE_o_REGB_26_port, 
      ID_EXE_o_REGB_25_port, ID_EXE_o_REGB_24_port, ID_EXE_o_REGB_23_port, 
      ID_EXE_o_REGB_22_port, ID_EXE_o_REGB_21_port, ID_EXE_o_REGB_20_port, 
      ID_EXE_o_REGB_19_port, ID_EXE_o_REGB_18_port, ID_EXE_o_REGB_17_port, 
      ID_EXE_o_REGB_16_port, ID_EXE_o_REGB_15_port, ID_EXE_o_REGB_14_port, 
      ID_EXE_o_REGB_13_port, ID_EXE_o_REGB_12_port, ID_EXE_o_REGB_11_port, 
      ID_EXE_o_REGB_10_port, ID_EXE_o_REGB_9_port, ID_EXE_o_REGB_8_port, 
      ID_EXE_o_REGB_7_port, ID_EXE_o_REGB_6_port, ID_EXE_o_REGB_5_port, 
      ID_EXE_o_REGB_4_port, ID_EXE_o_REGB_3_port, ID_EXE_o_REGB_2_port, 
      ID_EXE_o_REGB_1_port, ID_EXE_o_REGB_0_port, ID_EXE_o_SHAMT_4_port, 
      ID_EXE_o_SHAMT_3_port, ID_EXE_o_SHAMT_2_port, ID_EXE_o_SHAMT_1_port, 
      ID_EXE_o_SHAMT_0_port, ID_EXE_o_FUNCT_5_port, ID_EXE_o_FUNCT_4_port, 
      ID_EXE_o_FUNCT_3_port, ID_EXE_o_FUNCT_2_port, ID_EXE_o_FUNCT_1_port, 
      ID_EXE_o_FUNCT_0_port, ID_EXE_o_SIGN_EXTEND_31_port, 
      ID_EXE_o_SIGN_EXTEND_30_port, ID_EXE_o_SIGN_EXTEND_29_port, 
      ID_EXE_o_SIGN_EXTEND_28_port, ID_EXE_o_SIGN_EXTEND_27_port, 
      ID_EXE_o_SIGN_EXTEND_26_port, ID_EXE_o_SIGN_EXTEND_25_port, 
      ID_EXE_o_SIGN_EXTEND_24_port, ID_EXE_o_SIGN_EXTEND_23_port, 
      ID_EXE_o_SIGN_EXTEND_22_port, ID_EXE_o_SIGN_EXTEND_21_port, 
      ID_EXE_o_SIGN_EXTEND_20_port, ID_EXE_o_SIGN_EXTEND_19_port, 
      ID_EXE_o_SIGN_EXTEND_18_port, ID_EXE_o_SIGN_EXTEND_17_port, 
      ID_EXE_o_SIGN_EXTEND_16_port, ID_EXE_o_SIGN_EXTEND_15_port, 
      ID_EXE_o_SIGN_EXTEND_14_port, ID_EXE_o_SIGN_EXTEND_13_port, 
      ID_EXE_o_SIGN_EXTEND_12_port, ID_EXE_o_SIGN_EXTEND_11_port, 
      ID_EXE_o_SIGN_EXTEND_10_port, ID_EXE_o_SIGN_EXTEND_9_port, 
      ID_EXE_o_SIGN_EXTEND_8_port, ID_EXE_o_SIGN_EXTEND_7_port, 
      ID_EXE_o_SIGN_EXTEND_6_port, ID_EXE_o_SIGN_EXTEND_5_port, 
      ID_EXE_o_SIGN_EXTEND_4_port, ID_EXE_o_SIGN_EXTEND_3_port, 
      ID_EXE_o_SIGN_EXTEND_2_port, ID_EXE_o_SIGN_EXTEND_1_port, 
      ID_EXE_o_SIGN_EXTEND_0_port, ID_EXE_o_PC_PLUS1_11_port, 
      ID_EXE_o_PC_PLUS1_10_port, ID_EXE_o_PC_PLUS1_9_port, 
      ID_EXE_o_PC_PLUS1_8_port, ID_EXE_o_PC_PLUS1_7_port, 
      ID_EXE_o_PC_PLUS1_6_port, ID_EXE_o_PC_PLUS1_5_port, 
      ID_EXE_o_PC_PLUS1_4_port, ID_EXE_o_PC_PLUS1_3_port, 
      ID_EXE_o_PC_PLUS1_2_port, ID_EXE_o_PC_PLUS1_1_port, 
      ID_EXE_o_PC_PLUS1_0_port, ID_EXE_o_RS_4_port, ID_EXE_o_RS_3_port, 
      ID_EXE_o_RS_2_port, ID_EXE_o_RS_1_port, ID_EXE_o_RS_0_port, 
      ID_EXE_o_RT_4_port, ID_EXE_o_RT_3_port, ID_EXE_o_RT_2_port, 
      ID_EXE_o_RT_1_port, ID_EXE_o_RT_0_port, ID_EXE_o_RD_4_port, 
      ID_EXE_o_RD_3_port, ID_EXE_o_RD_2_port, ID_EXE_o_RD_1_port, 
      ID_EXE_o_RD_0_port, ID_EXE_o_ALUSRC_B_port, ID_EXE_o_MEMTOREG_port, 
      ID_EXE_o_REGWRITE_port, ID_EXE_o_MEMWEN_N_port, ID_EXE_o_CALU_OP_3_port, 
      ID_EXE_o_CALU_OP_2_port, ID_EXE_o_CALU_OP_1_port, ID_EXE_o_CALU_OP_0_port
      , ID_EXE_o_REGDST_port );
   
   id_exe_c_reg_REGA_31_inst : HS65_LH_DFPRQX9 port map( D => n144, CP => clk, 
                           RN => n164, Q => ID_EXE_o_REGA_31_port);
   id_exe_c_reg_REGA_30_inst : HS65_LH_DFPRQX9 port map( D => n143, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_30_port);
   id_exe_c_reg_REGA_29_inst : HS65_LH_DFPRQX9 port map( D => n142, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_29_port);
   id_exe_c_reg_REGA_28_inst : HS65_LH_DFPRQX9 port map( D => n141, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_28_port);
   id_exe_c_reg_REGA_27_inst : HS65_LH_DFPRQX9 port map( D => n140, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_27_port);
   id_exe_c_reg_REGA_26_inst : HS65_LH_DFPRQX9 port map( D => n139, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_26_port);
   id_exe_c_reg_REGA_25_inst : HS65_LH_DFPRQX9 port map( D => n138, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_25_port);
   id_exe_c_reg_REGA_24_inst : HS65_LH_DFPRQX9 port map( D => n137, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_24_port);
   id_exe_c_reg_REGA_23_inst : HS65_LH_DFPRQX9 port map( D => n136, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_23_port);
   id_exe_c_reg_REGA_22_inst : HS65_LH_DFPRQX9 port map( D => n135, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_22_port);
   id_exe_c_reg_REGA_21_inst : HS65_LH_DFPRQX9 port map( D => n134, CP => clk, 
                           RN => n175, Q => ID_EXE_o_REGA_21_port);
   id_exe_c_reg_REGA_20_inst : HS65_LH_DFPRQX9 port map( D => n133, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_20_port);
   id_exe_c_reg_REGA_19_inst : HS65_LH_DFPRQX9 port map( D => n132, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_19_port);
   id_exe_c_reg_REGA_18_inst : HS65_LH_DFPRQX9 port map( D => n131, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_18_port);
   id_exe_c_reg_REGA_17_inst : HS65_LH_DFPRQX9 port map( D => n130, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_17_port);
   id_exe_c_reg_REGA_16_inst : HS65_LH_DFPRQX9 port map( D => n129, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_16_port);
   id_exe_c_reg_REGA_15_inst : HS65_LH_DFPRQX9 port map( D => n128, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_15_port);
   id_exe_c_reg_REGA_14_inst : HS65_LH_DFPRQX9 port map( D => n127, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_14_port);
   id_exe_c_reg_REGA_13_inst : HS65_LH_DFPRQX9 port map( D => n126, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_13_port);
   id_exe_c_reg_REGA_12_inst : HS65_LH_DFPRQX9 port map( D => n125, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_12_port);
   id_exe_c_reg_REGA_11_inst : HS65_LH_DFPRQX9 port map( D => n124, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_11_port);
   id_exe_c_reg_REGA_10_inst : HS65_LH_DFPRQX9 port map( D => n123, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_10_port);
   id_exe_c_reg_REGA_9_inst : HS65_LH_DFPRQX9 port map( D => n122, CP => clk, 
                           RN => n174, Q => ID_EXE_o_REGA_9_port);
   id_exe_c_reg_REGA_8_inst : HS65_LH_DFPRQX9 port map( D => n121, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_8_port);
   id_exe_c_reg_REGA_7_inst : HS65_LH_DFPRQX9 port map( D => n120, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_7_port);
   id_exe_c_reg_REGA_6_inst : HS65_LH_DFPRQX9 port map( D => n119, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_6_port);
   id_exe_c_reg_REGA_5_inst : HS65_LH_DFPRQX9 port map( D => n118, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_5_port);
   id_exe_c_reg_REGA_4_inst : HS65_LH_DFPRQX9 port map( D => n117, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_4_port);
   id_exe_c_reg_REGA_3_inst : HS65_LH_DFPRQX9 port map( D => n116, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_3_port);
   id_exe_c_reg_REGA_2_inst : HS65_LH_DFPRQX9 port map( D => n115, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_2_port);
   id_exe_c_reg_REGA_1_inst : HS65_LH_DFPRQX9 port map( D => n114, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_1_port);
   id_exe_c_reg_REGA_0_inst : HS65_LH_DFPRQX9 port map( D => n113, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGA_0_port);
   id_exe_c_reg_REGB_31_inst : HS65_LH_DFPRQX9 port map( D => n112, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGB_31_port);
   id_exe_c_reg_REGB_30_inst : HS65_LH_DFPRQX9 port map( D => n111, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGB_30_port);
   id_exe_c_reg_REGB_29_inst : HS65_LH_DFPRQX9 port map( D => n110, CP => clk, 
                           RN => n173, Q => ID_EXE_o_REGB_29_port);
   id_exe_c_reg_REGB_28_inst : HS65_LH_DFPRQX9 port map( D => n109, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_28_port);
   id_exe_c_reg_REGB_27_inst : HS65_LH_DFPRQX9 port map( D => n108, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_27_port);
   id_exe_c_reg_REGB_26_inst : HS65_LH_DFPRQX9 port map( D => n107, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_26_port);
   id_exe_c_reg_REGB_25_inst : HS65_LH_DFPRQX9 port map( D => n106, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_25_port);
   id_exe_c_reg_REGB_24_inst : HS65_LH_DFPRQX9 port map( D => n105, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_24_port);
   id_exe_c_reg_REGB_23_inst : HS65_LH_DFPRQX9 port map( D => n104, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_23_port);
   id_exe_c_reg_REGB_22_inst : HS65_LH_DFPRQX9 port map( D => n103, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_22_port);
   id_exe_c_reg_REGB_21_inst : HS65_LH_DFPRQX9 port map( D => n102, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_21_port);
   id_exe_c_reg_REGB_20_inst : HS65_LH_DFPRQX9 port map( D => n101, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_20_port);
   id_exe_c_reg_REGB_19_inst : HS65_LH_DFPRQX9 port map( D => n100, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_19_port);
   id_exe_c_reg_REGB_18_inst : HS65_LH_DFPRQX9 port map( D => n99, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_18_port);
   id_exe_c_reg_REGB_17_inst : HS65_LH_DFPRQX9 port map( D => n98, CP => clk, 
                           RN => n172, Q => ID_EXE_o_REGB_17_port);
   id_exe_c_reg_REGB_16_inst : HS65_LH_DFPRQX9 port map( D => n97, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_16_port);
   id_exe_c_reg_REGB_15_inst : HS65_LH_DFPRQX9 port map( D => n96, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_15_port);
   id_exe_c_reg_REGB_14_inst : HS65_LH_DFPRQX9 port map( D => n95, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_14_port);
   id_exe_c_reg_REGB_13_inst : HS65_LH_DFPRQX9 port map( D => n94, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_13_port);
   id_exe_c_reg_REGB_12_inst : HS65_LH_DFPRQX9 port map( D => n93, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_12_port);
   id_exe_c_reg_REGB_11_inst : HS65_LH_DFPRQX9 port map( D => n92, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_11_port);
   id_exe_c_reg_REGB_10_inst : HS65_LH_DFPRQX9 port map( D => n91, CP => clk, 
                           RN => n171, Q => ID_EXE_o_REGB_10_port);
   id_exe_c_reg_REGB_9_inst : HS65_LH_DFPRQX9 port map( D => n90, CP => clk, RN
                           => n171, Q => ID_EXE_o_REGB_9_port);
   id_exe_c_reg_REGB_8_inst : HS65_LH_DFPRQX9 port map( D => n89, CP => clk, RN
                           => n171, Q => ID_EXE_o_REGB_8_port);
   id_exe_c_reg_REGB_7_inst : HS65_LH_DFPRQX9 port map( D => n88, CP => clk, RN
                           => n171, Q => ID_EXE_o_REGB_7_port);
   id_exe_c_reg_REGB_6_inst : HS65_LH_DFPRQX9 port map( D => n87, CP => clk, RN
                           => n171, Q => ID_EXE_o_REGB_6_port);
   id_exe_c_reg_REGB_5_inst : HS65_LH_DFPRQX9 port map( D => n86, CP => clk, RN
                           => n171, Q => ID_EXE_o_REGB_5_port);
   id_exe_c_reg_REGB_4_inst : HS65_LH_DFPRQX9 port map( D => n85, CP => clk, RN
                           => n170, Q => ID_EXE_o_REGB_4_port);
   id_exe_c_reg_REGB_3_inst : HS65_LH_DFPRQX9 port map( D => n84, CP => clk, RN
                           => n170, Q => ID_EXE_o_REGB_3_port);
   id_exe_c_reg_REGB_2_inst : HS65_LH_DFPRQX9 port map( D => n83, CP => clk, RN
                           => n170, Q => ID_EXE_o_REGB_2_port);
   id_exe_c_reg_REGB_1_inst : HS65_LH_DFPRQX9 port map( D => n82, CP => clk, RN
                           => n170, Q => ID_EXE_o_REGB_1_port);
   id_exe_c_reg_REGB_0_inst : HS65_LH_DFPRQX9 port map( D => n81, CP => clk, RN
                           => n170, Q => ID_EXE_o_REGB_0_port);
   id_exe_c_reg_SHAMT_4_inst : HS65_LH_DFPRQX9 port map( D => n80, CP => clk, 
                           RN => n170, Q => ID_EXE_o_SHAMT_4_port);
   id_exe_c_reg_SHAMT_3_inst : HS65_LH_DFPRQX9 port map( D => n79, CP => clk, 
                           RN => n170, Q => ID_EXE_o_SHAMT_3_port);
   id_exe_c_reg_SHAMT_2_inst : HS65_LH_DFPRQX9 port map( D => n78, CP => clk, 
                           RN => n170, Q => ID_EXE_o_SHAMT_2_port);
   id_exe_c_reg_SHAMT_1_inst : HS65_LH_DFPRQX9 port map( D => n77, CP => clk, 
                           RN => n170, Q => ID_EXE_o_SHAMT_1_port);
   id_exe_c_reg_SHAMT_0_inst : HS65_LH_DFPRQX9 port map( D => n76, CP => clk, 
                           RN => n170, Q => ID_EXE_o_SHAMT_0_port);
   id_exe_c_reg_FUNCT_5_inst : HS65_LH_DFPRQX9 port map( D => n75, CP => clk, 
                           RN => n170, Q => ID_EXE_o_FUNCT_5_port);
   id_exe_c_reg_FUNCT_4_inst : HS65_LH_DFPRQX9 port map( D => n74, CP => clk, 
                           RN => n170, Q => ID_EXE_o_FUNCT_4_port);
   id_exe_c_reg_FUNCT_3_inst : HS65_LH_DFPRQX9 port map( D => n73, CP => clk, 
                           RN => n169, Q => ID_EXE_o_FUNCT_3_port);
   id_exe_c_reg_FUNCT_2_inst : HS65_LH_DFPRQX9 port map( D => n72, CP => clk, 
                           RN => n169, Q => ID_EXE_o_FUNCT_2_port);
   id_exe_c_reg_FUNCT_1_inst : HS65_LH_DFPRQX9 port map( D => n71, CP => clk, 
                           RN => n169, Q => ID_EXE_o_FUNCT_1_port);
   id_exe_c_reg_FUNCT_0_inst : HS65_LH_DFPRQX9 port map( D => n70, CP => clk, 
                           RN => n169, Q => ID_EXE_o_FUNCT_0_port);
   id_exe_c_reg_SIGN_EXTEND_31_inst : HS65_LH_DFPRQX9 port map( D => n69, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_31_port);
   id_exe_c_reg_SIGN_EXTEND_30_inst : HS65_LH_DFPRQX9 port map( D => n68, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_30_port);
   id_exe_c_reg_SIGN_EXTEND_29_inst : HS65_LH_DFPRQX9 port map( D => n67, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_29_port);
   id_exe_c_reg_SIGN_EXTEND_28_inst : HS65_LH_DFPRQX9 port map( D => n66, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_28_port);
   id_exe_c_reg_SIGN_EXTEND_27_inst : HS65_LH_DFPRQX9 port map( D => n65, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_27_port);
   id_exe_c_reg_SIGN_EXTEND_26_inst : HS65_LH_DFPRQX9 port map( D => n64, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_26_port);
   id_exe_c_reg_SIGN_EXTEND_25_inst : HS65_LH_DFPRQX9 port map( D => n63, CP =>
                           clk, RN => n169, Q => ID_EXE_o_SIGN_EXTEND_25_port);
   id_exe_c_reg_SIGN_EXTEND_24_inst : HS65_LH_DFPRQX9 port map( D => n62, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_24_port);
   id_exe_c_reg_SIGN_EXTEND_23_inst : HS65_LH_DFPRQX9 port map( D => n61, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_23_port);
   id_exe_c_reg_SIGN_EXTEND_22_inst : HS65_LH_DFPRQX9 port map( D => n60, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_22_port);
   id_exe_c_reg_SIGN_EXTEND_21_inst : HS65_LH_DFPRQX9 port map( D => n59, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_21_port);
   id_exe_c_reg_SIGN_EXTEND_20_inst : HS65_LH_DFPRQX9 port map( D => n58, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_20_port);
   id_exe_c_reg_SIGN_EXTEND_19_inst : HS65_LH_DFPRQX9 port map( D => n57, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_19_port);
   id_exe_c_reg_SIGN_EXTEND_18_inst : HS65_LH_DFPRQX9 port map( D => n56, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_18_port);
   id_exe_c_reg_SIGN_EXTEND_17_inst : HS65_LH_DFPRQX9 port map( D => n55, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_17_port);
   id_exe_c_reg_SIGN_EXTEND_16_inst : HS65_LH_DFPRQX9 port map( D => n54, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_16_port);
   id_exe_c_reg_SIGN_EXTEND_15_inst : HS65_LH_DFPRQX9 port map( D => n53, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_15_port);
   id_exe_c_reg_SIGN_EXTEND_14_inst : HS65_LH_DFPRQX9 port map( D => n52, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_14_port);
   id_exe_c_reg_SIGN_EXTEND_13_inst : HS65_LH_DFPRQX9 port map( D => n51, CP =>
                           clk, RN => n168, Q => ID_EXE_o_SIGN_EXTEND_13_port);
   id_exe_c_reg_SIGN_EXTEND_12_inst : HS65_LH_DFPRQX9 port map( D => n50, CP =>
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_12_port);
   id_exe_c_reg_SIGN_EXTEND_11_inst : HS65_LH_DFPRQX9 port map( D => n49, CP =>
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_11_port);
   id_exe_c_reg_SIGN_EXTEND_10_inst : HS65_LH_DFPRQX9 port map( D => n48, CP =>
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_10_port);
   id_exe_c_reg_SIGN_EXTEND_9_inst : HS65_LH_DFPRQX9 port map( D => n47, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_9_port);
   id_exe_c_reg_SIGN_EXTEND_8_inst : HS65_LH_DFPRQX9 port map( D => n46, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_8_port);
   id_exe_c_reg_SIGN_EXTEND_7_inst : HS65_LH_DFPRQX9 port map( D => n45, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_7_port);
   id_exe_c_reg_SIGN_EXTEND_6_inst : HS65_LH_DFPRQX9 port map( D => n44, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_6_port);
   id_exe_c_reg_SIGN_EXTEND_5_inst : HS65_LH_DFPRQX9 port map( D => n43, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_5_port);
   id_exe_c_reg_SIGN_EXTEND_4_inst : HS65_LH_DFPRQX9 port map( D => n42, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_4_port);
   id_exe_c_reg_SIGN_EXTEND_3_inst : HS65_LH_DFPRQX9 port map( D => n41, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_3_port);
   id_exe_c_reg_SIGN_EXTEND_2_inst : HS65_LH_DFPRQX9 port map( D => n40, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_2_port);
   id_exe_c_reg_SIGN_EXTEND_1_inst : HS65_LH_DFPRQX9 port map( D => n39, CP => 
                           clk, RN => n167, Q => ID_EXE_o_SIGN_EXTEND_1_port);
   id_exe_c_reg_SIGN_EXTEND_0_inst : HS65_LH_DFPRQX9 port map( D => n38, CP => 
                           clk, RN => n166, Q => ID_EXE_o_SIGN_EXTEND_0_port);
   id_exe_c_reg_PC_PLUS1_11_inst : HS65_LH_DFPRQX9 port map( D => n37, CP => 
                           clk, RN => n166, Q => ID_EXE_o_PC_PLUS1_11_port);
   id_exe_c_reg_PC_PLUS1_10_inst : HS65_LH_DFPRQX9 port map( D => n36, CP => 
                           clk, RN => n166, Q => ID_EXE_o_PC_PLUS1_10_port);
   id_exe_c_reg_PC_PLUS1_9_inst : HS65_LH_DFPRQX9 port map( D => n35, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_9_port);
   id_exe_c_reg_PC_PLUS1_8_inst : HS65_LH_DFPRQX9 port map( D => n34, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_8_port);
   id_exe_c_reg_PC_PLUS1_7_inst : HS65_LH_DFPRQX9 port map( D => n33, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_7_port);
   id_exe_c_reg_PC_PLUS1_6_inst : HS65_LH_DFPRQX9 port map( D => n32, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_6_port);
   id_exe_c_reg_PC_PLUS1_5_inst : HS65_LH_DFPRQX9 port map( D => n31, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_5_port);
   id_exe_c_reg_PC_PLUS1_4_inst : HS65_LH_DFPRQX9 port map( D => n30, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_4_port);
   id_exe_c_reg_PC_PLUS1_3_inst : HS65_LH_DFPRQX9 port map( D => n29, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_3_port);
   id_exe_c_reg_PC_PLUS1_2_inst : HS65_LH_DFPRQX9 port map( D => n28, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_2_port);
   id_exe_c_reg_PC_PLUS1_1_inst : HS65_LH_DFPRQX9 port map( D => n27, CP => clk
                           , RN => n166, Q => ID_EXE_o_PC_PLUS1_1_port);
   id_exe_c_reg_PC_PLUS1_0_inst : HS65_LH_DFPRQX9 port map( D => n26, CP => clk
                           , RN => n165, Q => ID_EXE_o_PC_PLUS1_0_port);
   id_exe_c_reg_RS_4_inst : HS65_LH_DFPRQX9 port map( D => n25, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RS_4_port);
   id_exe_c_reg_RS_3_inst : HS65_LH_DFPRQX9 port map( D => n24, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RS_3_port);
   id_exe_c_reg_RS_2_inst : HS65_LH_DFPRQX9 port map( D => n23, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RS_2_port);
   id_exe_c_reg_RS_1_inst : HS65_LH_DFPRQX9 port map( D => n22, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RS_1_port);
   id_exe_c_reg_RS_0_inst : HS65_LH_DFPRQX9 port map( D => n21, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RS_0_port);
   id_exe_c_reg_RT_4_inst : HS65_LH_DFPRQX9 port map( D => n20, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RT_4_port);
   id_exe_c_reg_RT_3_inst : HS65_LH_DFPRQX9 port map( D => n19, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RT_3_port);
   id_exe_c_reg_RT_2_inst : HS65_LH_DFPRQX9 port map( D => n18, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RT_2_port);
   id_exe_c_reg_RT_1_inst : HS65_LH_DFPRQX9 port map( D => n17, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RT_1_port);
   id_exe_c_reg_RT_0_inst : HS65_LH_DFPRQX9 port map( D => n16, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RT_0_port);
   id_exe_c_reg_RD_4_inst : HS65_LH_DFPRQX9 port map( D => n15, CP => clk, RN 
                           => n165, Q => ID_EXE_o_RD_4_port);
   id_exe_c_reg_RD_3_inst : HS65_LH_DFPRQX9 port map( D => n14, CP => clk, RN 
                           => n164, Q => ID_EXE_o_RD_3_port);
   id_exe_c_reg_RD_2_inst : HS65_LH_DFPRQX9 port map( D => n13, CP => clk, RN 
                           => n164, Q => ID_EXE_o_RD_2_port);
   id_exe_c_reg_RD_1_inst : HS65_LH_DFPRQX9 port map( D => n12, CP => clk, RN 
                           => n164, Q => ID_EXE_o_RD_1_port);
   id_exe_c_reg_RD_0_inst : HS65_LH_DFPRQX9 port map( D => n11, CP => clk, RN 
                           => n164, Q => ID_EXE_o_RD_0_port);
   id_exe_c_reg_ALUSRC_B_inst : HS65_LH_DFPRQX9 port map( D => n10, CP => clk, 
                           RN => n164, Q => ID_EXE_o_ALUSRC_B_port);
   id_exe_c_reg_MEMTOREG_inst : HS65_LH_DFPRQX9 port map( D => n9, CP => clk, 
                           RN => n164, Q => ID_EXE_o_MEMTOREG_port);
   id_exe_c_reg_REGWRITE_inst : HS65_LH_DFPRQX9 port map( D => n8, CP => clk, 
                           RN => n164, Q => ID_EXE_o_REGWRITE_port);
   id_exe_c_reg_MEMWEN_N_inst : HS65_LH_DFPSQX9 port map( D => n7, CP => clk, 
                           SN => n175, Q => ID_EXE_o_MEMWEN_N_port);
   id_exe_c_reg_CALU_OP_3_inst : HS65_LH_DFPRQX9 port map( D => n6, CP => clk, 
                           RN => n164, Q => ID_EXE_o_CALU_OP_3_port);
   id_exe_c_reg_CALU_OP_2_inst : HS65_LH_DFPRQX9 port map( D => n5, CP => clk, 
                           RN => n164, Q => ID_EXE_o_CALU_OP_2_port);
   id_exe_c_reg_CALU_OP_1_inst : HS65_LH_DFPRQX9 port map( D => n4, CP => clk, 
                           RN => n164, Q => ID_EXE_o_CALU_OP_1_port);
   id_exe_c_reg_CALU_OP_0_inst : HS65_LH_DFPRQX9 port map( D => n3, CP => clk, 
                           RN => n164, Q => ID_EXE_o_CALU_OP_0_port);
   id_exe_c_reg_REGDST_inst : HS65_LH_DFPRQX9 port map( D => n2, CP => clk, RN 
                           => n169, Q => ID_EXE_o_REGDST_port);
   U2 : HS65_LH_BFX9 port map( A => n179, Z => n165);
   U3 : HS65_LH_BFX9 port map( A => n179, Z => n166);
   U4 : HS65_LH_BFX9 port map( A => n178, Z => n167);
   U5 : HS65_LH_BFX9 port map( A => n178, Z => n168);
   U6 : HS65_LH_BFX9 port map( A => n178, Z => n169);
   U7 : HS65_LH_BFX9 port map( A => n177, Z => n170);
   U8 : HS65_LH_BFX9 port map( A => n177, Z => n171);
   U9 : HS65_LH_BFX9 port map( A => n177, Z => n172);
   U10 : HS65_LH_BFX9 port map( A => n176, Z => n173);
   U11 : HS65_LH_BFX9 port map( A => n176, Z => n174);
   U12 : HS65_LH_BFX9 port map( A => n179, Z => n164);
   U13 : HS65_LH_BFX9 port map( A => n176, Z => n175);
   U14 : HS65_LH_BFX9 port map( A => n163, Z => n178);
   U15 : HS65_LH_BFX9 port map( A => n162, Z => n177);
   U16 : HS65_LH_BFX9 port map( A => n162, Z => n176);
   U17 : HS65_LH_BFX9 port map( A => n163, Z => n179);
   U18 : HS65_LH_BFX9 port map( A => n1, Z => n150);
   U19 : HS65_LH_BFX9 port map( A => n1, Z => n151);
   U20 : HS65_LH_BFX9 port map( A => n1, Z => n152);
   U21 : HS65_LH_BFX9 port map( A => n145, Z => n153);
   U22 : HS65_LH_BFX9 port map( A => n145, Z => n154);
   U23 : HS65_LH_BFX9 port map( A => n145, Z => n155);
   U24 : HS65_LH_BFX9 port map( A => n146, Z => n156);
   U25 : HS65_LH_BFX9 port map( A => n146, Z => n157);
   U26 : HS65_LH_BFX9 port map( A => n146, Z => n158);
   U27 : HS65_LH_BFX9 port map( A => n147, Z => n159);
   U28 : HS65_LH_BFX9 port map( A => n147, Z => n160);
   U29 : HS65_LH_BFX9 port map( A => n147, Z => n161);
   U30 : HS65_LH_BFX9 port map( A => rst_n, Z => n162);
   U31 : HS65_LH_BFX9 port map( A => rst_n, Z => n163);
   U32 : HS65_LH_BFX9 port map( A => n149, Z => n1);
   U33 : HS65_LH_BFX9 port map( A => n149, Z => n145);
   U34 : HS65_LH_BFX9 port map( A => n148, Z => n146);
   U35 : HS65_LH_BFX9 port map( A => n148, Z => n147);
   U36 : HS65_LH_BFX9 port map( A => n180, Z => n149);
   U37 : HS65_LH_BFX9 port map( A => n180, Z => n148);
   U38 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_0_port, B => halt_i, C => 
                           ID_EXE_i(111), D => n159, Z => n113);
   U39 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_1_port, B => halt_i, C => 
                           ID_EXE_i(112), D => n159, Z => n114);
   U40 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_2_port, B => halt_i, C => 
                           ID_EXE_i(113), D => n159, Z => n115);
   U41 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_3_port, B => halt_i, C => 
                           ID_EXE_i(114), D => n159, Z => n116);
   U42 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_4_port, B => halt_i, C => 
                           ID_EXE_i(115), D => n159, Z => n117);
   U43 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_5_port, B => halt_i, C => 
                           ID_EXE_i(116), D => n159, Z => n118);
   U44 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_6_port, B => halt_i, C => 
                           ID_EXE_i(117), D => n159, Z => n119);
   U45 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_7_port, B => halt_i, C => 
                           ID_EXE_i(118), D => n159, Z => n120);
   U46 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_8_port, B => halt_i, C => 
                           ID_EXE_i(119), D => n159, Z => n121);
   U47 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_9_port, B => halt_i, C => 
                           ID_EXE_i(120), D => n160, Z => n122);
   U48 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_10_port, B => halt_i, C =>
                           ID_EXE_i(121), D => n160, Z => n123);
   U49 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_11_port, B => halt_i, C =>
                           ID_EXE_i(122), D => n160, Z => n124);
   U50 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_12_port, B => halt_i, C =>
                           ID_EXE_i(123), D => n160, Z => n125);
   U51 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_13_port, B => halt_i, C =>
                           ID_EXE_i(124), D => n160, Z => n126);
   U52 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_14_port, B => halt_i, C =>
                           ID_EXE_i(125), D => n160, Z => n127);
   U53 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_15_port, B => halt_i, C =>
                           ID_EXE_i(126), D => n160, Z => n128);
   U54 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_16_port, B => halt_i, C =>
                           ID_EXE_i(127), D => n160, Z => n129);
   U55 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_17_port, B => halt_i, C =>
                           ID_EXE_i(128), D => n160, Z => n130);
   U56 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_18_port, B => halt_i, C =>
                           ID_EXE_i(129), D => n160, Z => n131);
   U57 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_19_port, B => halt_i, C =>
                           ID_EXE_i(130), D => n160, Z => n132);
   U58 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_20_port, B => halt_i, C =>
                           ID_EXE_i(131), D => n160, Z => n133);
   U59 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_21_port, B => halt_i, C =>
                           ID_EXE_i(132), D => n161, Z => n134);
   U60 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_22_port, B => halt_i, C =>
                           ID_EXE_i(133), D => n161, Z => n135);
   U61 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_23_port, B => halt_i, C =>
                           ID_EXE_i(134), D => n161, Z => n136);
   U62 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_24_port, B => halt_i, C =>
                           ID_EXE_i(135), D => n161, Z => n137);
   U63 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_25_port, B => halt_i, C =>
                           ID_EXE_i(136), D => n161, Z => n138);
   U64 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_26_port, B => halt_i, C =>
                           ID_EXE_i(137), D => n161, Z => n139);
   U65 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_27_port, B => halt_i, C =>
                           ID_EXE_i(138), D => n161, Z => n140);
   U66 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_28_port, B => halt_i, C =>
                           ID_EXE_i(139), D => n161, Z => n141);
   U67 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_29_port, B => halt_i, C =>
                           ID_EXE_i(140), D => n161, Z => n142);
   U68 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_30_port, B => halt_i, C =>
                           ID_EXE_i(141), D => n161, Z => n143);
   U69 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGA_31_port, B => halt_i, C =>
                           ID_EXE_i(142), D => n161, Z => n144);
   U70 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_0_port, B => halt_i, C => 
                           ID_EXE_i(79), D => n156, Z => n81);
   U71 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_1_port, B => halt_i, C => 
                           ID_EXE_i(80), D => n156, Z => n82);
   U72 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_2_port, B => halt_i, C => 
                           ID_EXE_i(81), D => n156, Z => n83);
   U73 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_3_port, B => halt_i, C => 
                           ID_EXE_i(82), D => n156, Z => n84);
   U74 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_4_port, B => halt_i, C => 
                           ID_EXE_i(83), D => n156, Z => n85);
   U75 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_5_port, B => halt_i, C => 
                           ID_EXE_i(84), D => n157, Z => n86);
   U76 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_6_port, B => halt_i, C => 
                           ID_EXE_i(85), D => n157, Z => n87);
   U77 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_7_port, B => halt_i, C => 
                           ID_EXE_i(86), D => n157, Z => n88);
   U78 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_8_port, B => halt_i, C => 
                           ID_EXE_i(87), D => n157, Z => n89);
   U79 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_9_port, B => halt_i, C => 
                           ID_EXE_i(88), D => n157, Z => n90);
   U80 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_11_port, B => halt_i, C =>
                           ID_EXE_i(90), D => n157, Z => n92);
   U81 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_12_port, B => halt_i, C =>
                           ID_EXE_i(91), D => n157, Z => n93);
   U82 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_13_port, B => halt_i, C =>
                           ID_EXE_i(92), D => n157, Z => n94);
   U83 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_14_port, B => halt_i, C =>
                           ID_EXE_i(93), D => n157, Z => n95);
   U84 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_15_port, B => halt_i, C =>
                           ID_EXE_i(94), D => n157, Z => n96);
   U85 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_16_port, B => halt_i, C =>
                           ID_EXE_i(95), D => n157, Z => n97);
   U86 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_17_port, B => halt_i, C =>
                           ID_EXE_i(96), D => n158, Z => n98);
   U87 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_18_port, B => halt_i, C =>
                           ID_EXE_i(97), D => n158, Z => n99);
   U88 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_19_port, B => halt_i, C =>
                           ID_EXE_i(98), D => n158, Z => n100);
   U89 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_20_port, B => halt_i, C =>
                           ID_EXE_i(99), D => n158, Z => n101);
   U90 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_21_port, B => halt_i, C =>
                           ID_EXE_i(100), D => n158, Z => n102);
   U91 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_22_port, B => halt_i, C =>
                           ID_EXE_i(101), D => n158, Z => n103);
   U92 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_23_port, B => halt_i, C =>
                           ID_EXE_i(102), D => n158, Z => n104);
   U93 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_24_port, B => halt_i, C =>
                           ID_EXE_i(103), D => n158, Z => n105);
   U94 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_25_port, B => halt_i, C =>
                           ID_EXE_i(104), D => n158, Z => n106);
   U95 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_26_port, B => halt_i, C =>
                           ID_EXE_i(105), D => n158, Z => n107);
   U96 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_27_port, B => halt_i, C =>
                           ID_EXE_i(106), D => n158, Z => n108);
   U97 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_28_port, B => halt_i, C =>
                           ID_EXE_i(107), D => n158, Z => n109);
   U98 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_29_port, B => halt_i, C =>
                           ID_EXE_i(108), D => n159, Z => n110);
   U99 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_30_port, B => halt_i, C =>
                           ID_EXE_i(109), D => n159, Z => n111);
   U100 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_31_port, B => halt_i, C 
                           => ID_EXE_i(110), D => n159, Z => n112);
   U101 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGB_10_port, B => halt_i, C 
                           => ID_EXE_i(89), D => n157, Z => n91);
   U102 : HS65_LH_AO22X9 port map( A => ID_EXE_o_ALUSRC_B_port, B => halt_i, C 
                           => ID_EXE_i(8), D => n150, Z => n10);
   U103 : HS65_LH_AO22X9 port map( A => ID_EXE_o_CALU_OP_0_port, B => halt_i, C
                           => ID_EXE_i(1), D => n150, Z => n3);
   U104 : HS65_LH_AO22X9 port map( A => ID_EXE_o_CALU_OP_2_port, B => halt_i, C
                           => ID_EXE_i(3), D => n150, Z => n5);
   U105 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RT_0_port, B => halt_i, C => 
                           ID_EXE_i(14), D => n151, Z => n16);
   U106 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RS_0_port, B => halt_i, C => 
                           ID_EXE_i(19), D => n151, Z => n21);
   U107 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RT_1_port, B => halt_i, C => 
                           ID_EXE_i(15), D => n151, Z => n17);
   U108 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RT_2_port, B => halt_i, C => 
                           ID_EXE_i(16), D => n151, Z => n18);
   U109 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RT_3_port, B => halt_i, C => 
                           ID_EXE_i(17), D => n151, Z => n19);
   U110 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RS_1_port, B => halt_i, C => 
                           ID_EXE_i(20), D => n151, Z => n22);
   U111 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RS_2_port, B => halt_i, C => 
                           ID_EXE_i(21), D => n151, Z => n23);
   U112 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RS_3_port, B => halt_i, C => 
                           ID_EXE_i(22), D => n151, Z => n24);
   U113 : HS65_LH_AO22X9 port map( A => ID_EXE_o_REGWRITE_port, B => halt_i, C 
                           => ID_EXE_i(6), D => n150, Z => n8);
   U114 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RT_4_port, B => halt_i, C => 
                           ID_EXE_i(18), D => n151, Z => n20);
   U115 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RS_4_port, B => halt_i, C => 
                           ID_EXE_i(23), D => n151, Z => n25);
   U116 : HS65_LH_AO22X9 port map( A => ID_EXE_o_MEMWEN_N_port, B => halt_i, C 
                           => ID_EXE_i(5), D => n150, Z => n7);
   U117 : HS65_LH_AO22X9 port map( A => ID_EXE_o_CALU_OP_1_port, B => halt_i, C
                           => ID_EXE_i(2), D => n150, Z => n4);
   U118 : HS65_LH_AO22X9 port map( A => halt_i, B => ID_EXE_o_REGDST_port, C =>
                           ID_EXE_i(0), D => n150, Z => n2);
   U119 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RD_4_port, B => halt_i, C => 
                           ID_EXE_i(13), D => n151, Z => n15);
   U120 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_15_port, B => 
                           halt_i, C => ID_EXE_i(51), D => n154, Z => n53);
   U121 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_16_port, B => 
                           halt_i, C => ID_EXE_i(52), D => n154, Z => n54);
   U122 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_17_port, B => 
                           halt_i, C => ID_EXE_i(53), D => n154, Z => n55);
   U123 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_18_port, B => 
                           halt_i, C => ID_EXE_i(54), D => n154, Z => n56);
   U124 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_19_port, B => 
                           halt_i, C => ID_EXE_i(55), D => n154, Z => n57);
   U125 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_20_port, B => 
                           halt_i, C => ID_EXE_i(56), D => n154, Z => n58);
   U126 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_21_port, B => 
                           halt_i, C => ID_EXE_i(57), D => n154, Z => n59);
   U127 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_22_port, B => 
                           halt_i, C => ID_EXE_i(58), D => n154, Z => n60);
   U128 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_23_port, B => 
                           halt_i, C => ID_EXE_i(59), D => n154, Z => n61);
   U129 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_24_port, B => 
                           halt_i, C => ID_EXE_i(60), D => n155, Z => n62);
   U130 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_25_port, B => 
                           halt_i, C => ID_EXE_i(61), D => n155, Z => n63);
   U131 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_26_port, B => 
                           halt_i, C => ID_EXE_i(62), D => n155, Z => n64);
   U132 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_27_port, B => 
                           halt_i, C => ID_EXE_i(63), D => n155, Z => n65);
   U133 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_28_port, B => 
                           halt_i, C => ID_EXE_i(64), D => n155, Z => n66);
   U134 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_29_port, B => 
                           halt_i, C => ID_EXE_i(65), D => n155, Z => n67);
   U135 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_30_port, B => 
                           halt_i, C => ID_EXE_i(66), D => n155, Z => n68);
   U136 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_31_port, B => 
                           halt_i, C => ID_EXE_i(67), D => n155, Z => n69);
   U137 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RD_0_port, B => halt_i, C => 
                           ID_EXE_i(9), D => n150, Z => n11);
   U138 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RD_1_port, B => halt_i, C => 
                           ID_EXE_i(10), D => n150, Z => n12);
   U139 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RD_2_port, B => halt_i, C => 
                           ID_EXE_i(11), D => n150, Z => n13);
   U140 : HS65_LH_AO22X9 port map( A => ID_EXE_o_RD_3_port, B => halt_i, C => 
                           ID_EXE_i(12), D => n151, Z => n14);
   U141 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_0_port, B => 
                           halt_i, C => ID_EXE_i(36), D => n153, Z => n38);
   U142 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_1_port, B => 
                           halt_i, C => ID_EXE_i(37), D => n153, Z => n39);
   U143 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_2_port, B => 
                           halt_i, C => ID_EXE_i(38), D => n153, Z => n40);
   U144 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_3_port, B => 
                           halt_i, C => ID_EXE_i(39), D => n153, Z => n41);
   U145 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_4_port, B => 
                           halt_i, C => ID_EXE_i(40), D => n153, Z => n42);
   U146 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_5_port, B => 
                           halt_i, C => ID_EXE_i(41), D => n153, Z => n43);
   U147 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_6_port, B => 
                           halt_i, C => ID_EXE_i(42), D => n153, Z => n44);
   U148 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_7_port, B => 
                           halt_i, C => ID_EXE_i(43), D => n153, Z => n45);
   U149 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_8_port, B => 
                           halt_i, C => ID_EXE_i(44), D => n153, Z => n46);
   U150 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_9_port, B => 
                           halt_i, C => ID_EXE_i(45), D => n153, Z => n47);
   U151 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_10_port, B => 
                           halt_i, C => ID_EXE_i(46), D => n153, Z => n48);
   U152 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_11_port, B => 
                           halt_i, C => ID_EXE_i(47), D => n153, Z => n49);
   U153 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_12_port, B => 
                           halt_i, C => ID_EXE_i(48), D => n154, Z => n50);
   U154 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_13_port, B => 
                           halt_i, C => ID_EXE_i(49), D => n154, Z => n51);
   U155 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SIGN_EXTEND_14_port, B => 
                           halt_i, C => ID_EXE_i(50), D => n154, Z => n52);
   U156 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_0_port, B => halt_i, C 
                           => ID_EXE_i(68), D => n155, Z => n70);
   U157 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_1_port, B => halt_i, C 
                           => ID_EXE_i(69), D => n155, Z => n71);
   U158 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_2_port, B => halt_i, C 
                           => ID_EXE_i(70), D => n155, Z => n72);
   U159 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_3_port, B => halt_i, C 
                           => ID_EXE_i(71), D => n155, Z => n73);
   U160 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_4_port, B => halt_i, C 
                           => ID_EXE_i(72), D => n156, Z => n74);
   U161 : HS65_LH_AO22X9 port map( A => ID_EXE_o_FUNCT_5_port, B => halt_i, C 
                           => ID_EXE_i(73), D => n156, Z => n75);
   U162 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SHAMT_0_port, B => halt_i, C 
                           => ID_EXE_i(74), D => n156, Z => n76);
   U163 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SHAMT_1_port, B => halt_i, C 
                           => ID_EXE_i(75), D => n156, Z => n77);
   U164 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SHAMT_2_port, B => halt_i, C 
                           => ID_EXE_i(76), D => n156, Z => n78);
   U165 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SHAMT_3_port, B => halt_i, C 
                           => ID_EXE_i(77), D => n156, Z => n79);
   U166 : HS65_LH_AO22X9 port map( A => ID_EXE_o_SHAMT_4_port, B => halt_i, C 
                           => ID_EXE_i(78), D => n156, Z => n80);
   U167 : HS65_LH_AO22X9 port map( A => ID_EXE_o_MEMTOREG_port, B => halt_i, C 
                           => ID_EXE_i(7), D => n150, Z => n9);
   U168 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_1_port, B => halt_i, 
                           C => ID_EXE_i(25), D => n152, Z => n27);
   U169 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_2_port, B => halt_i, 
                           C => ID_EXE_i(26), D => n152, Z => n28);
   U170 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_3_port, B => halt_i, 
                           C => ID_EXE_i(27), D => n152, Z => n29);
   U171 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_4_port, B => halt_i, 
                           C => ID_EXE_i(28), D => n152, Z => n30);
   U172 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_5_port, B => halt_i, 
                           C => ID_EXE_i(29), D => n152, Z => n31);
   U173 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_6_port, B => halt_i, 
                           C => ID_EXE_i(30), D => n152, Z => n32);
   U174 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_7_port, B => halt_i, 
                           C => ID_EXE_i(31), D => n152, Z => n33);
   U175 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_8_port, B => halt_i, 
                           C => ID_EXE_i(32), D => n152, Z => n34);
   U176 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_9_port, B => halt_i, 
                           C => ID_EXE_i(33), D => n152, Z => n35);
   U177 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_10_port, B => halt_i,
                           C => ID_EXE_i(34), D => n152, Z => n36);
   U178 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_11_port, B => halt_i,
                           C => ID_EXE_i(35), D => n152, Z => n37);
   U179 : HS65_LH_AO22X9 port map( A => ID_EXE_o_PC_PLUS1_0_port, B => halt_i, 
                           C => ID_EXE_i(24), D => n152, Z => n26);
   U180 : HS65_LH_AO22X9 port map( A => ID_EXE_o_CALU_OP_3_port, B => halt_i, C
                           => ID_EXE_i(4), D => n150, Z => n6);
   U181 : HS65_LH_IVX9 port map( A => halt_i, Z => n180);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity id_top is

   port( clk, rst_n : in std_logic;  id_top_i : in std_logic_vector (71 downto 
         0);  id_top_o : out std_logic_vector (127 downto 0));

end id_top;

architecture SYN_Behavioral of id_top is

   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component regfile
      port( clk, rst_n : in std_logic;  regfile_i : in std_logic_vector (49 
            downto 0);  regfile_o : out std_logic_vector (63 downto 0));
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96 : std_logic;

begin
   
   regfile_inst : regfile port map( clk => clk, rst_n => rst_n, regfile_i(49) 
                           => id_top_i(65), regfile_i(48) => id_top_i(64), 
                           regfile_i(47) => id_top_i(63), regfile_i(46) => 
                           id_top_i(62), regfile_i(45) => id_top_i(61), 
                           regfile_i(44) => id_top_i(60), regfile_i(43) => 
                           id_top_i(59), regfile_i(42) => id_top_i(58), 
                           regfile_i(41) => id_top_i(57), regfile_i(40) => 
                           id_top_i(56), regfile_i(39) => id_top_i(4), 
                           regfile_i(38) => id_top_i(3), regfile_i(37) => 
                           id_top_i(2), regfile_i(36) => id_top_i(1), 
                           regfile_i(35) => id_top_i(0), regfile_i(34) => n96, 
                           regfile_i(33) => n95, regfile_i(32) => n94, 
                           regfile_i(31) => n93, regfile_i(30) => n92, 
                           regfile_i(29) => n91, regfile_i(28) => n90, 
                           regfile_i(27) => n89, regfile_i(26) => n88, 
                           regfile_i(25) => n87, regfile_i(24) => n86, 
                           regfile_i(23) => n85, regfile_i(22) => n84, 
                           regfile_i(21) => n83, regfile_i(20) => n82, 
                           regfile_i(19) => n81, regfile_i(18) => n80, 
                           regfile_i(17) => n79, regfile_i(16) => n78, 
                           regfile_i(15) => n77, regfile_i(14) => n76, 
                           regfile_i(13) => n75, regfile_i(12) => n74, 
                           regfile_i(11) => n73, regfile_i(10) => n72, 
                           regfile_i(9) => n71, regfile_i(8) => n70, 
                           regfile_i(7) => n69, regfile_i(6) => n68, 
                           regfile_i(5) => n67, regfile_i(4) => n66, 
                           regfile_i(3) => n65, regfile_i(2) => id_top_i(7), 
                           regfile_i(1) => id_top_i(6), regfile_i(0) => 
                           id_top_i(5), regfile_o(63) => id_top_o(127), 
                           regfile_o(62) => id_top_o(126), regfile_o(61) => 
                           id_top_o(125), regfile_o(60) => id_top_o(124), 
                           regfile_o(59) => id_top_o(123), regfile_o(58) => 
                           id_top_o(122), regfile_o(57) => id_top_o(121), 
                           regfile_o(56) => id_top_o(120), regfile_o(55) => 
                           id_top_o(119), regfile_o(54) => id_top_o(118), 
                           regfile_o(53) => id_top_o(117), regfile_o(52) => 
                           id_top_o(116), regfile_o(51) => id_top_o(115), 
                           regfile_o(50) => id_top_o(114), regfile_o(49) => 
                           id_top_o(113), regfile_o(48) => id_top_o(112), 
                           regfile_o(47) => id_top_o(111), regfile_o(46) => 
                           id_top_o(110), regfile_o(45) => id_top_o(109), 
                           regfile_o(44) => id_top_o(108), regfile_o(43) => 
                           id_top_o(107), regfile_o(42) => id_top_o(106), 
                           regfile_o(41) => id_top_o(105), regfile_o(40) => 
                           id_top_o(104), regfile_o(39) => id_top_o(103), 
                           regfile_o(38) => id_top_o(102), regfile_o(37) => 
                           id_top_o(101), regfile_o(36) => id_top_o(100), 
                           regfile_o(35) => id_top_o(99), regfile_o(34) => 
                           id_top_o(98), regfile_o(33) => id_top_o(97), 
                           regfile_o(32) => id_top_o(96), regfile_o(31) => 
                           id_top_o(95), regfile_o(30) => id_top_o(94), 
                           regfile_o(29) => id_top_o(93), regfile_o(28) => 
                           id_top_o(92), regfile_o(27) => id_top_o(91), 
                           regfile_o(26) => id_top_o(90), regfile_o(25) => 
                           id_top_o(89), regfile_o(24) => id_top_o(88), 
                           regfile_o(23) => id_top_o(87), regfile_o(22) => 
                           id_top_o(86), regfile_o(21) => id_top_o(85), 
                           regfile_o(20) => id_top_o(84), regfile_o(19) => 
                           id_top_o(83), regfile_o(18) => id_top_o(82), 
                           regfile_o(17) => id_top_o(81), regfile_o(16) => 
                           id_top_o(80), regfile_o(15) => id_top_o(79), 
                           regfile_o(14) => id_top_o(78), regfile_o(13) => 
                           id_top_o(77), regfile_o(12) => id_top_o(76), 
                           regfile_o(11) => id_top_o(75), regfile_o(10) => 
                           id_top_o(74), regfile_o(9) => id_top_o(73), 
                           regfile_o(8) => id_top_o(72), regfile_o(7) => 
                           id_top_o(71), regfile_o(6) => id_top_o(70), 
                           regfile_o(5) => id_top_o(69), regfile_o(4) => 
                           id_top_o(68), regfile_o(3) => id_top_o(67), 
                           regfile_o(2) => id_top_o(66), regfile_o(1) => 
                           id_top_o(65), regfile_o(0) => id_top_o(64));
   U1 : HS65_LH_BFX9 port map( A => id_top_i(8), Z => n65);
   U2 : HS65_LH_BFX9 port map( A => id_top_i(9), Z => n66);
   U3 : HS65_LH_BFX9 port map( A => id_top_i(10), Z => n67);
   U4 : HS65_LH_BFX9 port map( A => id_top_i(11), Z => n68);
   U5 : HS65_LH_BFX9 port map( A => id_top_i(12), Z => n69);
   U6 : HS65_LH_BFX9 port map( A => id_top_i(13), Z => n70);
   U7 : HS65_LH_BFX9 port map( A => id_top_i(14), Z => n71);
   U8 : HS65_LH_BFX9 port map( A => id_top_i(15), Z => n72);
   U9 : HS65_LH_BFX9 port map( A => id_top_i(16), Z => n73);
   U10 : HS65_LH_BFX9 port map( A => id_top_i(17), Z => n74);
   U11 : HS65_LH_BFX9 port map( A => id_top_i(18), Z => n75);
   U12 : HS65_LH_BFX9 port map( A => id_top_i(19), Z => n76);
   U13 : HS65_LH_BFX9 port map( A => id_top_i(20), Z => n77);
   U14 : HS65_LH_BFX9 port map( A => id_top_i(21), Z => n78);
   U15 : HS65_LH_BFX9 port map( A => id_top_i(22), Z => n79);
   U16 : HS65_LH_BFX9 port map( A => id_top_i(23), Z => n80);
   U17 : HS65_LH_BFX9 port map( A => id_top_i(24), Z => n81);
   U18 : HS65_LH_BFX9 port map( A => id_top_i(25), Z => n82);
   U19 : HS65_LH_BFX9 port map( A => id_top_i(26), Z => n83);
   U20 : HS65_LH_BFX9 port map( A => id_top_i(27), Z => n84);
   U21 : HS65_LH_BFX9 port map( A => id_top_i(28), Z => n85);
   U22 : HS65_LH_BFX9 port map( A => id_top_i(29), Z => n86);
   U23 : HS65_LH_BFX9 port map( A => id_top_i(30), Z => n87);
   U24 : HS65_LH_BFX9 port map( A => id_top_i(31), Z => n88);
   U25 : HS65_LH_BFX9 port map( A => id_top_i(32), Z => n89);
   U26 : HS65_LH_BFX9 port map( A => id_top_i(33), Z => n90);
   U27 : HS65_LH_BFX9 port map( A => id_top_i(34), Z => n91);
   U28 : HS65_LH_BFX9 port map( A => id_top_i(35), Z => n92);
   U29 : HS65_LH_BFX9 port map( A => id_top_i(36), Z => n93);
   U30 : HS65_LH_BFX9 port map( A => id_top_i(37), Z => n94);
   U31 : HS65_LH_BFX9 port map( A => id_top_i(38), Z => n95);
   U32 : HS65_LH_BFX9 port map( A => id_top_i(39), Z => n96);
   U33 : HS65_LH_BFX9 port map( A => id_top_i(51), Z => id_top_o(43));
   U34 : HS65_LH_BFX9 port map( A => id_top_i(52), Z => id_top_o(44));
   U35 : HS65_LH_BFX9 port map( A => id_top_i(53), Z => id_top_o(45));
   U36 : HS65_LH_BFX9 port map( A => id_top_i(54), Z => id_top_o(46));
   U37 : HS65_LH_BFX9 port map( A => id_top_i(40), Z => id_top_o(0));
   U38 : HS65_LH_BFX9 port map( A => id_top_i(41), Z => id_top_o(1));
   U39 : HS65_LH_BFX9 port map( A => id_top_i(42), Z => id_top_o(2));
   U40 : HS65_LH_BFX9 port map( A => id_top_i(43), Z => id_top_o(3));
   U41 : HS65_LH_BFX9 port map( A => id_top_i(44), Z => id_top_o(4));
   U42 : HS65_LH_BFX9 port map( A => id_top_i(45), Z => id_top_o(5));
   U43 : HS65_LH_BFX9 port map( A => id_top_i(46), Z => id_top_o(6));
   U44 : HS65_LH_BFX9 port map( A => id_top_i(47), Z => id_top_o(7));
   U45 : HS65_LH_BFX9 port map( A => id_top_i(48), Z => id_top_o(8));
   U46 : HS65_LH_BFX9 port map( A => id_top_i(49), Z => id_top_o(9));
   U47 : HS65_LH_BFX9 port map( A => id_top_i(50), Z => id_top_o(10));
   U48 : HS65_LH_BFX9 port map( A => id_top_i(51), Z => id_top_o(11));
   U49 : HS65_LH_BFX9 port map( A => id_top_i(52), Z => id_top_o(12));
   U50 : HS65_LH_BFX9 port map( A => id_top_i(53), Z => id_top_o(13));
   U51 : HS65_LH_BFX9 port map( A => id_top_i(54), Z => id_top_o(14));
   U52 : HS65_LH_BFX9 port map( A => id_top_i(40), Z => id_top_o(32));
   U53 : HS65_LH_BFX9 port map( A => id_top_i(41), Z => id_top_o(33));
   U54 : HS65_LH_BFX9 port map( A => id_top_i(42), Z => id_top_o(34));
   U55 : HS65_LH_BFX9 port map( A => id_top_i(43), Z => id_top_o(35));
   U56 : HS65_LH_BFX9 port map( A => id_top_i(44), Z => id_top_o(36));
   U57 : HS65_LH_BFX9 port map( A => id_top_i(45), Z => id_top_o(37));
   U58 : HS65_LH_BFX9 port map( A => id_top_i(46), Z => id_top_o(38));
   U59 : HS65_LH_BFX9 port map( A => id_top_i(47), Z => id_top_o(39));
   U60 : HS65_LH_BFX9 port map( A => id_top_i(48), Z => id_top_o(40));
   U61 : HS65_LH_BFX9 port map( A => id_top_i(49), Z => id_top_o(41));
   U62 : HS65_LH_BFX9 port map( A => id_top_i(50), Z => id_top_o(42));
   U63 : HS65_LH_BFX9 port map( A => id_top_i(71), Z => id_top_o(63));
   U64 : HS65_LH_BFX9 port map( A => id_top_i(70), Z => id_top_o(62));
   U65 : HS65_LH_BFX9 port map( A => id_top_i(69), Z => id_top_o(61));
   U66 : HS65_LH_BFX9 port map( A => id_top_i(68), Z => id_top_o(60));
   U67 : HS65_LH_BFX9 port map( A => id_top_i(67), Z => id_top_o(59));
   U68 : HS65_LH_BFX9 port map( A => id_top_i(66), Z => id_top_o(58));
   U69 : HS65_LH_BFX9 port map( A => id_top_i(65), Z => id_top_o(57));
   U70 : HS65_LH_BFX9 port map( A => id_top_i(64), Z => id_top_o(56));
   U71 : HS65_LH_BFX9 port map( A => id_top_i(63), Z => id_top_o(55));
   U72 : HS65_LH_BFX9 port map( A => id_top_i(62), Z => id_top_o(54));
   U73 : HS65_LH_BFX9 port map( A => id_top_i(61), Z => id_top_o(53));
   U74 : HS65_LH_BFX9 port map( A => id_top_i(60), Z => id_top_o(52));
   U75 : HS65_LH_BFX9 port map( A => id_top_i(59), Z => id_top_o(51));
   U76 : HS65_LH_BFX9 port map( A => id_top_i(58), Z => id_top_o(50));
   U77 : HS65_LH_BFX9 port map( A => id_top_i(57), Z => id_top_o(49));
   U78 : HS65_LH_BFX9 port map( A => id_top_i(56), Z => id_top_o(48));
   U79 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(16));
   U80 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(17));
   U81 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(18));
   U82 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(19));
   U83 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(20));
   U84 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(21));
   U85 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(22));
   U86 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(23));
   U87 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(24));
   U88 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(25));
   U89 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(26));
   U90 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(27));
   U91 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(28));
   U92 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(29));
   U93 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(30));
   U94 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(31));
   U95 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(47));
   U96 : HS65_LH_BFX9 port map( A => id_top_i(55), Z => id_top_o(15));

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity if_id is

   port( clk, rst_n, halt_i : in std_logic;  IF_ID_i : in std_logic_vector (11 
         downto 0);  IF_ID_o : out std_logic_vector (11 downto 0));

end if_id;

architecture SYN_Behavioral of if_id is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_DFPRQX9
      port( D, CP, RN : in std_logic;  Q : out std_logic);
   end component;
   
   signal IF_ID_o_PC_PLUS1_11_port, IF_ID_o_PC_PLUS1_10_port, 
      IF_ID_o_PC_PLUS1_9_port, IF_ID_o_PC_PLUS1_8_port, IF_ID_o_PC_PLUS1_7_port
      , IF_ID_o_PC_PLUS1_6_port, IF_ID_o_PC_PLUS1_5_port, 
      IF_ID_o_PC_PLUS1_4_port, IF_ID_o_PC_PLUS1_3_port, IF_ID_o_PC_PLUS1_2_port
      , IF_ID_o_PC_PLUS1_1_port, IF_ID_o_PC_PLUS1_0_port, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n1 : std_logic;

begin
   IF_ID_o <= ( IF_ID_o_PC_PLUS1_11_port, IF_ID_o_PC_PLUS1_10_port, 
      IF_ID_o_PC_PLUS1_9_port, IF_ID_o_PC_PLUS1_8_port, IF_ID_o_PC_PLUS1_7_port
      , IF_ID_o_PC_PLUS1_6_port, IF_ID_o_PC_PLUS1_5_port, 
      IF_ID_o_PC_PLUS1_4_port, IF_ID_o_PC_PLUS1_3_port, IF_ID_o_PC_PLUS1_2_port
      , IF_ID_o_PC_PLUS1_1_port, IF_ID_o_PC_PLUS1_0_port );
   
   if_id_c_reg_PC_PLUS1_11_inst : HS65_LH_DFPRQX9 port map( D => n13, CP => clk
                           , RN => rst_n, Q => IF_ID_o_PC_PLUS1_11_port);
   if_id_c_reg_PC_PLUS1_10_inst : HS65_LH_DFPRQX9 port map( D => n12, CP => clk
                           , RN => rst_n, Q => IF_ID_o_PC_PLUS1_10_port);
   if_id_c_reg_PC_PLUS1_9_inst : HS65_LH_DFPRQX9 port map( D => n11, CP => clk,
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_9_port);
   if_id_c_reg_PC_PLUS1_8_inst : HS65_LH_DFPRQX9 port map( D => n10, CP => clk,
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_8_port);
   if_id_c_reg_PC_PLUS1_7_inst : HS65_LH_DFPRQX9 port map( D => n9, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_7_port);
   if_id_c_reg_PC_PLUS1_6_inst : HS65_LH_DFPRQX9 port map( D => n8, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_6_port);
   if_id_c_reg_PC_PLUS1_5_inst : HS65_LH_DFPRQX9 port map( D => n7, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_5_port);
   if_id_c_reg_PC_PLUS1_4_inst : HS65_LH_DFPRQX9 port map( D => n6, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_4_port);
   if_id_c_reg_PC_PLUS1_3_inst : HS65_LH_DFPRQX9 port map( D => n5, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_3_port);
   if_id_c_reg_PC_PLUS1_2_inst : HS65_LH_DFPRQX9 port map( D => n4, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_2_port);
   if_id_c_reg_PC_PLUS1_1_inst : HS65_LH_DFPRQX9 port map( D => n3, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_1_port);
   if_id_c_reg_PC_PLUS1_0_inst : HS65_LH_DFPRQX9 port map( D => n2, CP => clk, 
                           RN => rst_n, Q => IF_ID_o_PC_PLUS1_0_port);
   U2 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_11_port, B => halt_i, C 
                           => IF_ID_i(11), D => n1, Z => n13);
   U3 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_7_port, B => halt_i, C 
                           => IF_ID_i(7), D => n1, Z => n9);
   U4 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_8_port, B => halt_i, C 
                           => IF_ID_i(8), D => n1, Z => n10);
   U5 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_9_port, B => halt_i, C 
                           => IF_ID_i(9), D => n1, Z => n11);
   U6 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_10_port, B => halt_i, C 
                           => IF_ID_i(10), D => n1, Z => n12);
   U7 : HS65_LH_AO22X9 port map( A => halt_i, B => IF_ID_o_PC_PLUS1_0_port, C 
                           => IF_ID_i(0), D => n1, Z => n2);
   U8 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_1_port, B => halt_i, C 
                           => IF_ID_i(1), D => n1, Z => n3);
   U9 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_2_port, B => halt_i, C 
                           => IF_ID_i(2), D => n1, Z => n4);
   U10 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_3_port, B => halt_i, C 
                           => IF_ID_i(3), D => n1, Z => n5);
   U11 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_4_port, B => halt_i, C 
                           => IF_ID_i(4), D => n1, Z => n6);
   U12 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_5_port, B => halt_i, C 
                           => IF_ID_i(5), D => n1, Z => n7);
   U13 : HS65_LH_AO22X9 port map( A => IF_ID_o_PC_PLUS1_6_port, B => halt_i, C 
                           => IF_ID_i(6), D => n1, Z => n8);
   U14 : HS65_LH_IVX9 port map( A => halt_i, Z => n1);

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity if_top is

   port( clk, rst_n : in std_logic;  if_top_i : in std_logic_vector (13 downto 
         0);  if_top_o : out std_logic_vector (23 downto 0));

end if_top;

architecture SYN_behavioral of if_top is

   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component if_top_DW01_inc_0
      port( A : in std_logic_vector (11 downto 0);  SUM : out std_logic_vector 
            (11 downto 0));
   end component;
   
   component pc
      port( clk, rst_n, halt_i : in std_logic;  npc_i : in std_logic_vector (11
            downto 0);  pc_o : out std_logic_vector (11 downto 0));
   end component;
   
   signal if_top_o_IMEM_ADDR_11_port, if_top_o_IMEM_ADDR_10_port, 
      if_top_o_IMEM_ADDR_9_port, if_top_o_IMEM_ADDR_8_port, 
      if_top_o_IMEM_ADDR_7_port, if_top_o_IMEM_ADDR_6_port, 
      if_top_o_IMEM_ADDR_5_port, if_top_o_IMEM_ADDR_4_port, 
      if_top_o_IMEM_ADDR_3_port, if_top_o_IMEM_ADDR_2_port, 
      if_top_o_IMEM_ADDR_1_port, if_top_o_IMEM_ADDR_0_port, 
      if_top_o_PC_PLUS1_11_port, if_top_o_PC_PLUS1_10_port, 
      if_top_o_PC_PLUS1_9_port, if_top_o_PC_PLUS1_8_port, 
      if_top_o_PC_PLUS1_7_port, if_top_o_PC_PLUS1_6_port, 
      if_top_o_PC_PLUS1_5_port, if_top_o_PC_PLUS1_4_port, 
      if_top_o_PC_PLUS1_3_port, if_top_o_PC_PLUS1_2_port, 
      if_top_o_PC_PLUS1_1_port, if_top_o_PC_PLUS1_0_port, s_npc_11_port, 
      s_npc_10_port, s_npc_9_port, s_npc_8_port, s_npc_7_port, s_npc_6_port, 
      s_npc_5_port, s_npc_4_port, s_npc_3_port, s_npc_2_port, s_npc_1_port, 
      s_npc_0_port, n1 : std_logic;

begin
   if_top_o <= ( if_top_o_IMEM_ADDR_11_port, if_top_o_IMEM_ADDR_10_port, 
      if_top_o_IMEM_ADDR_9_port, if_top_o_IMEM_ADDR_8_port, 
      if_top_o_IMEM_ADDR_7_port, if_top_o_IMEM_ADDR_6_port, 
      if_top_o_IMEM_ADDR_5_port, if_top_o_IMEM_ADDR_4_port, 
      if_top_o_IMEM_ADDR_3_port, if_top_o_IMEM_ADDR_2_port, 
      if_top_o_IMEM_ADDR_1_port, if_top_o_IMEM_ADDR_0_port, 
      if_top_o_PC_PLUS1_11_port, if_top_o_PC_PLUS1_10_port, 
      if_top_o_PC_PLUS1_9_port, if_top_o_PC_PLUS1_8_port, 
      if_top_o_PC_PLUS1_7_port, if_top_o_PC_PLUS1_6_port, 
      if_top_o_PC_PLUS1_5_port, if_top_o_PC_PLUS1_4_port, 
      if_top_o_PC_PLUS1_3_port, if_top_o_PC_PLUS1_2_port, 
      if_top_o_PC_PLUS1_1_port, if_top_o_PC_PLUS1_0_port );
   
   pc_inst : pc port map( clk => clk, rst_n => rst_n, halt_i => if_top_i(13), 
                           npc_i(11) => s_npc_11_port, npc_i(10) => 
                           s_npc_10_port, npc_i(9) => s_npc_9_port, npc_i(8) =>
                           s_npc_8_port, npc_i(7) => s_npc_7_port, npc_i(6) => 
                           s_npc_6_port, npc_i(5) => s_npc_5_port, npc_i(4) => 
                           s_npc_4_port, npc_i(3) => s_npc_3_port, npc_i(2) => 
                           s_npc_2_port, npc_i(1) => s_npc_1_port, npc_i(0) => 
                           s_npc_0_port, pc_o(11) => if_top_o_IMEM_ADDR_11_port
                           , pc_o(10) => if_top_o_IMEM_ADDR_10_port, pc_o(9) =>
                           if_top_o_IMEM_ADDR_9_port, pc_o(8) => 
                           if_top_o_IMEM_ADDR_8_port, pc_o(7) => 
                           if_top_o_IMEM_ADDR_7_port, pc_o(6) => 
                           if_top_o_IMEM_ADDR_6_port, pc_o(5) => 
                           if_top_o_IMEM_ADDR_5_port, pc_o(4) => 
                           if_top_o_IMEM_ADDR_4_port, pc_o(3) => 
                           if_top_o_IMEM_ADDR_3_port, pc_o(2) => 
                           if_top_o_IMEM_ADDR_2_port, pc_o(1) => 
                           if_top_o_IMEM_ADDR_1_port, pc_o(0) => 
                           if_top_o_IMEM_ADDR_0_port);
   add_37 : if_top_DW01_inc_0 port map( A(11) => if_top_o_IMEM_ADDR_11_port, 
                           A(10) => if_top_o_IMEM_ADDR_10_port, A(9) => 
                           if_top_o_IMEM_ADDR_9_port, A(8) => 
                           if_top_o_IMEM_ADDR_8_port, A(7) => 
                           if_top_o_IMEM_ADDR_7_port, A(6) => 
                           if_top_o_IMEM_ADDR_6_port, A(5) => 
                           if_top_o_IMEM_ADDR_5_port, A(4) => 
                           if_top_o_IMEM_ADDR_4_port, A(3) => 
                           if_top_o_IMEM_ADDR_3_port, A(2) => 
                           if_top_o_IMEM_ADDR_2_port, A(1) => 
                           if_top_o_IMEM_ADDR_1_port, A(0) => 
                           if_top_o_IMEM_ADDR_0_port, SUM(11) => 
                           if_top_o_PC_PLUS1_11_port, SUM(10) => 
                           if_top_o_PC_PLUS1_10_port, SUM(9) => 
                           if_top_o_PC_PLUS1_9_port, SUM(8) => 
                           if_top_o_PC_PLUS1_8_port, SUM(7) => 
                           if_top_o_PC_PLUS1_7_port, SUM(6) => 
                           if_top_o_PC_PLUS1_6_port, SUM(5) => 
                           if_top_o_PC_PLUS1_5_port, SUM(4) => 
                           if_top_o_PC_PLUS1_4_port, SUM(3) => 
                           if_top_o_PC_PLUS1_3_port, SUM(2) => 
                           if_top_o_PC_PLUS1_2_port, SUM(1) => 
                           if_top_o_PC_PLUS1_1_port, SUM(0) => 
                           if_top_o_PC_PLUS1_0_port);
   U2 : HS65_LH_IVX9 port map( A => if_top_i(0), Z => n1);
   U3 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_9_port, B => n1, C => 
                           if_top_i(0), D => if_top_i(10), Z => s_npc_9_port);
   U4 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_0_port, B => n1, C => 
                           if_top_i(1), D => if_top_i(0), Z => s_npc_0_port);
   U5 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_1_port, B => n1, C => 
                           if_top_i(2), D => if_top_i(0), Z => s_npc_1_port);
   U6 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_2_port, B => n1, C => 
                           if_top_i(3), D => if_top_i(0), Z => s_npc_2_port);
   U7 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_3_port, B => n1, C => 
                           if_top_i(4), D => if_top_i(0), Z => s_npc_3_port);
   U8 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_4_port, B => n1, C => 
                           if_top_i(5), D => if_top_i(0), Z => s_npc_4_port);
   U9 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_5_port, B => n1, C => 
                           if_top_i(6), D => if_top_i(0), Z => s_npc_5_port);
   U10 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_6_port, B => n1, C => 
                           if_top_i(7), D => if_top_i(0), Z => s_npc_6_port);
   U11 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_7_port, B => n1, C => 
                           if_top_i(8), D => if_top_i(0), Z => s_npc_7_port);
   U12 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_8_port, B => n1, C => 
                           if_top_i(9), D => if_top_i(0), Z => s_npc_8_port);
   U13 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_10_port, B => n1, C =>
                           if_top_i(11), D => if_top_i(0), Z => s_npc_10_port);
   U14 : HS65_LH_AO22X9 port map( A => if_top_o_PC_PLUS1_11_port, B => n1, C =>
                           if_top_i(12), D => if_top_i(0), Z => s_npc_11_port);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity controller is

   port( ctrl_i : in std_logic_vector (5 downto 0);  ctrl_o : out 
         std_logic_vector (9 downto 0));

end controller;

architecture SYN_behavioral of controller is

   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CB4I6X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_CBI4I1X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3X4
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND4ABX3
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR4ABX2
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI21X3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_OAI31X5
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR3AX2
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND3X5
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NAND2X7
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal ctrl_o_REGDST_port, ctrl_o_ALUSRC_B_port, ctrl_o_MEMTOREG_port, 
      ctrl_o_REGWRITE_port, ctrl_o_MEMWEN_N_port, ctrl_o_BRANCH_port, 
      ctrl_o_CALU_OP_2_port, ctrl_o_CALU_OP_1_port, ctrl_o_CALU_OP_0_port, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      ctrl_o_CALU_OP_3_port, n2, n3, n4, n5, n6, n7, n8, n24 : std_logic;

begin
   ctrl_o <= ( ctrl_o_REGDST_port, ctrl_o_ALUSRC_B_port, ctrl_o_MEMTOREG_port, 
      ctrl_o_REGWRITE_port, ctrl_o_MEMWEN_N_port, ctrl_o_BRANCH_port, 
      ctrl_o_CALU_OP_3_port, ctrl_o_CALU_OP_2_port, ctrl_o_CALU_OP_1_port, 
      ctrl_o_CALU_OP_0_port );
   
   U3 : HS65_LH_IVX9 port map( A => n2, Z => ctrl_o_CALU_OP_3_port);
   n2 <= '1';
   U5 : HS65_LH_OAI31X5 port map( A => n22, B => n14, C => n15, D => n8, Z => 
                           n21);
   U6 : HS65_LH_NOR2X6 port map( A => n24, B => n4, Z => n22);
   U7 : HS65_LH_NAND2X7 port map( A => n17, B => n8, Z => n10);
   U8 : HS65_LH_NAND2X7 port map( A => n19, B => n16, Z => n11);
   U9 : HS65_LH_IVX9 port map( A => n19, Z => n4);
   U10 : HS65_LH_NOR4ABX2 port map( A => n16, B => n5, C => n7, D => ctrl_i(2),
                           Z => n15);
   U11 : HS65_LH_NOR3AX2 port map( A => n23, B => ctrl_i(1), C => ctrl_i(2), Z 
                           => n14);
   U12 : HS65_LH_NOR3X4 port map( A => n7, B => ctrl_i(2), C => n5, Z => n19);
   U13 : HS65_LH_NAND3X5 port map( A => n23, B => ctrl_i(1), C => ctrl_i(2), Z 
                           => n12);
   U14 : HS65_LH_NOR4ABX2 port map( A => n16, B => n5, C => ctrl_i(1), D => 
                           ctrl_i(2), Z => n13);
   U15 : HS65_LH_NOR3X4 port map( A => n24, B => ctrl_i(3), C => n4, Z => n17);
   U16 : HS65_LH_NAND3X5 port map( A => n16, B => n7, C => ctrl_i(2), Z => n20)
                           ;
   U17 : HS65_LH_NOR3AX2 port map( A => ctrl_i(3), B => n5, C => ctrl_i(5), Z 
                           => n23);
   U18 : HS65_LH_NOR2X6 port map( A => ctrl_i(5), B => ctrl_i(3), Z => n16);
   U19 : HS65_LH_IVX9 port map( A => ctrl_i(4), Z => n8);
   U20 : HS65_LH_OAI21X3 port map( A => ctrl_i(4), B => n11, C => n6, Z => 
                           ctrl_o_CALU_OP_2_port);
   U21 : HS65_LH_IVX9 port map( A => ctrl_i(1), Z => n7);
   U22 : HS65_LH_IVX9 port map( A => ctrl_i(5), Z => n24);
   U23 : HS65_LH_IVX9 port map( A => ctrl_o_BRANCH_port, Z => n6);
   U24 : HS65_LH_NOR2X6 port map( A => n20, B => ctrl_i(4), Z => 
                           ctrl_o_BRANCH_port);
   U25 : HS65_LH_IVX9 port map( A => ctrl_i(0), Z => n5);
   U26 : HS65_LH_OAI21X3 port map( A => ctrl_i(4), B => n12, C => n21, Z => 
                           ctrl_o_ALUSRC_B_port);
   U27 : HS65_LH_OAI31X5 port map( A => n20, B => ctrl_i(4), C => n5, D => n21,
                           Z => ctrl_o_CALU_OP_0_port);
   U28 : HS65_LH_OAI21X3 port map( A => ctrl_i(4), B => n9, C => n10, Z => 
                           ctrl_o_REGWRITE_port);
   U29 : HS65_LH_NOR4ABX2 port map( A => n11, B => n12, C => n13, D => n14, Z 
                           => n9);
   U30 : HS65_LH_NAND4ABX3 port map( A => n17, B => ctrl_i(2), C => n8, D => 
                           n18, Z => ctrl_o_MEMWEN_N_port);
   U31 : HS65_LH_NOR3X4 port map( A => n5, B => n24, C => n7, Z => n18);
   U32 : HS65_LH_CBI4I1X5 port map( A => n3, B => n12, C => ctrl_i(4), D => n6,
                           Z => ctrl_o_CALU_OP_1_port);
   U33 : HS65_LH_IVX9 port map( A => n15, Z => n3);
   U34 : HS65_LH_CB4I6X9 port map( A => n13, B => n15, C => n8, D => 
                           ctrl_o_CALU_OP_2_port, Z => ctrl_o_REGDST_port);
   U35 : HS65_LH_IVX9 port map( A => n10, Z => ctrl_o_MEMTOREG_port);

end SYN_behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity mini_mips_pipeline is

   port( clk, rst_n : in std_logic;  mini_mips_i : in std_logic_vector (63 
         downto 0);  mini_mips_o : out std_logic_vector (56 downto 0));

end mini_mips_pipeline;

architecture SYN_Behavioral of mini_mips_pipeline is

   component HS65_LH_BFX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO222X4
      port( A, B, C, D, E, F : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AO22X9
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_NOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_IVX9
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LH_AND2X4
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HS65_LHS_XNOR2X6
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component mem_wb
      port( clk, rst_n, halt_i : in std_logic;  MEM_WB_i : in std_logic_vector 
            (38 downto 0);  MEM_WB_o : out std_logic_vector (38 downto 0));
   end component;
   
   component exe_mem
      port( clk, rst_n, halt_i : in std_logic;  EXE_MEM_i : in std_logic_vector
            (71 downto 0);  EXE_MEM_o : out std_logic_vector (71 downto 0));
   end component;
   
   component forwarding_unit
      port( forwarding_unit_i : in std_logic_vector (31 downto 0);  
            forwarding_unit_o : out std_logic_vector (5 downto 0));
   end component;
   
   component exe_top
      port( clk, rst_n : in std_logic;  exe_top_i : in std_logic_vector (134 
            downto 0);  exe_top_o : out std_logic_vector (81 downto 0));
   end component;
   
   component id_exe
      port( clk, rst_n, halt_i : in std_logic;  ID_EXE_i : in std_logic_vector 
            (142 downto 0);  ID_EXE_o : out std_logic_vector (142 downto 0));
   end component;
   
   component id_top
      port( clk, rst_n : in std_logic;  id_top_i : in std_logic_vector (71 
            downto 0);  id_top_o : out std_logic_vector (127 downto 0));
   end component;
   
   component if_id
      port( clk, rst_n, halt_i : in std_logic;  IF_ID_i : in std_logic_vector 
            (11 downto 0);  IF_ID_o : out std_logic_vector (11 downto 0));
   end component;
   
   component if_top
      port( clk, rst_n : in std_logic;  if_top_i : in std_logic_vector (13 
            downto 0);  if_top_o : out std_logic_vector (23 downto 0));
   end component;
   
   component controller
      port( ctrl_i : in std_logic_vector (5 downto 0);  ctrl_o : out 
            std_logic_vector (9 downto 0));
   end component;
   
   signal X_Logic0_port, mini_mips_o_DMEM_ADDR_11_port, 
      mini_mips_o_DMEM_ADDR_10_port, mini_mips_o_DMEM_ADDR_9_port, 
      mini_mips_o_DMEM_ADDR_8_port, mini_mips_o_DMEM_ADDR_7_port, 
      mini_mips_o_DMEM_ADDR_6_port, mini_mips_o_DMEM_ADDR_5_port, 
      mini_mips_o_DMEM_ADDR_4_port, mini_mips_o_DMEM_ADDR_3_port, 
      mini_mips_o_DMEM_ADDR_2_port, mini_mips_o_DMEM_ADDR_1_port, 
      mini_mips_o_DMEM_ADDR_0_port, mini_mips_o_DMEM_DATA_31_port, 
      mini_mips_o_DMEM_DATA_30_port, mini_mips_o_DMEM_DATA_29_port, 
      mini_mips_o_DMEM_DATA_28_port, mini_mips_o_DMEM_DATA_27_port, 
      mini_mips_o_DMEM_DATA_26_port, mini_mips_o_DMEM_DATA_25_port, 
      mini_mips_o_DMEM_DATA_24_port, mini_mips_o_DMEM_DATA_23_port, 
      mini_mips_o_DMEM_DATA_22_port, mini_mips_o_DMEM_DATA_21_port, 
      mini_mips_o_DMEM_DATA_20_port, mini_mips_o_DMEM_DATA_19_port, 
      mini_mips_o_DMEM_DATA_18_port, mini_mips_o_DMEM_DATA_17_port, 
      mini_mips_o_DMEM_DATA_16_port, mini_mips_o_DMEM_DATA_15_port, 
      mini_mips_o_DMEM_DATA_14_port, mini_mips_o_DMEM_DATA_13_port, 
      mini_mips_o_DMEM_DATA_12_port, mini_mips_o_DMEM_DATA_11_port, 
      mini_mips_o_DMEM_DATA_10_port, mini_mips_o_DMEM_DATA_9_port, 
      mini_mips_o_DMEM_DATA_8_port, mini_mips_o_DMEM_DATA_7_port, 
      mini_mips_o_DMEM_DATA_6_port, mini_mips_o_DMEM_DATA_5_port, 
      mini_mips_o_DMEM_DATA_4_port, mini_mips_o_DMEM_DATA_3_port, 
      mini_mips_o_DMEM_DATA_2_port, mini_mips_o_DMEM_DATA_1_port, 
      mini_mips_o_DMEM_DATA_0_port, mini_mips_o_IMEM_ADDR_11_port, 
      mini_mips_o_IMEM_ADDR_10_port, mini_mips_o_IMEM_ADDR_9_port, 
      mini_mips_o_IMEM_ADDR_8_port, mini_mips_o_IMEM_ADDR_7_port, 
      mini_mips_o_IMEM_ADDR_6_port, mini_mips_o_IMEM_ADDR_5_port, 
      mini_mips_o_IMEM_ADDR_4_port, mini_mips_o_IMEM_ADDR_3_port, 
      mini_mips_o_IMEM_ADDR_2_port, mini_mips_o_IMEM_ADDR_1_port, 
      mini_mips_o_IMEM_ADDR_0_port, mini_mips_o_DMEM_WEN_N_port, 
      s_id_out_pc_plus1_p_11_port, s_id_out_pc_plus1_p_10_port, 
      s_id_out_pc_plus1_p_9_port, s_id_out_pc_plus1_p_8_port, 
      s_id_out_pc_plus1_p_7_port, s_id_out_pc_plus1_p_6_port, 
      s_id_out_pc_plus1_p_5_port, s_id_out_pc_plus1_p_4_port, 
      s_id_out_pc_plus1_p_3_port, s_id_out_pc_plus1_p_2_port, 
      s_id_out_pc_plus1_p_1_port, s_id_out_pc_plus1_p_0_port, s_if_PCSrc, 
      s_exe_out_memtoReg_p, s_exe_out_regWrite_p, s_exe_out_memWen_n_p, 
      s_mem_out_memtoReg_p, s_mem_out_regWrite_p, s_mem_out_write_reg_p_4_port,
      s_mem_out_write_reg_p_3_port, s_mem_out_write_reg_p_2_port, 
      s_mem_out_write_reg_p_1_port, s_mem_out_write_reg_p_0_port, 
      s_mem_out_alu_res_p_31_port, s_mem_out_alu_res_p_30_port, 
      s_mem_out_alu_res_p_29_port, s_mem_out_alu_res_p_28_port, 
      s_mem_out_alu_res_p_27_port, s_mem_out_alu_res_p_26_port, 
      s_mem_out_alu_res_p_25_port, s_mem_out_alu_res_p_24_port, 
      s_mem_out_alu_res_p_23_port, s_mem_out_alu_res_p_22_port, 
      s_mem_out_alu_res_p_21_port, s_mem_out_alu_res_p_20_port, 
      s_mem_out_alu_res_p_19_port, s_mem_out_alu_res_p_18_port, 
      s_mem_out_alu_res_p_17_port, s_mem_out_alu_res_p_16_port, 
      s_mem_out_alu_res_p_15_port, s_mem_out_alu_res_p_14_port, 
      s_mem_out_alu_res_p_13_port, s_mem_out_alu_res_p_12_port, 
      s_wb_in_memtoReg_p, s_writeback_data_31_port, s_writeback_data_30_port, 
      s_writeback_data_29_port, s_writeback_data_28_port, 
      s_writeback_data_27_port, s_writeback_data_26_port, 
      s_writeback_data_25_port, s_writeback_data_24_port, 
      s_writeback_data_23_port, s_writeback_data_22_port, 
      s_writeback_data_21_port, s_writeback_data_20_port, 
      s_writeback_data_19_port, s_writeback_data_18_port, 
      s_writeback_data_17_port, s_writeback_data_16_port, 
      s_writeback_data_15_port, s_writeback_data_14_port, 
      s_writeback_data_13_port, s_writeback_data_12_port, 
      s_writeback_data_11_port, s_writeback_data_10_port, 
      s_writeback_data_9_port, s_writeback_data_8_port, s_writeback_data_7_port
      , s_writeback_data_6_port, s_writeback_data_5_port, 
      s_writeback_data_4_port, s_writeback_data_3_port, s_writeback_data_2_port
      , s_writeback_data_1_port, s_writeback_data_0_port, 
      s_wb_in_alu_res_p_31_port, s_wb_in_alu_res_p_30_port, 
      s_wb_in_alu_res_p_29_port, s_wb_in_alu_res_p_28_port, 
      s_wb_in_alu_res_p_27_port, s_wb_in_alu_res_p_26_port, 
      s_wb_in_alu_res_p_25_port, s_wb_in_alu_res_p_24_port, 
      s_wb_in_alu_res_p_23_port, s_wb_in_alu_res_p_22_port, 
      s_wb_in_alu_res_p_21_port, s_wb_in_alu_res_p_20_port, 
      s_wb_in_alu_res_p_19_port, s_wb_in_alu_res_p_18_port, 
      s_wb_in_alu_res_p_17_port, s_wb_in_alu_res_p_16_port, 
      s_wb_in_alu_res_p_15_port, s_wb_in_alu_res_p_14_port, 
      s_wb_in_alu_res_p_13_port, s_wb_in_alu_res_p_12_port, 
      s_wb_in_alu_res_p_11_port, s_wb_in_alu_res_p_10_port, 
      s_wb_in_alu_res_p_9_port, s_wb_in_alu_res_p_8_port, 
      s_wb_in_alu_res_p_7_port, s_wb_in_alu_res_p_6_port, 
      s_wb_in_alu_res_p_5_port, s_wb_in_alu_res_p_4_port, 
      s_wb_in_alu_res_p_3_port, s_wb_in_alu_res_p_2_port, 
      s_wb_in_alu_res_p_1_port, s_wb_in_alu_res_p_0_port, s_forward_A_1_port, 
      s_forward_A_0_port, s_src_a_31_port, s_src_a_30_port, s_src_a_29_port, 
      s_src_a_28_port, s_src_a_27_port, s_src_a_26_port, s_src_a_25_port, 
      s_src_a_24_port, s_src_a_23_port, s_src_a_22_port, s_src_a_21_port, 
      s_src_a_20_port, s_src_a_19_port, s_src_a_18_port, s_src_a_17_port, 
      s_src_a_16_port, s_src_a_15_port, s_src_a_14_port, s_src_a_13_port, 
      s_src_a_12_port, s_src_a_11_port, s_src_a_10_port, s_src_a_9_port, 
      s_src_a_8_port, s_src_a_7_port, s_src_a_6_port, s_src_a_5_port, 
      s_src_a_4_port, s_src_a_3_port, s_src_a_2_port, s_src_a_1_port, 
      s_src_a_0_port, s_exe_in_regA_p_31_port, s_exe_in_regA_p_30_port, 
      s_exe_in_regA_p_29_port, s_exe_in_regA_p_28_port, s_exe_in_regA_p_27_port
      , s_exe_in_regA_p_26_port, s_exe_in_regA_p_25_port, 
      s_exe_in_regA_p_24_port, s_exe_in_regA_p_23_port, s_exe_in_regA_p_22_port
      , s_exe_in_regA_p_21_port, s_exe_in_regA_p_20_port, 
      s_exe_in_regA_p_19_port, s_exe_in_regA_p_18_port, s_exe_in_regA_p_17_port
      , s_exe_in_regA_p_16_port, s_exe_in_regA_p_15_port, 
      s_exe_in_regA_p_14_port, s_exe_in_regA_p_13_port, s_exe_in_regA_p_12_port
      , s_exe_in_regA_p_11_port, s_exe_in_regA_p_10_port, 
      s_exe_in_regA_p_9_port, s_exe_in_regA_p_8_port, s_exe_in_regA_p_7_port, 
      s_exe_in_regA_p_6_port, s_exe_in_regA_p_5_port, s_exe_in_regA_p_4_port, 
      s_exe_in_regA_p_3_port, s_exe_in_regA_p_2_port, s_exe_in_regA_p_1_port, 
      s_exe_in_regA_p_0_port, s_forward_B_1_port, s_forward_B_0_port, 
      s_src_b_31_port, s_src_b_30_port, s_src_b_29_port, s_src_b_28_port, 
      s_src_b_27_port, s_src_b_26_port, s_src_b_25_port, s_src_b_24_port, 
      s_src_b_23_port, s_src_b_22_port, s_src_b_21_port, s_src_b_20_port, 
      s_src_b_19_port, s_src_b_18_port, s_src_b_17_port, s_src_b_16_port, 
      s_src_b_15_port, s_src_b_14_port, s_src_b_13_port, s_src_b_12_port, 
      s_src_b_11_port, s_src_b_10_port, s_src_b_9_port, s_src_b_8_port, 
      s_src_b_7_port, s_src_b_6_port, s_src_b_5_port, s_src_b_4_port, 
      s_src_b_3_port, s_src_b_2_port, s_src_b_1_port, s_src_b_0_port, 
      s_exe_in_regB_p_31_port, s_exe_in_regB_p_30_port, s_exe_in_regB_p_29_port
      , s_exe_in_regB_p_28_port, s_exe_in_regB_p_27_port, 
      s_exe_in_regB_p_26_port, s_exe_in_regB_p_25_port, s_exe_in_regB_p_24_port
      , s_exe_in_regB_p_23_port, s_exe_in_regB_p_22_port, 
      s_exe_in_regB_p_21_port, s_exe_in_regB_p_20_port, s_exe_in_regB_p_19_port
      , s_exe_in_regB_p_18_port, s_exe_in_regB_p_17_port, 
      s_exe_in_regB_p_16_port, s_exe_in_regB_p_15_port, s_exe_in_regB_p_14_port
      , s_exe_in_regB_p_13_port, s_exe_in_regB_p_12_port, 
      s_exe_in_regB_p_11_port, s_exe_in_regB_p_10_port, s_exe_in_regB_p_9_port,
      s_exe_in_regB_p_8_port, s_exe_in_regB_p_7_port, s_exe_in_regB_p_6_port, 
      s_exe_in_regB_p_5_port, s_exe_in_regB_p_4_port, s_exe_in_regB_p_3_port, 
      s_exe_in_regB_p_2_port, s_exe_in_regB_p_1_port, s_exe_in_regB_p_0_port, 
      s_id_ctrl_opcode_5_port, s_id_ctrl_opcode_4_port, s_id_ctrl_opcode_3_port
      , s_id_ctrl_opcode_2_port, s_id_ctrl_opcode_1_port, 
      s_id_ctrl_opcode_0_port, s_ctrl_out_RegDst_p, s_ctrl_out_ALUsrc_B_p, 
      s_ctrl_out_memtoReg_p, s_ctrl_out_regWrite_p, s_ctrl_out_memWen_n_p, 
      s_ctrl_out_cALU_OP_p_3_port, s_ctrl_out_cALU_OP_p_2_port, 
      s_ctrl_out_cALU_OP_p_1_port, s_ctrl_out_cALU_OP_p_0_port, 
      s_exe_if_branch_pc_11_port, s_exe_if_branch_pc_10_port, 
      s_exe_if_branch_pc_9_port, s_exe_if_branch_pc_8_port, 
      s_exe_if_branch_pc_7_port, s_exe_if_branch_pc_6_port, 
      s_exe_if_branch_pc_5_port, s_exe_if_branch_pc_4_port, 
      s_exe_if_branch_pc_3_port, s_exe_if_branch_pc_2_port, 
      s_exe_if_branch_pc_1_port, s_exe_if_branch_pc_0_port, 
      s_if_out_pc_plus1_p_11_port, s_if_out_pc_plus1_p_10_port, 
      s_if_out_pc_plus1_p_9_port, s_if_out_pc_plus1_p_8_port, 
      s_if_out_pc_plus1_p_7_port, s_if_out_pc_plus1_p_6_port, 
      s_if_out_pc_plus1_p_5_port, s_if_out_pc_plus1_p_4_port, 
      s_if_out_pc_plus1_p_3_port, s_if_out_pc_plus1_p_2_port, 
      s_if_out_pc_plus1_p_1_port, s_if_out_pc_plus1_p_0_port, 
      s_regfile_forward_A, s_regfile_forward_B, s_wb_in_regWrite_p, 
      s_wb_in_write_reg_p_4_port, s_wb_in_write_reg_p_3_port, 
      s_wb_in_write_reg_p_2_port, s_wb_in_write_reg_p_1_port, 
      s_wb_in_write_reg_p_0_port, s_id_out_regA_p_31_port, 
      s_id_out_regA_p_30_port, s_id_out_regA_p_29_port, s_id_out_regA_p_28_port
      , s_id_out_regA_p_27_port, s_id_out_regA_p_26_port, 
      s_id_out_regA_p_25_port, s_id_out_regA_p_24_port, s_id_out_regA_p_23_port
      , s_id_out_regA_p_22_port, s_id_out_regA_p_21_port, 
      s_id_out_regA_p_20_port, s_id_out_regA_p_19_port, s_id_out_regA_p_18_port
      , s_id_out_regA_p_17_port, s_id_out_regA_p_16_port, 
      s_id_out_regA_p_15_port, s_id_out_regA_p_14_port, s_id_out_regA_p_13_port
      , s_id_out_regA_p_12_port, s_id_out_regA_p_11_port, 
      s_id_out_regA_p_10_port, s_id_out_regA_p_9_port, s_id_out_regA_p_8_port, 
      s_id_out_regA_p_7_port, s_id_out_regA_p_6_port, s_id_out_regA_p_5_port, 
      s_id_out_regA_p_4_port, s_id_out_regA_p_3_port, s_id_out_regA_p_2_port, 
      s_id_out_regA_p_1_port, s_id_out_regA_p_0_port, s_id_out_regB_p_31_port, 
      s_id_out_regB_p_30_port, s_id_out_regB_p_29_port, s_id_out_regB_p_28_port
      , s_id_out_regB_p_27_port, s_id_out_regB_p_26_port, 
      s_id_out_regB_p_25_port, s_id_out_regB_p_24_port, s_id_out_regB_p_23_port
      , s_id_out_regB_p_22_port, s_id_out_regB_p_21_port, 
      s_id_out_regB_p_20_port, s_id_out_regB_p_19_port, s_id_out_regB_p_18_port
      , s_id_out_regB_p_17_port, s_id_out_regB_p_16_port, 
      s_id_out_regB_p_15_port, s_id_out_regB_p_14_port, s_id_out_regB_p_13_port
      , s_id_out_regB_p_12_port, s_id_out_regB_p_11_port, 
      s_id_out_regB_p_10_port, s_id_out_regB_p_9_port, s_id_out_regB_p_8_port, 
      s_id_out_regB_p_7_port, s_id_out_regB_p_6_port, s_id_out_regB_p_5_port, 
      s_id_out_regB_p_4_port, s_id_out_regB_p_3_port, s_id_out_regB_p_2_port, 
      s_id_out_regB_p_1_port, s_id_out_regB_p_0_port, s_id_out_RS_p_4_port, 
      s_id_out_RS_p_3_port, s_id_out_RS_p_2_port, s_id_out_RS_p_1_port, 
      s_id_out_RS_p_0_port, s_id_out_RT_p_4_port, s_id_out_RT_p_3_port, 
      s_id_out_RT_p_2_port, s_id_out_RT_p_1_port, s_id_out_RT_p_0_port, 
      s_id_out_RD_p_4_port, s_id_out_RD_p_3_port, s_id_out_RD_p_2_port, 
      s_id_out_RD_p_1_port, s_id_out_RD_p_0_port, s_id_out_shamt_p_4_port, 
      s_id_out_shamt_p_3_port, s_id_out_shamt_p_2_port, s_id_out_shamt_p_1_port
      , s_id_out_shamt_p_0_port, s_id_out_funct_p_5_port, 
      s_id_out_funct_p_4_port, s_id_out_funct_p_3_port, s_id_out_funct_p_2_port
      , s_id_out_funct_p_1_port, s_id_out_funct_p_0_port, 
      s_id_out_sign_extend_p_31_port, s_id_out_sign_extend_p_30_port, 
      s_id_out_sign_extend_p_29_port, s_id_out_sign_extend_p_28_port, 
      s_id_out_sign_extend_p_27_port, s_id_out_sign_extend_p_26_port, 
      s_id_out_sign_extend_p_25_port, s_id_out_sign_extend_p_24_port, 
      s_id_out_sign_extend_p_23_port, s_id_out_sign_extend_p_22_port, 
      s_id_out_sign_extend_p_21_port, s_id_out_sign_extend_p_20_port, 
      s_id_out_sign_extend_p_19_port, s_id_out_sign_extend_p_18_port, 
      s_id_out_sign_extend_p_17_port, s_id_out_sign_extend_p_16_port, 
      s_id_out_sign_extend_p_15_port, s_id_out_sign_extend_p_14_port, 
      s_id_out_sign_extend_p_13_port, s_id_out_sign_extend_p_12_port, 
      s_id_out_sign_extend_p_11_port, s_id_out_sign_extend_p_10_port, 
      s_id_out_sign_extend_p_9_port, s_id_out_sign_extend_p_8_port, 
      s_id_out_sign_extend_p_7_port, s_id_out_sign_extend_p_6_port, 
      s_id_out_sign_extend_p_5_port, s_id_out_sign_extend_p_4_port, 
      s_id_out_sign_extend_p_3_port, s_id_out_sign_extend_p_2_port, 
      s_id_out_sign_extend_p_1_port, s_id_out_sign_extend_p_0_port, 
      s_exe_in_shamt_p_4_port, s_exe_in_shamt_p_3_port, s_exe_in_shamt_p_2_port
      , s_exe_in_shamt_p_1_port, s_exe_in_shamt_p_0_port, 
      s_exe_in_funct_p_5_port, s_exe_in_funct_p_4_port, s_exe_in_funct_p_3_port
      , s_exe_in_funct_p_2_port, s_exe_in_funct_p_1_port, 
      s_exe_in_funct_p_0_port, s_exe_in_sign_extend_p_31_port, 
      s_exe_in_sign_extend_p_30_port, s_exe_in_sign_extend_p_29_port, 
      s_exe_in_sign_extend_p_28_port, s_exe_in_sign_extend_p_27_port, 
      s_exe_in_sign_extend_p_26_port, s_exe_in_sign_extend_p_25_port, 
      s_exe_in_sign_extend_p_24_port, s_exe_in_sign_extend_p_23_port, 
      s_exe_in_sign_extend_p_22_port, s_exe_in_sign_extend_p_21_port, 
      s_exe_in_sign_extend_p_20_port, s_exe_in_sign_extend_p_19_port, 
      s_exe_in_sign_extend_p_18_port, s_exe_in_sign_extend_p_17_port, 
      s_exe_in_sign_extend_p_16_port, s_exe_in_sign_extend_p_15_port, 
      s_exe_in_sign_extend_p_14_port, s_exe_in_sign_extend_p_13_port, 
      s_exe_in_sign_extend_p_12_port, s_exe_in_sign_extend_p_11_port, 
      s_exe_in_sign_extend_p_10_port, s_exe_in_sign_extend_p_9_port, 
      s_exe_in_sign_extend_p_8_port, s_exe_in_sign_extend_p_7_port, 
      s_exe_in_sign_extend_p_6_port, s_exe_in_sign_extend_p_5_port, 
      s_exe_in_sign_extend_p_4_port, s_exe_in_sign_extend_p_3_port, 
      s_exe_in_sign_extend_p_2_port, s_exe_in_sign_extend_p_1_port, 
      s_exe_in_sign_extend_p_0_port, s_exe_in_pc_plus1_p_11_port, 
      s_exe_in_pc_plus1_p_10_port, s_exe_in_pc_plus1_p_9_port, 
      s_exe_in_pc_plus1_p_8_port, s_exe_in_pc_plus1_p_7_port, 
      s_exe_in_pc_plus1_p_6_port, s_exe_in_pc_plus1_p_5_port, 
      s_exe_in_pc_plus1_p_4_port, s_exe_in_pc_plus1_p_3_port, 
      s_exe_in_pc_plus1_p_2_port, s_exe_in_pc_plus1_p_1_port, 
      s_exe_in_pc_plus1_p_0_port, s_exe_in_RS_p_4_port, s_exe_in_RS_p_3_port, 
      s_exe_in_RS_p_2_port, s_exe_in_RS_p_1_port, s_exe_in_RS_p_0_port, 
      s_exe_in_RT_p_4_port, s_exe_in_RT_p_3_port, s_exe_in_RT_p_2_port, 
      s_exe_in_RT_p_1_port, s_exe_in_RT_p_0_port, s_exe_in_RD_p_4_port, 
      s_exe_in_RD_p_3_port, s_exe_in_RD_p_2_port, s_exe_in_RD_p_1_port, 
      s_exe_in_RD_p_0_port, s_exe_in_ALUsrc_B_p, s_exe_in_cALU_OP_p_3_port, 
      s_exe_in_cALU_OP_p_2_port, s_exe_in_cALU_OP_p_1_port, 
      s_exe_in_cALU_OP_p_0_port, s_exe_in_RegDst_p, s_exe_out_alu_res_p_31_port
      , s_exe_out_alu_res_p_30_port, s_exe_out_alu_res_p_29_port, 
      s_exe_out_alu_res_p_28_port, s_exe_out_alu_res_p_27_port, 
      s_exe_out_alu_res_p_26_port, s_exe_out_alu_res_p_25_port, 
      s_exe_out_alu_res_p_24_port, s_exe_out_alu_res_p_23_port, 
      s_exe_out_alu_res_p_22_port, s_exe_out_alu_res_p_21_port, 
      s_exe_out_alu_res_p_20_port, s_exe_out_alu_res_p_19_port, 
      s_exe_out_alu_res_p_18_port, s_exe_out_alu_res_p_17_port, 
      s_exe_out_alu_res_p_16_port, s_exe_out_alu_res_p_15_port, 
      s_exe_out_alu_res_p_14_port, s_exe_out_alu_res_p_13_port, 
      s_exe_out_alu_res_p_12_port, s_exe_out_alu_res_p_11_port, 
      s_exe_out_alu_res_p_10_port, s_exe_out_alu_res_p_9_port, 
      s_exe_out_alu_res_p_8_port, s_exe_out_alu_res_p_7_port, 
      s_exe_out_alu_res_p_6_port, s_exe_out_alu_res_p_5_port, 
      s_exe_out_alu_res_p_4_port, s_exe_out_alu_res_p_3_port, 
      s_exe_out_alu_res_p_2_port, s_exe_out_alu_res_p_1_port, 
      s_exe_out_alu_res_p_0_port, s_exe_out_write_reg_p_4_port, 
      s_exe_out_write_reg_p_3_port, s_exe_out_write_reg_p_2_port, 
      s_exe_out_write_reg_p_1_port, s_exe_out_write_reg_p_0_port, 
      s_exe_out_dmem_data_p_31_port, s_exe_out_dmem_data_p_30_port, 
      s_exe_out_dmem_data_p_29_port, s_exe_out_dmem_data_p_28_port, 
      s_exe_out_dmem_data_p_27_port, s_exe_out_dmem_data_p_26_port, 
      s_exe_out_dmem_data_p_25_port, s_exe_out_dmem_data_p_24_port, 
      s_exe_out_dmem_data_p_23_port, s_exe_out_dmem_data_p_22_port, 
      s_exe_out_dmem_data_p_21_port, s_exe_out_dmem_data_p_20_port, 
      s_exe_out_dmem_data_p_19_port, s_exe_out_dmem_data_p_18_port, 
      s_exe_out_dmem_data_p_17_port, s_exe_out_dmem_data_p_16_port, 
      s_exe_out_dmem_data_p_15_port, s_exe_out_dmem_data_p_14_port, 
      s_exe_out_dmem_data_p_13_port, s_exe_out_dmem_data_p_12_port, 
      s_exe_out_dmem_data_p_11_port, s_exe_out_dmem_data_p_10_port, 
      s_exe_out_dmem_data_p_9_port, s_exe_out_dmem_data_p_8_port, 
      s_exe_out_dmem_data_p_7_port, s_exe_out_dmem_data_p_6_port, 
      s_exe_out_dmem_data_p_5_port, s_exe_out_dmem_data_p_4_port, 
      s_exe_out_dmem_data_p_3_port, s_exe_out_dmem_data_p_2_port, 
      s_exe_out_dmem_data_p_1_port, s_exe_out_dmem_data_p_0_port, n4, n6, n7, 
      n9, n1, n2, n3, n5, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n_1021, n_1022 : std_logic;

begin
   mini_mips_o <= ( mini_mips_o_DMEM_ADDR_11_port, 
      mini_mips_o_DMEM_ADDR_10_port, mini_mips_o_DMEM_ADDR_9_port, 
      mini_mips_o_DMEM_ADDR_8_port, mini_mips_o_DMEM_ADDR_7_port, 
      mini_mips_o_DMEM_ADDR_6_port, mini_mips_o_DMEM_ADDR_5_port, 
      mini_mips_o_DMEM_ADDR_4_port, mini_mips_o_DMEM_ADDR_3_port, 
      mini_mips_o_DMEM_ADDR_2_port, mini_mips_o_DMEM_ADDR_1_port, 
      mini_mips_o_DMEM_ADDR_0_port, mini_mips_o_DMEM_DATA_31_port, 
      mini_mips_o_DMEM_DATA_30_port, mini_mips_o_DMEM_DATA_29_port, 
      mini_mips_o_DMEM_DATA_28_port, mini_mips_o_DMEM_DATA_27_port, 
      mini_mips_o_DMEM_DATA_26_port, mini_mips_o_DMEM_DATA_25_port, 
      mini_mips_o_DMEM_DATA_24_port, mini_mips_o_DMEM_DATA_23_port, 
      mini_mips_o_DMEM_DATA_22_port, mini_mips_o_DMEM_DATA_21_port, 
      mini_mips_o_DMEM_DATA_20_port, mini_mips_o_DMEM_DATA_19_port, 
      mini_mips_o_DMEM_DATA_18_port, mini_mips_o_DMEM_DATA_17_port, 
      mini_mips_o_DMEM_DATA_16_port, mini_mips_o_DMEM_DATA_15_port, 
      mini_mips_o_DMEM_DATA_14_port, mini_mips_o_DMEM_DATA_13_port, 
      mini_mips_o_DMEM_DATA_12_port, mini_mips_o_DMEM_DATA_11_port, 
      mini_mips_o_DMEM_DATA_10_port, mini_mips_o_DMEM_DATA_9_port, 
      mini_mips_o_DMEM_DATA_8_port, mini_mips_o_DMEM_DATA_7_port, 
      mini_mips_o_DMEM_DATA_6_port, mini_mips_o_DMEM_DATA_5_port, 
      mini_mips_o_DMEM_DATA_4_port, mini_mips_o_DMEM_DATA_3_port, 
      mini_mips_o_DMEM_DATA_2_port, mini_mips_o_DMEM_DATA_1_port, 
      mini_mips_o_DMEM_DATA_0_port, mini_mips_o_IMEM_ADDR_11_port, 
      mini_mips_o_IMEM_ADDR_10_port, mini_mips_o_IMEM_ADDR_9_port, 
      mini_mips_o_IMEM_ADDR_8_port, mini_mips_o_IMEM_ADDR_7_port, 
      mini_mips_o_IMEM_ADDR_6_port, mini_mips_o_IMEM_ADDR_5_port, 
      mini_mips_o_IMEM_ADDR_4_port, mini_mips_o_IMEM_ADDR_3_port, 
      mini_mips_o_IMEM_ADDR_2_port, mini_mips_o_IMEM_ADDR_1_port, 
      mini_mips_o_IMEM_ADDR_0_port, mini_mips_o_DMEM_WEN_N_port );
   
   X_Logic0_port <= '0';
   ctrl_inst : controller port map( ctrl_i(5) => s_id_ctrl_opcode_5_port, 
                           ctrl_i(4) => s_id_ctrl_opcode_4_port, ctrl_i(3) => 
                           s_id_ctrl_opcode_3_port, ctrl_i(2) => 
                           s_id_ctrl_opcode_2_port, ctrl_i(1) => 
                           s_id_ctrl_opcode_1_port, ctrl_i(0) => 
                           s_id_ctrl_opcode_0_port, ctrl_o(9) => 
                           s_ctrl_out_RegDst_p, ctrl_o(8) => 
                           s_ctrl_out_ALUsrc_B_p, ctrl_o(7) => 
                           s_ctrl_out_memtoReg_p, ctrl_o(6) => 
                           s_ctrl_out_regWrite_p, ctrl_o(5) => 
                           s_ctrl_out_memWen_n_p, ctrl_o(4) => n_1021, 
                           ctrl_o(3) => n_1022, ctrl_o(2) => 
                           s_ctrl_out_cALU_OP_p_2_port, ctrl_o(1) => 
                           s_ctrl_out_cALU_OP_p_1_port, ctrl_o(0) => 
                           s_ctrl_out_cALU_OP_p_0_port);
   if_top_inst : if_top port map( clk => clk, rst_n => n35, if_top_i(13) => 
                           X_Logic0_port, if_top_i(12) => 
                           s_exe_if_branch_pc_11_port, if_top_i(11) => 
                           s_exe_if_branch_pc_10_port, if_top_i(10) => 
                           s_exe_if_branch_pc_9_port, if_top_i(9) => 
                           s_exe_if_branch_pc_8_port, if_top_i(8) => 
                           s_exe_if_branch_pc_7_port, if_top_i(7) => 
                           s_exe_if_branch_pc_6_port, if_top_i(6) => 
                           s_exe_if_branch_pc_5_port, if_top_i(5) => 
                           s_exe_if_branch_pc_4_port, if_top_i(4) => 
                           s_exe_if_branch_pc_3_port, if_top_i(3) => 
                           s_exe_if_branch_pc_2_port, if_top_i(2) => 
                           s_exe_if_branch_pc_1_port, if_top_i(1) => 
                           s_exe_if_branch_pc_0_port, if_top_i(0) => s_if_PCSrc
                           , if_top_o(23) => mini_mips_o_IMEM_ADDR_11_port, 
                           if_top_o(22) => mini_mips_o_IMEM_ADDR_10_port, 
                           if_top_o(21) => mini_mips_o_IMEM_ADDR_9_port, 
                           if_top_o(20) => mini_mips_o_IMEM_ADDR_8_port, 
                           if_top_o(19) => mini_mips_o_IMEM_ADDR_7_port, 
                           if_top_o(18) => mini_mips_o_IMEM_ADDR_6_port, 
                           if_top_o(17) => mini_mips_o_IMEM_ADDR_5_port, 
                           if_top_o(16) => mini_mips_o_IMEM_ADDR_4_port, 
                           if_top_o(15) => mini_mips_o_IMEM_ADDR_3_port, 
                           if_top_o(14) => mini_mips_o_IMEM_ADDR_2_port, 
                           if_top_o(13) => mini_mips_o_IMEM_ADDR_1_port, 
                           if_top_o(12) => mini_mips_o_IMEM_ADDR_0_port, 
                           if_top_o(11) => s_if_out_pc_plus1_p_11_port, 
                           if_top_o(10) => s_if_out_pc_plus1_p_10_port, 
                           if_top_o(9) => s_if_out_pc_plus1_p_9_port, 
                           if_top_o(8) => s_if_out_pc_plus1_p_8_port, 
                           if_top_o(7) => s_if_out_pc_plus1_p_7_port, 
                           if_top_o(6) => s_if_out_pc_plus1_p_6_port, 
                           if_top_o(5) => s_if_out_pc_plus1_p_5_port, 
                           if_top_o(4) => s_if_out_pc_plus1_p_4_port, 
                           if_top_o(3) => s_if_out_pc_plus1_p_3_port, 
                           if_top_o(2) => s_if_out_pc_plus1_p_2_port, 
                           if_top_o(1) => s_if_out_pc_plus1_p_1_port, 
                           if_top_o(0) => s_if_out_pc_plus1_p_0_port);
   if_id_inst : if_id port map( clk => clk, rst_n => n34, halt_i => 
                           X_Logic0_port, IF_ID_i(11) => 
                           s_if_out_pc_plus1_p_11_port, IF_ID_i(10) => 
                           s_if_out_pc_plus1_p_10_port, IF_ID_i(9) => 
                           s_if_out_pc_plus1_p_9_port, IF_ID_i(8) => 
                           s_if_out_pc_plus1_p_8_port, IF_ID_i(7) => 
                           s_if_out_pc_plus1_p_7_port, IF_ID_i(6) => 
                           s_if_out_pc_plus1_p_6_port, IF_ID_i(5) => 
                           s_if_out_pc_plus1_p_5_port, IF_ID_i(4) => 
                           s_if_out_pc_plus1_p_4_port, IF_ID_i(3) => 
                           s_if_out_pc_plus1_p_3_port, IF_ID_i(2) => 
                           s_if_out_pc_plus1_p_2_port, IF_ID_i(1) => 
                           s_if_out_pc_plus1_p_1_port, IF_ID_i(0) => 
                           s_if_out_pc_plus1_p_0_port, IF_ID_o(11) => 
                           s_id_out_pc_plus1_p_11_port, IF_ID_o(10) => 
                           s_id_out_pc_plus1_p_10_port, IF_ID_o(9) => 
                           s_id_out_pc_plus1_p_9_port, IF_ID_o(8) => 
                           s_id_out_pc_plus1_p_8_port, IF_ID_o(7) => 
                           s_id_out_pc_plus1_p_7_port, IF_ID_o(6) => 
                           s_id_out_pc_plus1_p_6_port, IF_ID_o(5) => 
                           s_id_out_pc_plus1_p_5_port, IF_ID_o(4) => 
                           s_id_out_pc_plus1_p_4_port, IF_ID_o(3) => 
                           s_id_out_pc_plus1_p_3_port, IF_ID_o(2) => 
                           s_id_out_pc_plus1_p_2_port, IF_ID_o(1) => 
                           s_id_out_pc_plus1_p_1_port, IF_ID_o(0) => 
                           s_id_out_pc_plus1_p_0_port);
   id_top_inst : id_top port map( clk => clk, rst_n => n33, id_top_i(71) => 
                           mini_mips_i(31), id_top_i(70) => mini_mips_i(30), 
                           id_top_i(69) => mini_mips_i(29), id_top_i(68) => 
                           mini_mips_i(28), id_top_i(67) => mini_mips_i(27), 
                           id_top_i(66) => mini_mips_i(26), id_top_i(65) => 
                           mini_mips_i(25), id_top_i(64) => mini_mips_i(24), 
                           id_top_i(63) => mini_mips_i(23), id_top_i(62) => 
                           mini_mips_i(22), id_top_i(61) => mini_mips_i(21), 
                           id_top_i(60) => mini_mips_i(20), id_top_i(59) => 
                           mini_mips_i(19), id_top_i(58) => mini_mips_i(18), 
                           id_top_i(57) => mini_mips_i(17), id_top_i(56) => 
                           mini_mips_i(16), id_top_i(55) => mini_mips_i(15), 
                           id_top_i(54) => mini_mips_i(14), id_top_i(53) => 
                           mini_mips_i(13), id_top_i(52) => mini_mips_i(12), 
                           id_top_i(51) => mini_mips_i(11), id_top_i(50) => 
                           mini_mips_i(10), id_top_i(49) => mini_mips_i(9), 
                           id_top_i(48) => mini_mips_i(8), id_top_i(47) => 
                           mini_mips_i(7), id_top_i(46) => mini_mips_i(6), 
                           id_top_i(45) => mini_mips_i(5), id_top_i(44) => 
                           mini_mips_i(4), id_top_i(43) => mini_mips_i(3), 
                           id_top_i(42) => mini_mips_i(2), id_top_i(41) => 
                           mini_mips_i(1), id_top_i(40) => mini_mips_i(0), 
                           id_top_i(39) => s_writeback_data_31_port, 
                           id_top_i(38) => s_writeback_data_30_port, 
                           id_top_i(37) => s_writeback_data_29_port, 
                           id_top_i(36) => s_writeback_data_28_port, 
                           id_top_i(35) => s_writeback_data_27_port, 
                           id_top_i(34) => s_writeback_data_26_port, 
                           id_top_i(33) => s_writeback_data_25_port, 
                           id_top_i(32) => s_writeback_data_24_port, 
                           id_top_i(31) => s_writeback_data_23_port, 
                           id_top_i(30) => s_writeback_data_22_port, 
                           id_top_i(29) => s_writeback_data_21_port, 
                           id_top_i(28) => s_writeback_data_20_port, 
                           id_top_i(27) => s_writeback_data_19_port, 
                           id_top_i(26) => s_writeback_data_18_port, 
                           id_top_i(25) => s_writeback_data_17_port, 
                           id_top_i(24) => s_writeback_data_16_port, 
                           id_top_i(23) => s_writeback_data_15_port, 
                           id_top_i(22) => s_writeback_data_14_port, 
                           id_top_i(21) => s_writeback_data_13_port, 
                           id_top_i(20) => s_writeback_data_12_port, 
                           id_top_i(19) => s_writeback_data_11_port, 
                           id_top_i(18) => s_writeback_data_10_port, 
                           id_top_i(17) => s_writeback_data_9_port, 
                           id_top_i(16) => s_writeback_data_8_port, 
                           id_top_i(15) => s_writeback_data_7_port, 
                           id_top_i(14) => s_writeback_data_6_port, 
                           id_top_i(13) => s_writeback_data_5_port, 
                           id_top_i(12) => s_writeback_data_4_port, 
                           id_top_i(11) => s_writeback_data_3_port, 
                           id_top_i(10) => s_writeback_data_2_port, id_top_i(9)
                           => s_writeback_data_1_port, id_top_i(8) => 
                           s_writeback_data_0_port, id_top_i(7) => 
                           s_regfile_forward_A, id_top_i(6) => 
                           s_regfile_forward_B, id_top_i(5) => 
                           s_wb_in_regWrite_p, id_top_i(4) => 
                           s_wb_in_write_reg_p_4_port, id_top_i(3) => 
                           s_wb_in_write_reg_p_3_port, id_top_i(2) => 
                           s_wb_in_write_reg_p_2_port, id_top_i(1) => 
                           s_wb_in_write_reg_p_1_port, id_top_i(0) => 
                           s_wb_in_write_reg_p_0_port, id_top_o(127) => 
                           s_id_out_regA_p_31_port, id_top_o(126) => 
                           s_id_out_regA_p_30_port, id_top_o(125) => 
                           s_id_out_regA_p_29_port, id_top_o(124) => 
                           s_id_out_regA_p_28_port, id_top_o(123) => 
                           s_id_out_regA_p_27_port, id_top_o(122) => 
                           s_id_out_regA_p_26_port, id_top_o(121) => 
                           s_id_out_regA_p_25_port, id_top_o(120) => 
                           s_id_out_regA_p_24_port, id_top_o(119) => 
                           s_id_out_regA_p_23_port, id_top_o(118) => 
                           s_id_out_regA_p_22_port, id_top_o(117) => 
                           s_id_out_regA_p_21_port, id_top_o(116) => 
                           s_id_out_regA_p_20_port, id_top_o(115) => 
                           s_id_out_regA_p_19_port, id_top_o(114) => 
                           s_id_out_regA_p_18_port, id_top_o(113) => 
                           s_id_out_regA_p_17_port, id_top_o(112) => 
                           s_id_out_regA_p_16_port, id_top_o(111) => 
                           s_id_out_regA_p_15_port, id_top_o(110) => 
                           s_id_out_regA_p_14_port, id_top_o(109) => 
                           s_id_out_regA_p_13_port, id_top_o(108) => 
                           s_id_out_regA_p_12_port, id_top_o(107) => 
                           s_id_out_regA_p_11_port, id_top_o(106) => 
                           s_id_out_regA_p_10_port, id_top_o(105) => 
                           s_id_out_regA_p_9_port, id_top_o(104) => 
                           s_id_out_regA_p_8_port, id_top_o(103) => 
                           s_id_out_regA_p_7_port, id_top_o(102) => 
                           s_id_out_regA_p_6_port, id_top_o(101) => 
                           s_id_out_regA_p_5_port, id_top_o(100) => 
                           s_id_out_regA_p_4_port, id_top_o(99) => 
                           s_id_out_regA_p_3_port, id_top_o(98) => 
                           s_id_out_regA_p_2_port, id_top_o(97) => 
                           s_id_out_regA_p_1_port, id_top_o(96) => 
                           s_id_out_regA_p_0_port, id_top_o(95) => 
                           s_id_out_regB_p_31_port, id_top_o(94) => 
                           s_id_out_regB_p_30_port, id_top_o(93) => 
                           s_id_out_regB_p_29_port, id_top_o(92) => 
                           s_id_out_regB_p_28_port, id_top_o(91) => 
                           s_id_out_regB_p_27_port, id_top_o(90) => 
                           s_id_out_regB_p_26_port, id_top_o(89) => 
                           s_id_out_regB_p_25_port, id_top_o(88) => 
                           s_id_out_regB_p_24_port, id_top_o(87) => 
                           s_id_out_regB_p_23_port, id_top_o(86) => 
                           s_id_out_regB_p_22_port, id_top_o(85) => 
                           s_id_out_regB_p_21_port, id_top_o(84) => 
                           s_id_out_regB_p_20_port, id_top_o(83) => 
                           s_id_out_regB_p_19_port, id_top_o(82) => 
                           s_id_out_regB_p_18_port, id_top_o(81) => 
                           s_id_out_regB_p_17_port, id_top_o(80) => 
                           s_id_out_regB_p_16_port, id_top_o(79) => 
                           s_id_out_regB_p_15_port, id_top_o(78) => 
                           s_id_out_regB_p_14_port, id_top_o(77) => 
                           s_id_out_regB_p_13_port, id_top_o(76) => 
                           s_id_out_regB_p_12_port, id_top_o(75) => 
                           s_id_out_regB_p_11_port, id_top_o(74) => 
                           s_id_out_regB_p_10_port, id_top_o(73) => 
                           s_id_out_regB_p_9_port, id_top_o(72) => 
                           s_id_out_regB_p_8_port, id_top_o(71) => 
                           s_id_out_regB_p_7_port, id_top_o(70) => 
                           s_id_out_regB_p_6_port, id_top_o(69) => 
                           s_id_out_regB_p_5_port, id_top_o(68) => 
                           s_id_out_regB_p_4_port, id_top_o(67) => 
                           s_id_out_regB_p_3_port, id_top_o(66) => 
                           s_id_out_regB_p_2_port, id_top_o(65) => 
                           s_id_out_regB_p_1_port, id_top_o(64) => 
                           s_id_out_regB_p_0_port, id_top_o(63) => 
                           s_id_ctrl_opcode_5_port, id_top_o(62) => 
                           s_id_ctrl_opcode_4_port, id_top_o(61) => 
                           s_id_ctrl_opcode_3_port, id_top_o(60) => 
                           s_id_ctrl_opcode_2_port, id_top_o(59) => 
                           s_id_ctrl_opcode_1_port, id_top_o(58) => 
                           s_id_ctrl_opcode_0_port, id_top_o(57) => 
                           s_id_out_RS_p_4_port, id_top_o(56) => 
                           s_id_out_RS_p_3_port, id_top_o(55) => 
                           s_id_out_RS_p_2_port, id_top_o(54) => 
                           s_id_out_RS_p_1_port, id_top_o(53) => 
                           s_id_out_RS_p_0_port, id_top_o(52) => 
                           s_id_out_RT_p_4_port, id_top_o(51) => 
                           s_id_out_RT_p_3_port, id_top_o(50) => 
                           s_id_out_RT_p_2_port, id_top_o(49) => 
                           s_id_out_RT_p_1_port, id_top_o(48) => 
                           s_id_out_RT_p_0_port, id_top_o(47) => 
                           s_id_out_RD_p_4_port, id_top_o(46) => 
                           s_id_out_RD_p_3_port, id_top_o(45) => 
                           s_id_out_RD_p_2_port, id_top_o(44) => 
                           s_id_out_RD_p_1_port, id_top_o(43) => 
                           s_id_out_RD_p_0_port, id_top_o(42) => 
                           s_id_out_shamt_p_4_port, id_top_o(41) => 
                           s_id_out_shamt_p_3_port, id_top_o(40) => 
                           s_id_out_shamt_p_2_port, id_top_o(39) => 
                           s_id_out_shamt_p_1_port, id_top_o(38) => 
                           s_id_out_shamt_p_0_port, id_top_o(37) => 
                           s_id_out_funct_p_5_port, id_top_o(36) => 
                           s_id_out_funct_p_4_port, id_top_o(35) => 
                           s_id_out_funct_p_3_port, id_top_o(34) => 
                           s_id_out_funct_p_2_port, id_top_o(33) => 
                           s_id_out_funct_p_1_port, id_top_o(32) => 
                           s_id_out_funct_p_0_port, id_top_o(31) => 
                           s_id_out_sign_extend_p_31_port, id_top_o(30) => 
                           s_id_out_sign_extend_p_30_port, id_top_o(29) => 
                           s_id_out_sign_extend_p_29_port, id_top_o(28) => 
                           s_id_out_sign_extend_p_28_port, id_top_o(27) => 
                           s_id_out_sign_extend_p_27_port, id_top_o(26) => 
                           s_id_out_sign_extend_p_26_port, id_top_o(25) => 
                           s_id_out_sign_extend_p_25_port, id_top_o(24) => 
                           s_id_out_sign_extend_p_24_port, id_top_o(23) => 
                           s_id_out_sign_extend_p_23_port, id_top_o(22) => 
                           s_id_out_sign_extend_p_22_port, id_top_o(21) => 
                           s_id_out_sign_extend_p_21_port, id_top_o(20) => 
                           s_id_out_sign_extend_p_20_port, id_top_o(19) => 
                           s_id_out_sign_extend_p_19_port, id_top_o(18) => 
                           s_id_out_sign_extend_p_18_port, id_top_o(17) => 
                           s_id_out_sign_extend_p_17_port, id_top_o(16) => 
                           s_id_out_sign_extend_p_16_port, id_top_o(15) => 
                           s_id_out_sign_extend_p_15_port, id_top_o(14) => 
                           s_id_out_sign_extend_p_14_port, id_top_o(13) => 
                           s_id_out_sign_extend_p_13_port, id_top_o(12) => 
                           s_id_out_sign_extend_p_12_port, id_top_o(11) => 
                           s_id_out_sign_extend_p_11_port, id_top_o(10) => 
                           s_id_out_sign_extend_p_10_port, id_top_o(9) => 
                           s_id_out_sign_extend_p_9_port, id_top_o(8) => 
                           s_id_out_sign_extend_p_8_port, id_top_o(7) => 
                           s_id_out_sign_extend_p_7_port, id_top_o(6) => 
                           s_id_out_sign_extend_p_6_port, id_top_o(5) => 
                           s_id_out_sign_extend_p_5_port, id_top_o(4) => 
                           s_id_out_sign_extend_p_4_port, id_top_o(3) => 
                           s_id_out_sign_extend_p_3_port, id_top_o(2) => 
                           s_id_out_sign_extend_p_2_port, id_top_o(1) => 
                           s_id_out_sign_extend_p_1_port, id_top_o(0) => 
                           s_id_out_sign_extend_p_0_port);
   id_exe_inst : id_exe port map( clk => clk, rst_n => n34, halt_i => 
                           X_Logic0_port, ID_EXE_i(142) => 
                           s_id_out_regA_p_31_port, ID_EXE_i(141) => 
                           s_id_out_regA_p_30_port, ID_EXE_i(140) => 
                           s_id_out_regA_p_29_port, ID_EXE_i(139) => 
                           s_id_out_regA_p_28_port, ID_EXE_i(138) => 
                           s_id_out_regA_p_27_port, ID_EXE_i(137) => 
                           s_id_out_regA_p_26_port, ID_EXE_i(136) => 
                           s_id_out_regA_p_25_port, ID_EXE_i(135) => 
                           s_id_out_regA_p_24_port, ID_EXE_i(134) => 
                           s_id_out_regA_p_23_port, ID_EXE_i(133) => 
                           s_id_out_regA_p_22_port, ID_EXE_i(132) => 
                           s_id_out_regA_p_21_port, ID_EXE_i(131) => 
                           s_id_out_regA_p_20_port, ID_EXE_i(130) => 
                           s_id_out_regA_p_19_port, ID_EXE_i(129) => 
                           s_id_out_regA_p_18_port, ID_EXE_i(128) => 
                           s_id_out_regA_p_17_port, ID_EXE_i(127) => 
                           s_id_out_regA_p_16_port, ID_EXE_i(126) => 
                           s_id_out_regA_p_15_port, ID_EXE_i(125) => 
                           s_id_out_regA_p_14_port, ID_EXE_i(124) => 
                           s_id_out_regA_p_13_port, ID_EXE_i(123) => 
                           s_id_out_regA_p_12_port, ID_EXE_i(122) => 
                           s_id_out_regA_p_11_port, ID_EXE_i(121) => 
                           s_id_out_regA_p_10_port, ID_EXE_i(120) => 
                           s_id_out_regA_p_9_port, ID_EXE_i(119) => 
                           s_id_out_regA_p_8_port, ID_EXE_i(118) => 
                           s_id_out_regA_p_7_port, ID_EXE_i(117) => 
                           s_id_out_regA_p_6_port, ID_EXE_i(116) => 
                           s_id_out_regA_p_5_port, ID_EXE_i(115) => 
                           s_id_out_regA_p_4_port, ID_EXE_i(114) => 
                           s_id_out_regA_p_3_port, ID_EXE_i(113) => 
                           s_id_out_regA_p_2_port, ID_EXE_i(112) => 
                           s_id_out_regA_p_1_port, ID_EXE_i(111) => 
                           s_id_out_regA_p_0_port, ID_EXE_i(110) => 
                           s_id_out_regB_p_31_port, ID_EXE_i(109) => 
                           s_id_out_regB_p_30_port, ID_EXE_i(108) => 
                           s_id_out_regB_p_29_port, ID_EXE_i(107) => 
                           s_id_out_regB_p_28_port, ID_EXE_i(106) => 
                           s_id_out_regB_p_27_port, ID_EXE_i(105) => 
                           s_id_out_regB_p_26_port, ID_EXE_i(104) => 
                           s_id_out_regB_p_25_port, ID_EXE_i(103) => 
                           s_id_out_regB_p_24_port, ID_EXE_i(102) => 
                           s_id_out_regB_p_23_port, ID_EXE_i(101) => 
                           s_id_out_regB_p_22_port, ID_EXE_i(100) => 
                           s_id_out_regB_p_21_port, ID_EXE_i(99) => 
                           s_id_out_regB_p_20_port, ID_EXE_i(98) => 
                           s_id_out_regB_p_19_port, ID_EXE_i(97) => 
                           s_id_out_regB_p_18_port, ID_EXE_i(96) => 
                           s_id_out_regB_p_17_port, ID_EXE_i(95) => 
                           s_id_out_regB_p_16_port, ID_EXE_i(94) => 
                           s_id_out_regB_p_15_port, ID_EXE_i(93) => 
                           s_id_out_regB_p_14_port, ID_EXE_i(92) => 
                           s_id_out_regB_p_13_port, ID_EXE_i(91) => 
                           s_id_out_regB_p_12_port, ID_EXE_i(90) => 
                           s_id_out_regB_p_11_port, ID_EXE_i(89) => 
                           s_id_out_regB_p_10_port, ID_EXE_i(88) => 
                           s_id_out_regB_p_9_port, ID_EXE_i(87) => 
                           s_id_out_regB_p_8_port, ID_EXE_i(86) => 
                           s_id_out_regB_p_7_port, ID_EXE_i(85) => 
                           s_id_out_regB_p_6_port, ID_EXE_i(84) => 
                           s_id_out_regB_p_5_port, ID_EXE_i(83) => 
                           s_id_out_regB_p_4_port, ID_EXE_i(82) => 
                           s_id_out_regB_p_3_port, ID_EXE_i(81) => 
                           s_id_out_regB_p_2_port, ID_EXE_i(80) => 
                           s_id_out_regB_p_1_port, ID_EXE_i(79) => 
                           s_id_out_regB_p_0_port, ID_EXE_i(78) => 
                           s_id_out_shamt_p_4_port, ID_EXE_i(77) => 
                           s_id_out_shamt_p_3_port, ID_EXE_i(76) => 
                           s_id_out_shamt_p_2_port, ID_EXE_i(75) => 
                           s_id_out_shamt_p_1_port, ID_EXE_i(74) => 
                           s_id_out_shamt_p_0_port, ID_EXE_i(73) => 
                           s_id_out_funct_p_5_port, ID_EXE_i(72) => 
                           s_id_out_funct_p_4_port, ID_EXE_i(71) => 
                           s_id_out_funct_p_3_port, ID_EXE_i(70) => 
                           s_id_out_funct_p_2_port, ID_EXE_i(69) => 
                           s_id_out_funct_p_1_port, ID_EXE_i(68) => 
                           s_id_out_funct_p_0_port, ID_EXE_i(67) => 
                           s_id_out_sign_extend_p_31_port, ID_EXE_i(66) => 
                           s_id_out_sign_extend_p_30_port, ID_EXE_i(65) => 
                           s_id_out_sign_extend_p_29_port, ID_EXE_i(64) => 
                           s_id_out_sign_extend_p_28_port, ID_EXE_i(63) => 
                           s_id_out_sign_extend_p_27_port, ID_EXE_i(62) => 
                           s_id_out_sign_extend_p_26_port, ID_EXE_i(61) => 
                           s_id_out_sign_extend_p_25_port, ID_EXE_i(60) => 
                           s_id_out_sign_extend_p_24_port, ID_EXE_i(59) => 
                           s_id_out_sign_extend_p_23_port, ID_EXE_i(58) => 
                           s_id_out_sign_extend_p_22_port, ID_EXE_i(57) => 
                           s_id_out_sign_extend_p_21_port, ID_EXE_i(56) => 
                           s_id_out_sign_extend_p_20_port, ID_EXE_i(55) => 
                           s_id_out_sign_extend_p_19_port, ID_EXE_i(54) => 
                           s_id_out_sign_extend_p_18_port, ID_EXE_i(53) => 
                           s_id_out_sign_extend_p_17_port, ID_EXE_i(52) => 
                           s_id_out_sign_extend_p_16_port, ID_EXE_i(51) => 
                           s_id_out_sign_extend_p_15_port, ID_EXE_i(50) => 
                           s_id_out_sign_extend_p_14_port, ID_EXE_i(49) => 
                           s_id_out_sign_extend_p_13_port, ID_EXE_i(48) => 
                           s_id_out_sign_extend_p_12_port, ID_EXE_i(47) => 
                           s_id_out_sign_extend_p_11_port, ID_EXE_i(46) => 
                           s_id_out_sign_extend_p_10_port, ID_EXE_i(45) => 
                           s_id_out_sign_extend_p_9_port, ID_EXE_i(44) => 
                           s_id_out_sign_extend_p_8_port, ID_EXE_i(43) => 
                           s_id_out_sign_extend_p_7_port, ID_EXE_i(42) => 
                           s_id_out_sign_extend_p_6_port, ID_EXE_i(41) => 
                           s_id_out_sign_extend_p_5_port, ID_EXE_i(40) => 
                           s_id_out_sign_extend_p_4_port, ID_EXE_i(39) => 
                           s_id_out_sign_extend_p_3_port, ID_EXE_i(38) => 
                           s_id_out_sign_extend_p_2_port, ID_EXE_i(37) => 
                           s_id_out_sign_extend_p_1_port, ID_EXE_i(36) => 
                           s_id_out_sign_extend_p_0_port, ID_EXE_i(35) => 
                           s_id_out_pc_plus1_p_11_port, ID_EXE_i(34) => 
                           s_id_out_pc_plus1_p_10_port, ID_EXE_i(33) => 
                           s_id_out_pc_plus1_p_9_port, ID_EXE_i(32) => 
                           s_id_out_pc_plus1_p_8_port, ID_EXE_i(31) => 
                           s_id_out_pc_plus1_p_7_port, ID_EXE_i(30) => 
                           s_id_out_pc_plus1_p_6_port, ID_EXE_i(29) => 
                           s_id_out_pc_plus1_p_5_port, ID_EXE_i(28) => 
                           s_id_out_pc_plus1_p_4_port, ID_EXE_i(27) => 
                           s_id_out_pc_plus1_p_3_port, ID_EXE_i(26) => 
                           s_id_out_pc_plus1_p_2_port, ID_EXE_i(25) => 
                           s_id_out_pc_plus1_p_1_port, ID_EXE_i(24) => 
                           s_id_out_pc_plus1_p_0_port, ID_EXE_i(23) => 
                           s_id_out_RS_p_4_port, ID_EXE_i(22) => 
                           s_id_out_RS_p_3_port, ID_EXE_i(21) => 
                           s_id_out_RS_p_2_port, ID_EXE_i(20) => 
                           s_id_out_RS_p_1_port, ID_EXE_i(19) => 
                           s_id_out_RS_p_0_port, ID_EXE_i(18) => 
                           s_id_out_RT_p_4_port, ID_EXE_i(17) => 
                           s_id_out_RT_p_3_port, ID_EXE_i(16) => 
                           s_id_out_RT_p_2_port, ID_EXE_i(15) => 
                           s_id_out_RT_p_1_port, ID_EXE_i(14) => 
                           s_id_out_RT_p_0_port, ID_EXE_i(13) => 
                           s_id_out_RD_p_4_port, ID_EXE_i(12) => 
                           s_id_out_RD_p_3_port, ID_EXE_i(11) => 
                           s_id_out_RD_p_2_port, ID_EXE_i(10) => 
                           s_id_out_RD_p_1_port, ID_EXE_i(9) => 
                           s_id_out_RD_p_0_port, ID_EXE_i(8) => 
                           s_ctrl_out_ALUsrc_B_p, ID_EXE_i(7) => 
                           s_ctrl_out_memtoReg_p, ID_EXE_i(6) => 
                           s_ctrl_out_regWrite_p, ID_EXE_i(5) => 
                           s_ctrl_out_memWen_n_p, ID_EXE_i(4) => 
                           s_ctrl_out_cALU_OP_p_3_port, ID_EXE_i(3) => 
                           s_ctrl_out_cALU_OP_p_2_port, ID_EXE_i(2) => 
                           s_ctrl_out_cALU_OP_p_1_port, ID_EXE_i(1) => 
                           s_ctrl_out_cALU_OP_p_0_port, ID_EXE_i(0) => 
                           s_ctrl_out_RegDst_p, ID_EXE_o(142) => 
                           s_exe_in_regA_p_31_port, ID_EXE_o(141) => 
                           s_exe_in_regA_p_30_port, ID_EXE_o(140) => 
                           s_exe_in_regA_p_29_port, ID_EXE_o(139) => 
                           s_exe_in_regA_p_28_port, ID_EXE_o(138) => 
                           s_exe_in_regA_p_27_port, ID_EXE_o(137) => 
                           s_exe_in_regA_p_26_port, ID_EXE_o(136) => 
                           s_exe_in_regA_p_25_port, ID_EXE_o(135) => 
                           s_exe_in_regA_p_24_port, ID_EXE_o(134) => 
                           s_exe_in_regA_p_23_port, ID_EXE_o(133) => 
                           s_exe_in_regA_p_22_port, ID_EXE_o(132) => 
                           s_exe_in_regA_p_21_port, ID_EXE_o(131) => 
                           s_exe_in_regA_p_20_port, ID_EXE_o(130) => 
                           s_exe_in_regA_p_19_port, ID_EXE_o(129) => 
                           s_exe_in_regA_p_18_port, ID_EXE_o(128) => 
                           s_exe_in_regA_p_17_port, ID_EXE_o(127) => 
                           s_exe_in_regA_p_16_port, ID_EXE_o(126) => 
                           s_exe_in_regA_p_15_port, ID_EXE_o(125) => 
                           s_exe_in_regA_p_14_port, ID_EXE_o(124) => 
                           s_exe_in_regA_p_13_port, ID_EXE_o(123) => 
                           s_exe_in_regA_p_12_port, ID_EXE_o(122) => 
                           s_exe_in_regA_p_11_port, ID_EXE_o(121) => 
                           s_exe_in_regA_p_10_port, ID_EXE_o(120) => 
                           s_exe_in_regA_p_9_port, ID_EXE_o(119) => 
                           s_exe_in_regA_p_8_port, ID_EXE_o(118) => 
                           s_exe_in_regA_p_7_port, ID_EXE_o(117) => 
                           s_exe_in_regA_p_6_port, ID_EXE_o(116) => 
                           s_exe_in_regA_p_5_port, ID_EXE_o(115) => 
                           s_exe_in_regA_p_4_port, ID_EXE_o(114) => 
                           s_exe_in_regA_p_3_port, ID_EXE_o(113) => 
                           s_exe_in_regA_p_2_port, ID_EXE_o(112) => 
                           s_exe_in_regA_p_1_port, ID_EXE_o(111) => 
                           s_exe_in_regA_p_0_port, ID_EXE_o(110) => 
                           s_exe_in_regB_p_31_port, ID_EXE_o(109) => 
                           s_exe_in_regB_p_30_port, ID_EXE_o(108) => 
                           s_exe_in_regB_p_29_port, ID_EXE_o(107) => 
                           s_exe_in_regB_p_28_port, ID_EXE_o(106) => 
                           s_exe_in_regB_p_27_port, ID_EXE_o(105) => 
                           s_exe_in_regB_p_26_port, ID_EXE_o(104) => 
                           s_exe_in_regB_p_25_port, ID_EXE_o(103) => 
                           s_exe_in_regB_p_24_port, ID_EXE_o(102) => 
                           s_exe_in_regB_p_23_port, ID_EXE_o(101) => 
                           s_exe_in_regB_p_22_port, ID_EXE_o(100) => 
                           s_exe_in_regB_p_21_port, ID_EXE_o(99) => 
                           s_exe_in_regB_p_20_port, ID_EXE_o(98) => 
                           s_exe_in_regB_p_19_port, ID_EXE_o(97) => 
                           s_exe_in_regB_p_18_port, ID_EXE_o(96) => 
                           s_exe_in_regB_p_17_port, ID_EXE_o(95) => 
                           s_exe_in_regB_p_16_port, ID_EXE_o(94) => 
                           s_exe_in_regB_p_15_port, ID_EXE_o(93) => 
                           s_exe_in_regB_p_14_port, ID_EXE_o(92) => 
                           s_exe_in_regB_p_13_port, ID_EXE_o(91) => 
                           s_exe_in_regB_p_12_port, ID_EXE_o(90) => 
                           s_exe_in_regB_p_11_port, ID_EXE_o(89) => 
                           s_exe_in_regB_p_10_port, ID_EXE_o(88) => 
                           s_exe_in_regB_p_9_port, ID_EXE_o(87) => 
                           s_exe_in_regB_p_8_port, ID_EXE_o(86) => 
                           s_exe_in_regB_p_7_port, ID_EXE_o(85) => 
                           s_exe_in_regB_p_6_port, ID_EXE_o(84) => 
                           s_exe_in_regB_p_5_port, ID_EXE_o(83) => 
                           s_exe_in_regB_p_4_port, ID_EXE_o(82) => 
                           s_exe_in_regB_p_3_port, ID_EXE_o(81) => 
                           s_exe_in_regB_p_2_port, ID_EXE_o(80) => 
                           s_exe_in_regB_p_1_port, ID_EXE_o(79) => 
                           s_exe_in_regB_p_0_port, ID_EXE_o(78) => 
                           s_exe_in_shamt_p_4_port, ID_EXE_o(77) => 
                           s_exe_in_shamt_p_3_port, ID_EXE_o(76) => 
                           s_exe_in_shamt_p_2_port, ID_EXE_o(75) => 
                           s_exe_in_shamt_p_1_port, ID_EXE_o(74) => 
                           s_exe_in_shamt_p_0_port, ID_EXE_o(73) => 
                           s_exe_in_funct_p_5_port, ID_EXE_o(72) => 
                           s_exe_in_funct_p_4_port, ID_EXE_o(71) => 
                           s_exe_in_funct_p_3_port, ID_EXE_o(70) => 
                           s_exe_in_funct_p_2_port, ID_EXE_o(69) => 
                           s_exe_in_funct_p_1_port, ID_EXE_o(68) => 
                           s_exe_in_funct_p_0_port, ID_EXE_o(67) => 
                           s_exe_in_sign_extend_p_31_port, ID_EXE_o(66) => 
                           s_exe_in_sign_extend_p_30_port, ID_EXE_o(65) => 
                           s_exe_in_sign_extend_p_29_port, ID_EXE_o(64) => 
                           s_exe_in_sign_extend_p_28_port, ID_EXE_o(63) => 
                           s_exe_in_sign_extend_p_27_port, ID_EXE_o(62) => 
                           s_exe_in_sign_extend_p_26_port, ID_EXE_o(61) => 
                           s_exe_in_sign_extend_p_25_port, ID_EXE_o(60) => 
                           s_exe_in_sign_extend_p_24_port, ID_EXE_o(59) => 
                           s_exe_in_sign_extend_p_23_port, ID_EXE_o(58) => 
                           s_exe_in_sign_extend_p_22_port, ID_EXE_o(57) => 
                           s_exe_in_sign_extend_p_21_port, ID_EXE_o(56) => 
                           s_exe_in_sign_extend_p_20_port, ID_EXE_o(55) => 
                           s_exe_in_sign_extend_p_19_port, ID_EXE_o(54) => 
                           s_exe_in_sign_extend_p_18_port, ID_EXE_o(53) => 
                           s_exe_in_sign_extend_p_17_port, ID_EXE_o(52) => 
                           s_exe_in_sign_extend_p_16_port, ID_EXE_o(51) => 
                           s_exe_in_sign_extend_p_15_port, ID_EXE_o(50) => 
                           s_exe_in_sign_extend_p_14_port, ID_EXE_o(49) => 
                           s_exe_in_sign_extend_p_13_port, ID_EXE_o(48) => 
                           s_exe_in_sign_extend_p_12_port, ID_EXE_o(47) => 
                           s_exe_in_sign_extend_p_11_port, ID_EXE_o(46) => 
                           s_exe_in_sign_extend_p_10_port, ID_EXE_o(45) => 
                           s_exe_in_sign_extend_p_9_port, ID_EXE_o(44) => 
                           s_exe_in_sign_extend_p_8_port, ID_EXE_o(43) => 
                           s_exe_in_sign_extend_p_7_port, ID_EXE_o(42) => 
                           s_exe_in_sign_extend_p_6_port, ID_EXE_o(41) => 
                           s_exe_in_sign_extend_p_5_port, ID_EXE_o(40) => 
                           s_exe_in_sign_extend_p_4_port, ID_EXE_o(39) => 
                           s_exe_in_sign_extend_p_3_port, ID_EXE_o(38) => 
                           s_exe_in_sign_extend_p_2_port, ID_EXE_o(37) => 
                           s_exe_in_sign_extend_p_1_port, ID_EXE_o(36) => 
                           s_exe_in_sign_extend_p_0_port, ID_EXE_o(35) => 
                           s_exe_in_pc_plus1_p_11_port, ID_EXE_o(34) => 
                           s_exe_in_pc_plus1_p_10_port, ID_EXE_o(33) => 
                           s_exe_in_pc_plus1_p_9_port, ID_EXE_o(32) => 
                           s_exe_in_pc_plus1_p_8_port, ID_EXE_o(31) => 
                           s_exe_in_pc_plus1_p_7_port, ID_EXE_o(30) => 
                           s_exe_in_pc_plus1_p_6_port, ID_EXE_o(29) => 
                           s_exe_in_pc_plus1_p_5_port, ID_EXE_o(28) => 
                           s_exe_in_pc_plus1_p_4_port, ID_EXE_o(27) => 
                           s_exe_in_pc_plus1_p_3_port, ID_EXE_o(26) => 
                           s_exe_in_pc_plus1_p_2_port, ID_EXE_o(25) => 
                           s_exe_in_pc_plus1_p_1_port, ID_EXE_o(24) => 
                           s_exe_in_pc_plus1_p_0_port, ID_EXE_o(23) => 
                           s_exe_in_RS_p_4_port, ID_EXE_o(22) => 
                           s_exe_in_RS_p_3_port, ID_EXE_o(21) => 
                           s_exe_in_RS_p_2_port, ID_EXE_o(20) => 
                           s_exe_in_RS_p_1_port, ID_EXE_o(19) => 
                           s_exe_in_RS_p_0_port, ID_EXE_o(18) => 
                           s_exe_in_RT_p_4_port, ID_EXE_o(17) => 
                           s_exe_in_RT_p_3_port, ID_EXE_o(16) => 
                           s_exe_in_RT_p_2_port, ID_EXE_o(15) => 
                           s_exe_in_RT_p_1_port, ID_EXE_o(14) => 
                           s_exe_in_RT_p_0_port, ID_EXE_o(13) => 
                           s_exe_in_RD_p_4_port, ID_EXE_o(12) => 
                           s_exe_in_RD_p_3_port, ID_EXE_o(11) => 
                           s_exe_in_RD_p_2_port, ID_EXE_o(10) => 
                           s_exe_in_RD_p_1_port, ID_EXE_o(9) => 
                           s_exe_in_RD_p_0_port, ID_EXE_o(8) => 
                           s_exe_in_ALUsrc_B_p, ID_EXE_o(7) => 
                           s_exe_out_memtoReg_p, ID_EXE_o(6) => 
                           s_exe_out_regWrite_p, ID_EXE_o(5) => 
                           s_exe_out_memWen_n_p, ID_EXE_o(4) => 
                           s_exe_in_cALU_OP_p_3_port, ID_EXE_o(3) => 
                           s_exe_in_cALU_OP_p_2_port, ID_EXE_o(2) => 
                           s_exe_in_cALU_OP_p_1_port, ID_EXE_o(1) => 
                           s_exe_in_cALU_OP_p_0_port, ID_EXE_o(0) => 
                           s_exe_in_RegDst_p);
   exe_top_inst : exe_top port map( clk => clk, rst_n => n33, exe_top_i(134) =>
                           s_exe_in_shamt_p_4_port, exe_top_i(133) => 
                           s_exe_in_shamt_p_3_port, exe_top_i(132) => 
                           s_exe_in_shamt_p_2_port, exe_top_i(131) => 
                           s_exe_in_shamt_p_1_port, exe_top_i(130) => 
                           s_exe_in_shamt_p_0_port, exe_top_i(129) => 
                           s_src_a_31_port, exe_top_i(128) => s_src_a_30_port, 
                           exe_top_i(127) => s_src_a_29_port, exe_top_i(126) =>
                           s_src_a_28_port, exe_top_i(125) => s_src_a_27_port, 
                           exe_top_i(124) => s_src_a_26_port, exe_top_i(123) =>
                           s_src_a_25_port, exe_top_i(122) => s_src_a_24_port, 
                           exe_top_i(121) => s_src_a_23_port, exe_top_i(120) =>
                           s_src_a_22_port, exe_top_i(119) => s_src_a_21_port, 
                           exe_top_i(118) => s_src_a_20_port, exe_top_i(117) =>
                           s_src_a_19_port, exe_top_i(116) => s_src_a_18_port, 
                           exe_top_i(115) => s_src_a_17_port, exe_top_i(114) =>
                           s_src_a_16_port, exe_top_i(113) => s_src_a_15_port, 
                           exe_top_i(112) => s_src_a_14_port, exe_top_i(111) =>
                           s_src_a_13_port, exe_top_i(110) => s_src_a_12_port, 
                           exe_top_i(109) => s_src_a_11_port, exe_top_i(108) =>
                           s_src_a_10_port, exe_top_i(107) => s_src_a_9_port, 
                           exe_top_i(106) => s_src_a_8_port, exe_top_i(105) => 
                           s_src_a_7_port, exe_top_i(104) => s_src_a_6_port, 
                           exe_top_i(103) => s_src_a_5_port, exe_top_i(102) => 
                           s_src_a_4_port, exe_top_i(101) => s_src_a_3_port, 
                           exe_top_i(100) => s_src_a_2_port, exe_top_i(99) => 
                           s_src_a_1_port, exe_top_i(98) => s_src_a_0_port, 
                           exe_top_i(97) => s_src_b_31_port, exe_top_i(96) => 
                           s_src_b_30_port, exe_top_i(95) => s_src_b_29_port, 
                           exe_top_i(94) => s_src_b_28_port, exe_top_i(93) => 
                           s_src_b_27_port, exe_top_i(92) => s_src_b_26_port, 
                           exe_top_i(91) => s_src_b_25_port, exe_top_i(90) => 
                           s_src_b_24_port, exe_top_i(89) => s_src_b_23_port, 
                           exe_top_i(88) => s_src_b_22_port, exe_top_i(87) => 
                           s_src_b_21_port, exe_top_i(86) => s_src_b_20_port, 
                           exe_top_i(85) => s_src_b_19_port, exe_top_i(84) => 
                           s_src_b_18_port, exe_top_i(83) => s_src_b_17_port, 
                           exe_top_i(82) => s_src_b_16_port, exe_top_i(81) => 
                           s_src_b_15_port, exe_top_i(80) => s_src_b_14_port, 
                           exe_top_i(79) => s_src_b_13_port, exe_top_i(78) => 
                           s_src_b_12_port, exe_top_i(77) => s_src_b_11_port, 
                           exe_top_i(76) => s_src_b_10_port, exe_top_i(75) => 
                           s_src_b_9_port, exe_top_i(74) => s_src_b_8_port, 
                           exe_top_i(73) => s_src_b_7_port, exe_top_i(72) => 
                           s_src_b_6_port, exe_top_i(71) => s_src_b_5_port, 
                           exe_top_i(70) => s_src_b_4_port, exe_top_i(69) => 
                           s_src_b_3_port, exe_top_i(68) => s_src_b_2_port, 
                           exe_top_i(67) => s_src_b_1_port, exe_top_i(66) => 
                           s_src_b_0_port, exe_top_i(65) => s_exe_in_ALUsrc_B_p
                           , exe_top_i(64) => s_exe_in_sign_extend_p_31_port, 
                           exe_top_i(63) => s_exe_in_sign_extend_p_30_port, 
                           exe_top_i(62) => s_exe_in_sign_extend_p_29_port, 
                           exe_top_i(61) => s_exe_in_sign_extend_p_28_port, 
                           exe_top_i(60) => s_exe_in_sign_extend_p_27_port, 
                           exe_top_i(59) => s_exe_in_sign_extend_p_26_port, 
                           exe_top_i(58) => s_exe_in_sign_extend_p_25_port, 
                           exe_top_i(57) => s_exe_in_sign_extend_p_24_port, 
                           exe_top_i(56) => s_exe_in_sign_extend_p_23_port, 
                           exe_top_i(55) => s_exe_in_sign_extend_p_22_port, 
                           exe_top_i(54) => s_exe_in_sign_extend_p_21_port, 
                           exe_top_i(53) => s_exe_in_sign_extend_p_20_port, 
                           exe_top_i(52) => s_exe_in_sign_extend_p_19_port, 
                           exe_top_i(51) => s_exe_in_sign_extend_p_18_port, 
                           exe_top_i(50) => s_exe_in_sign_extend_p_17_port, 
                           exe_top_i(49) => s_exe_in_sign_extend_p_16_port, 
                           exe_top_i(48) => s_exe_in_sign_extend_p_15_port, 
                           exe_top_i(47) => s_exe_in_sign_extend_p_14_port, 
                           exe_top_i(46) => s_exe_in_sign_extend_p_13_port, 
                           exe_top_i(45) => s_exe_in_sign_extend_p_12_port, 
                           exe_top_i(44) => s_exe_in_sign_extend_p_11_port, 
                           exe_top_i(43) => s_exe_in_sign_extend_p_10_port, 
                           exe_top_i(42) => s_exe_in_sign_extend_p_9_port, 
                           exe_top_i(41) => s_exe_in_sign_extend_p_8_port, 
                           exe_top_i(40) => s_exe_in_sign_extend_p_7_port, 
                           exe_top_i(39) => s_exe_in_sign_extend_p_6_port, 
                           exe_top_i(38) => s_exe_in_sign_extend_p_5_port, 
                           exe_top_i(37) => s_exe_in_sign_extend_p_4_port, 
                           exe_top_i(36) => s_exe_in_sign_extend_p_3_port, 
                           exe_top_i(35) => s_exe_in_sign_extend_p_2_port, 
                           exe_top_i(34) => s_exe_in_sign_extend_p_1_port, 
                           exe_top_i(33) => s_exe_in_sign_extend_p_0_port, 
                           exe_top_i(32) => s_exe_in_cALU_OP_p_3_port, 
                           exe_top_i(31) => s_exe_in_cALU_OP_p_2_port, 
                           exe_top_i(30) => s_exe_in_cALU_OP_p_1_port, 
                           exe_top_i(29) => s_exe_in_cALU_OP_p_0_port, 
                           exe_top_i(28) => s_exe_in_funct_p_5_port, 
                           exe_top_i(27) => s_exe_in_funct_p_4_port, 
                           exe_top_i(26) => s_exe_in_funct_p_3_port, 
                           exe_top_i(25) => s_exe_in_funct_p_2_port, 
                           exe_top_i(24) => s_exe_in_funct_p_1_port, 
                           exe_top_i(23) => s_exe_in_funct_p_0_port, 
                           exe_top_i(22) => s_exe_in_pc_plus1_p_11_port, 
                           exe_top_i(21) => s_exe_in_pc_plus1_p_10_port, 
                           exe_top_i(20) => s_exe_in_pc_plus1_p_9_port, 
                           exe_top_i(19) => s_exe_in_pc_plus1_p_8_port, 
                           exe_top_i(18) => s_exe_in_pc_plus1_p_7_port, 
                           exe_top_i(17) => s_exe_in_pc_plus1_p_6_port, 
                           exe_top_i(16) => s_exe_in_pc_plus1_p_5_port, 
                           exe_top_i(15) => s_exe_in_pc_plus1_p_4_port, 
                           exe_top_i(14) => s_exe_in_pc_plus1_p_3_port, 
                           exe_top_i(13) => s_exe_in_pc_plus1_p_2_port, 
                           exe_top_i(12) => s_exe_in_pc_plus1_p_1_port, 
                           exe_top_i(11) => s_exe_in_pc_plus1_p_0_port, 
                           exe_top_i(10) => s_exe_in_RegDst_p, exe_top_i(9) => 
                           s_exe_in_RT_p_4_port, exe_top_i(8) => 
                           s_exe_in_RT_p_3_port, exe_top_i(7) => 
                           s_exe_in_RT_p_2_port, exe_top_i(6) => 
                           s_exe_in_RT_p_1_port, exe_top_i(5) => 
                           s_exe_in_RT_p_0_port, exe_top_i(4) => 
                           s_exe_in_RD_p_4_port, exe_top_i(3) => 
                           s_exe_in_RD_p_3_port, exe_top_i(2) => 
                           s_exe_in_RD_p_2_port, exe_top_i(1) => 
                           s_exe_in_RD_p_1_port, exe_top_i(0) => 
                           s_exe_in_RD_p_0_port, exe_top_o(81) => s_if_PCSrc, 
                           exe_top_o(80) => s_exe_if_branch_pc_11_port, 
                           exe_top_o(79) => s_exe_if_branch_pc_10_port, 
                           exe_top_o(78) => s_exe_if_branch_pc_9_port, 
                           exe_top_o(77) => s_exe_if_branch_pc_8_port, 
                           exe_top_o(76) => s_exe_if_branch_pc_7_port, 
                           exe_top_o(75) => s_exe_if_branch_pc_6_port, 
                           exe_top_o(74) => s_exe_if_branch_pc_5_port, 
                           exe_top_o(73) => s_exe_if_branch_pc_4_port, 
                           exe_top_o(72) => s_exe_if_branch_pc_3_port, 
                           exe_top_o(71) => s_exe_if_branch_pc_2_port, 
                           exe_top_o(70) => s_exe_if_branch_pc_1_port, 
                           exe_top_o(69) => s_exe_if_branch_pc_0_port, 
                           exe_top_o(68) => s_exe_out_alu_res_p_31_port, 
                           exe_top_o(67) => s_exe_out_alu_res_p_30_port, 
                           exe_top_o(66) => s_exe_out_alu_res_p_29_port, 
                           exe_top_o(65) => s_exe_out_alu_res_p_28_port, 
                           exe_top_o(64) => s_exe_out_alu_res_p_27_port, 
                           exe_top_o(63) => s_exe_out_alu_res_p_26_port, 
                           exe_top_o(62) => s_exe_out_alu_res_p_25_port, 
                           exe_top_o(61) => s_exe_out_alu_res_p_24_port, 
                           exe_top_o(60) => s_exe_out_alu_res_p_23_port, 
                           exe_top_o(59) => s_exe_out_alu_res_p_22_port, 
                           exe_top_o(58) => s_exe_out_alu_res_p_21_port, 
                           exe_top_o(57) => s_exe_out_alu_res_p_20_port, 
                           exe_top_o(56) => s_exe_out_alu_res_p_19_port, 
                           exe_top_o(55) => s_exe_out_alu_res_p_18_port, 
                           exe_top_o(54) => s_exe_out_alu_res_p_17_port, 
                           exe_top_o(53) => s_exe_out_alu_res_p_16_port, 
                           exe_top_o(52) => s_exe_out_alu_res_p_15_port, 
                           exe_top_o(51) => s_exe_out_alu_res_p_14_port, 
                           exe_top_o(50) => s_exe_out_alu_res_p_13_port, 
                           exe_top_o(49) => s_exe_out_alu_res_p_12_port, 
                           exe_top_o(48) => s_exe_out_alu_res_p_11_port, 
                           exe_top_o(47) => s_exe_out_alu_res_p_10_port, 
                           exe_top_o(46) => s_exe_out_alu_res_p_9_port, 
                           exe_top_o(45) => s_exe_out_alu_res_p_8_port, 
                           exe_top_o(44) => s_exe_out_alu_res_p_7_port, 
                           exe_top_o(43) => s_exe_out_alu_res_p_6_port, 
                           exe_top_o(42) => s_exe_out_alu_res_p_5_port, 
                           exe_top_o(41) => s_exe_out_alu_res_p_4_port, 
                           exe_top_o(40) => s_exe_out_alu_res_p_3_port, 
                           exe_top_o(39) => s_exe_out_alu_res_p_2_port, 
                           exe_top_o(38) => s_exe_out_alu_res_p_1_port, 
                           exe_top_o(37) => s_exe_out_alu_res_p_0_port, 
                           exe_top_o(36) => s_exe_out_write_reg_p_4_port, 
                           exe_top_o(35) => s_exe_out_write_reg_p_3_port, 
                           exe_top_o(34) => s_exe_out_write_reg_p_2_port, 
                           exe_top_o(33) => s_exe_out_write_reg_p_1_port, 
                           exe_top_o(32) => s_exe_out_write_reg_p_0_port, 
                           exe_top_o(31) => s_exe_out_dmem_data_p_31_port, 
                           exe_top_o(30) => s_exe_out_dmem_data_p_30_port, 
                           exe_top_o(29) => s_exe_out_dmem_data_p_29_port, 
                           exe_top_o(28) => s_exe_out_dmem_data_p_28_port, 
                           exe_top_o(27) => s_exe_out_dmem_data_p_27_port, 
                           exe_top_o(26) => s_exe_out_dmem_data_p_26_port, 
                           exe_top_o(25) => s_exe_out_dmem_data_p_25_port, 
                           exe_top_o(24) => s_exe_out_dmem_data_p_24_port, 
                           exe_top_o(23) => s_exe_out_dmem_data_p_23_port, 
                           exe_top_o(22) => s_exe_out_dmem_data_p_22_port, 
                           exe_top_o(21) => s_exe_out_dmem_data_p_21_port, 
                           exe_top_o(20) => s_exe_out_dmem_data_p_20_port, 
                           exe_top_o(19) => s_exe_out_dmem_data_p_19_port, 
                           exe_top_o(18) => s_exe_out_dmem_data_p_18_port, 
                           exe_top_o(17) => s_exe_out_dmem_data_p_17_port, 
                           exe_top_o(16) => s_exe_out_dmem_data_p_16_port, 
                           exe_top_o(15) => s_exe_out_dmem_data_p_15_port, 
                           exe_top_o(14) => s_exe_out_dmem_data_p_14_port, 
                           exe_top_o(13) => s_exe_out_dmem_data_p_13_port, 
                           exe_top_o(12) => s_exe_out_dmem_data_p_12_port, 
                           exe_top_o(11) => s_exe_out_dmem_data_p_11_port, 
                           exe_top_o(10) => s_exe_out_dmem_data_p_10_port, 
                           exe_top_o(9) => s_exe_out_dmem_data_p_9_port, 
                           exe_top_o(8) => s_exe_out_dmem_data_p_8_port, 
                           exe_top_o(7) => s_exe_out_dmem_data_p_7_port, 
                           exe_top_o(6) => s_exe_out_dmem_data_p_6_port, 
                           exe_top_o(5) => s_exe_out_dmem_data_p_5_port, 
                           exe_top_o(4) => s_exe_out_dmem_data_p_4_port, 
                           exe_top_o(3) => s_exe_out_dmem_data_p_3_port, 
                           exe_top_o(2) => s_exe_out_dmem_data_p_2_port, 
                           exe_top_o(1) => s_exe_out_dmem_data_p_1_port, 
                           exe_top_o(0) => s_exe_out_dmem_data_p_0_port);
   forwarding_unit_inst : forwarding_unit port map( forwarding_unit_i(31) => 
                           s_exe_in_RS_p_4_port, forwarding_unit_i(30) => 
                           s_exe_in_RS_p_3_port, forwarding_unit_i(29) => 
                           s_exe_in_RS_p_2_port, forwarding_unit_i(28) => 
                           s_exe_in_RS_p_1_port, forwarding_unit_i(27) => 
                           s_exe_in_RS_p_0_port, forwarding_unit_i(26) => 
                           s_exe_in_RT_p_4_port, forwarding_unit_i(25) => 
                           s_exe_in_RT_p_3_port, forwarding_unit_i(24) => 
                           s_exe_in_RT_p_2_port, forwarding_unit_i(23) => 
                           s_exe_in_RT_p_1_port, forwarding_unit_i(22) => 
                           s_exe_in_RT_p_0_port, forwarding_unit_i(21) => 
                           s_id_out_RS_p_4_port, forwarding_unit_i(20) => 
                           s_id_out_RS_p_3_port, forwarding_unit_i(19) => 
                           s_id_out_RS_p_2_port, forwarding_unit_i(18) => 
                           s_id_out_RS_p_1_port, forwarding_unit_i(17) => 
                           s_id_out_RS_p_0_port, forwarding_unit_i(16) => 
                           s_id_out_RT_p_4_port, forwarding_unit_i(15) => 
                           s_id_out_RT_p_3_port, forwarding_unit_i(14) => 
                           s_id_out_RT_p_2_port, forwarding_unit_i(13) => 
                           s_id_out_RT_p_1_port, forwarding_unit_i(12) => 
                           s_id_out_RT_p_0_port, forwarding_unit_i(11) => 
                           s_mem_out_write_reg_p_4_port, forwarding_unit_i(10) 
                           => s_mem_out_write_reg_p_3_port, 
                           forwarding_unit_i(9) => s_mem_out_write_reg_p_2_port
                           , forwarding_unit_i(8) => 
                           s_mem_out_write_reg_p_1_port, forwarding_unit_i(7) 
                           => s_mem_out_write_reg_p_0_port, 
                           forwarding_unit_i(6) => s_wb_in_write_reg_p_4_port, 
                           forwarding_unit_i(5) => s_wb_in_write_reg_p_3_port, 
                           forwarding_unit_i(4) => s_wb_in_write_reg_p_2_port, 
                           forwarding_unit_i(3) => s_wb_in_write_reg_p_1_port, 
                           forwarding_unit_i(2) => s_wb_in_write_reg_p_0_port, 
                           forwarding_unit_i(1) => s_mem_out_regWrite_p, 
                           forwarding_unit_i(0) => s_wb_in_regWrite_p, 
                           forwarding_unit_o(5) => s_forward_A_1_port, 
                           forwarding_unit_o(4) => s_forward_A_0_port, 
                           forwarding_unit_o(3) => s_forward_B_1_port, 
                           forwarding_unit_o(2) => s_forward_B_0_port, 
                           forwarding_unit_o(1) => s_regfile_forward_A, 
                           forwarding_unit_o(0) => s_regfile_forward_B);
   exe_mem_inst : exe_mem port map( clk => clk, rst_n => n33, halt_i => 
                           X_Logic0_port, EXE_MEM_i(71) => 
                           s_exe_out_alu_res_p_31_port, EXE_MEM_i(70) => 
                           s_exe_out_alu_res_p_30_port, EXE_MEM_i(69) => 
                           s_exe_out_alu_res_p_29_port, EXE_MEM_i(68) => 
                           s_exe_out_alu_res_p_28_port, EXE_MEM_i(67) => 
                           s_exe_out_alu_res_p_27_port, EXE_MEM_i(66) => 
                           s_exe_out_alu_res_p_26_port, EXE_MEM_i(65) => 
                           s_exe_out_alu_res_p_25_port, EXE_MEM_i(64) => 
                           s_exe_out_alu_res_p_24_port, EXE_MEM_i(63) => 
                           s_exe_out_alu_res_p_23_port, EXE_MEM_i(62) => 
                           s_exe_out_alu_res_p_22_port, EXE_MEM_i(61) => 
                           s_exe_out_alu_res_p_21_port, EXE_MEM_i(60) => 
                           s_exe_out_alu_res_p_20_port, EXE_MEM_i(59) => 
                           s_exe_out_alu_res_p_19_port, EXE_MEM_i(58) => 
                           s_exe_out_alu_res_p_18_port, EXE_MEM_i(57) => 
                           s_exe_out_alu_res_p_17_port, EXE_MEM_i(56) => 
                           s_exe_out_alu_res_p_16_port, EXE_MEM_i(55) => 
                           s_exe_out_alu_res_p_15_port, EXE_MEM_i(54) => 
                           s_exe_out_alu_res_p_14_port, EXE_MEM_i(53) => 
                           s_exe_out_alu_res_p_13_port, EXE_MEM_i(52) => 
                           s_exe_out_alu_res_p_12_port, EXE_MEM_i(51) => 
                           s_exe_out_alu_res_p_11_port, EXE_MEM_i(50) => 
                           s_exe_out_alu_res_p_10_port, EXE_MEM_i(49) => 
                           s_exe_out_alu_res_p_9_port, EXE_MEM_i(48) => 
                           s_exe_out_alu_res_p_8_port, EXE_MEM_i(47) => 
                           s_exe_out_alu_res_p_7_port, EXE_MEM_i(46) => 
                           s_exe_out_alu_res_p_6_port, EXE_MEM_i(45) => 
                           s_exe_out_alu_res_p_5_port, EXE_MEM_i(44) => 
                           s_exe_out_alu_res_p_4_port, EXE_MEM_i(43) => 
                           s_exe_out_alu_res_p_3_port, EXE_MEM_i(42) => 
                           s_exe_out_alu_res_p_2_port, EXE_MEM_i(41) => 
                           s_exe_out_alu_res_p_1_port, EXE_MEM_i(40) => 
                           s_exe_out_alu_res_p_0_port, EXE_MEM_i(39) => 
                           s_exe_out_dmem_data_p_31_port, EXE_MEM_i(38) => 
                           s_exe_out_dmem_data_p_30_port, EXE_MEM_i(37) => 
                           s_exe_out_dmem_data_p_29_port, EXE_MEM_i(36) => 
                           s_exe_out_dmem_data_p_28_port, EXE_MEM_i(35) => 
                           s_exe_out_dmem_data_p_27_port, EXE_MEM_i(34) => 
                           s_exe_out_dmem_data_p_26_port, EXE_MEM_i(33) => 
                           s_exe_out_dmem_data_p_25_port, EXE_MEM_i(32) => 
                           s_exe_out_dmem_data_p_24_port, EXE_MEM_i(31) => 
                           s_exe_out_dmem_data_p_23_port, EXE_MEM_i(30) => 
                           s_exe_out_dmem_data_p_22_port, EXE_MEM_i(29) => 
                           s_exe_out_dmem_data_p_21_port, EXE_MEM_i(28) => 
                           s_exe_out_dmem_data_p_20_port, EXE_MEM_i(27) => 
                           s_exe_out_dmem_data_p_19_port, EXE_MEM_i(26) => 
                           s_exe_out_dmem_data_p_18_port, EXE_MEM_i(25) => 
                           s_exe_out_dmem_data_p_17_port, EXE_MEM_i(24) => 
                           s_exe_out_dmem_data_p_16_port, EXE_MEM_i(23) => 
                           s_exe_out_dmem_data_p_15_port, EXE_MEM_i(22) => 
                           s_exe_out_dmem_data_p_14_port, EXE_MEM_i(21) => 
                           s_exe_out_dmem_data_p_13_port, EXE_MEM_i(20) => 
                           s_exe_out_dmem_data_p_12_port, EXE_MEM_i(19) => 
                           s_exe_out_dmem_data_p_11_port, EXE_MEM_i(18) => 
                           s_exe_out_dmem_data_p_10_port, EXE_MEM_i(17) => 
                           s_exe_out_dmem_data_p_9_port, EXE_MEM_i(16) => 
                           s_exe_out_dmem_data_p_8_port, EXE_MEM_i(15) => 
                           s_exe_out_dmem_data_p_7_port, EXE_MEM_i(14) => 
                           s_exe_out_dmem_data_p_6_port, EXE_MEM_i(13) => 
                           s_exe_out_dmem_data_p_5_port, EXE_MEM_i(12) => 
                           s_exe_out_dmem_data_p_4_port, EXE_MEM_i(11) => 
                           s_exe_out_dmem_data_p_3_port, EXE_MEM_i(10) => 
                           s_exe_out_dmem_data_p_2_port, EXE_MEM_i(9) => 
                           s_exe_out_dmem_data_p_1_port, EXE_MEM_i(8) => 
                           s_exe_out_dmem_data_p_0_port, EXE_MEM_i(7) => 
                           s_exe_out_write_reg_p_4_port, EXE_MEM_i(6) => 
                           s_exe_out_write_reg_p_3_port, EXE_MEM_i(5) => 
                           s_exe_out_write_reg_p_2_port, EXE_MEM_i(4) => 
                           s_exe_out_write_reg_p_1_port, EXE_MEM_i(3) => 
                           s_exe_out_write_reg_p_0_port, EXE_MEM_i(2) => 
                           s_exe_out_memtoReg_p, EXE_MEM_i(1) => 
                           s_exe_out_regWrite_p, EXE_MEM_i(0) => 
                           s_exe_out_memWen_n_p, EXE_MEM_o(71) => 
                           s_mem_out_alu_res_p_31_port, EXE_MEM_o(70) => 
                           s_mem_out_alu_res_p_30_port, EXE_MEM_o(69) => 
                           s_mem_out_alu_res_p_29_port, EXE_MEM_o(68) => 
                           s_mem_out_alu_res_p_28_port, EXE_MEM_o(67) => 
                           s_mem_out_alu_res_p_27_port, EXE_MEM_o(66) => 
                           s_mem_out_alu_res_p_26_port, EXE_MEM_o(65) => 
                           s_mem_out_alu_res_p_25_port, EXE_MEM_o(64) => 
                           s_mem_out_alu_res_p_24_port, EXE_MEM_o(63) => 
                           s_mem_out_alu_res_p_23_port, EXE_MEM_o(62) => 
                           s_mem_out_alu_res_p_22_port, EXE_MEM_o(61) => 
                           s_mem_out_alu_res_p_21_port, EXE_MEM_o(60) => 
                           s_mem_out_alu_res_p_20_port, EXE_MEM_o(59) => 
                           s_mem_out_alu_res_p_19_port, EXE_MEM_o(58) => 
                           s_mem_out_alu_res_p_18_port, EXE_MEM_o(57) => 
                           s_mem_out_alu_res_p_17_port, EXE_MEM_o(56) => 
                           s_mem_out_alu_res_p_16_port, EXE_MEM_o(55) => 
                           s_mem_out_alu_res_p_15_port, EXE_MEM_o(54) => 
                           s_mem_out_alu_res_p_14_port, EXE_MEM_o(53) => 
                           s_mem_out_alu_res_p_13_port, EXE_MEM_o(52) => 
                           s_mem_out_alu_res_p_12_port, EXE_MEM_o(51) => 
                           mini_mips_o_DMEM_ADDR_11_port, EXE_MEM_o(50) => 
                           mini_mips_o_DMEM_ADDR_10_port, EXE_MEM_o(49) => 
                           mini_mips_o_DMEM_ADDR_9_port, EXE_MEM_o(48) => 
                           mini_mips_o_DMEM_ADDR_8_port, EXE_MEM_o(47) => 
                           mini_mips_o_DMEM_ADDR_7_port, EXE_MEM_o(46) => 
                           mini_mips_o_DMEM_ADDR_6_port, EXE_MEM_o(45) => 
                           mini_mips_o_DMEM_ADDR_5_port, EXE_MEM_o(44) => 
                           mini_mips_o_DMEM_ADDR_4_port, EXE_MEM_o(43) => 
                           mini_mips_o_DMEM_ADDR_3_port, EXE_MEM_o(42) => 
                           mini_mips_o_DMEM_ADDR_2_port, EXE_MEM_o(41) => 
                           mini_mips_o_DMEM_ADDR_1_port, EXE_MEM_o(40) => 
                           mini_mips_o_DMEM_ADDR_0_port, EXE_MEM_o(39) => 
                           mini_mips_o_DMEM_DATA_31_port, EXE_MEM_o(38) => 
                           mini_mips_o_DMEM_DATA_30_port, EXE_MEM_o(37) => 
                           mini_mips_o_DMEM_DATA_29_port, EXE_MEM_o(36) => 
                           mini_mips_o_DMEM_DATA_28_port, EXE_MEM_o(35) => 
                           mini_mips_o_DMEM_DATA_27_port, EXE_MEM_o(34) => 
                           mini_mips_o_DMEM_DATA_26_port, EXE_MEM_o(33) => 
                           mini_mips_o_DMEM_DATA_25_port, EXE_MEM_o(32) => 
                           mini_mips_o_DMEM_DATA_24_port, EXE_MEM_o(31) => 
                           mini_mips_o_DMEM_DATA_23_port, EXE_MEM_o(30) => 
                           mini_mips_o_DMEM_DATA_22_port, EXE_MEM_o(29) => 
                           mini_mips_o_DMEM_DATA_21_port, EXE_MEM_o(28) => 
                           mini_mips_o_DMEM_DATA_20_port, EXE_MEM_o(27) => 
                           mini_mips_o_DMEM_DATA_19_port, EXE_MEM_o(26) => 
                           mini_mips_o_DMEM_DATA_18_port, EXE_MEM_o(25) => 
                           mini_mips_o_DMEM_DATA_17_port, EXE_MEM_o(24) => 
                           mini_mips_o_DMEM_DATA_16_port, EXE_MEM_o(23) => 
                           mini_mips_o_DMEM_DATA_15_port, EXE_MEM_o(22) => 
                           mini_mips_o_DMEM_DATA_14_port, EXE_MEM_o(21) => 
                           mini_mips_o_DMEM_DATA_13_port, EXE_MEM_o(20) => 
                           mini_mips_o_DMEM_DATA_12_port, EXE_MEM_o(19) => 
                           mini_mips_o_DMEM_DATA_11_port, EXE_MEM_o(18) => 
                           mini_mips_o_DMEM_DATA_10_port, EXE_MEM_o(17) => 
                           mini_mips_o_DMEM_DATA_9_port, EXE_MEM_o(16) => 
                           mini_mips_o_DMEM_DATA_8_port, EXE_MEM_o(15) => 
                           mini_mips_o_DMEM_DATA_7_port, EXE_MEM_o(14) => 
                           mini_mips_o_DMEM_DATA_6_port, EXE_MEM_o(13) => 
                           mini_mips_o_DMEM_DATA_5_port, EXE_MEM_o(12) => 
                           mini_mips_o_DMEM_DATA_4_port, EXE_MEM_o(11) => 
                           mini_mips_o_DMEM_DATA_3_port, EXE_MEM_o(10) => 
                           mini_mips_o_DMEM_DATA_2_port, EXE_MEM_o(9) => 
                           mini_mips_o_DMEM_DATA_1_port, EXE_MEM_o(8) => 
                           mini_mips_o_DMEM_DATA_0_port, EXE_MEM_o(7) => 
                           s_mem_out_write_reg_p_4_port, EXE_MEM_o(6) => 
                           s_mem_out_write_reg_p_3_port, EXE_MEM_o(5) => 
                           s_mem_out_write_reg_p_2_port, EXE_MEM_o(4) => 
                           s_mem_out_write_reg_p_1_port, EXE_MEM_o(3) => 
                           s_mem_out_write_reg_p_0_port, EXE_MEM_o(2) => 
                           s_mem_out_memtoReg_p, EXE_MEM_o(1) => 
                           s_mem_out_regWrite_p, EXE_MEM_o(0) => 
                           mini_mips_o_DMEM_WEN_N_port);
   mem_wb_inst : mem_wb port map( clk => clk, rst_n => n34, halt_i => 
                           X_Logic0_port, MEM_WB_i(38) => 
                           s_mem_out_alu_res_p_31_port, MEM_WB_i(37) => 
                           s_mem_out_alu_res_p_30_port, MEM_WB_i(36) => 
                           s_mem_out_alu_res_p_29_port, MEM_WB_i(35) => 
                           s_mem_out_alu_res_p_28_port, MEM_WB_i(34) => 
                           s_mem_out_alu_res_p_27_port, MEM_WB_i(33) => 
                           s_mem_out_alu_res_p_26_port, MEM_WB_i(32) => 
                           s_mem_out_alu_res_p_25_port, MEM_WB_i(31) => 
                           s_mem_out_alu_res_p_24_port, MEM_WB_i(30) => 
                           s_mem_out_alu_res_p_23_port, MEM_WB_i(29) => 
                           s_mem_out_alu_res_p_22_port, MEM_WB_i(28) => 
                           s_mem_out_alu_res_p_21_port, MEM_WB_i(27) => 
                           s_mem_out_alu_res_p_20_port, MEM_WB_i(26) => 
                           s_mem_out_alu_res_p_19_port, MEM_WB_i(25) => 
                           s_mem_out_alu_res_p_18_port, MEM_WB_i(24) => 
                           s_mem_out_alu_res_p_17_port, MEM_WB_i(23) => 
                           s_mem_out_alu_res_p_16_port, MEM_WB_i(22) => 
                           s_mem_out_alu_res_p_15_port, MEM_WB_i(21) => 
                           s_mem_out_alu_res_p_14_port, MEM_WB_i(20) => 
                           s_mem_out_alu_res_p_13_port, MEM_WB_i(19) => 
                           s_mem_out_alu_res_p_12_port, MEM_WB_i(18) => 
                           mini_mips_o_DMEM_ADDR_11_port, MEM_WB_i(17) => 
                           mini_mips_o_DMEM_ADDR_10_port, MEM_WB_i(16) => 
                           mini_mips_o_DMEM_ADDR_9_port, MEM_WB_i(15) => 
                           mini_mips_o_DMEM_ADDR_8_port, MEM_WB_i(14) => 
                           mini_mips_o_DMEM_ADDR_7_port, MEM_WB_i(13) => 
                           mini_mips_o_DMEM_ADDR_6_port, MEM_WB_i(12) => 
                           mini_mips_o_DMEM_ADDR_5_port, MEM_WB_i(11) => 
                           mini_mips_o_DMEM_ADDR_4_port, MEM_WB_i(10) => 
                           mini_mips_o_DMEM_ADDR_3_port, MEM_WB_i(9) => 
                           mini_mips_o_DMEM_ADDR_2_port, MEM_WB_i(8) => 
                           mini_mips_o_DMEM_ADDR_1_port, MEM_WB_i(7) => 
                           mini_mips_o_DMEM_ADDR_0_port, MEM_WB_i(6) => 
                           s_mem_out_write_reg_p_4_port, MEM_WB_i(5) => 
                           s_mem_out_write_reg_p_3_port, MEM_WB_i(4) => 
                           s_mem_out_write_reg_p_2_port, MEM_WB_i(3) => 
                           s_mem_out_write_reg_p_1_port, MEM_WB_i(2) => 
                           s_mem_out_write_reg_p_0_port, MEM_WB_i(1) => 
                           s_mem_out_memtoReg_p, MEM_WB_i(0) => 
                           s_mem_out_regWrite_p, MEM_WB_o(38) => 
                           s_wb_in_alu_res_p_31_port, MEM_WB_o(37) => 
                           s_wb_in_alu_res_p_30_port, MEM_WB_o(36) => 
                           s_wb_in_alu_res_p_29_port, MEM_WB_o(35) => 
                           s_wb_in_alu_res_p_28_port, MEM_WB_o(34) => 
                           s_wb_in_alu_res_p_27_port, MEM_WB_o(33) => 
                           s_wb_in_alu_res_p_26_port, MEM_WB_o(32) => 
                           s_wb_in_alu_res_p_25_port, MEM_WB_o(31) => 
                           s_wb_in_alu_res_p_24_port, MEM_WB_o(30) => 
                           s_wb_in_alu_res_p_23_port, MEM_WB_o(29) => 
                           s_wb_in_alu_res_p_22_port, MEM_WB_o(28) => 
                           s_wb_in_alu_res_p_21_port, MEM_WB_o(27) => 
                           s_wb_in_alu_res_p_20_port, MEM_WB_o(26) => 
                           s_wb_in_alu_res_p_19_port, MEM_WB_o(25) => 
                           s_wb_in_alu_res_p_18_port, MEM_WB_o(24) => 
                           s_wb_in_alu_res_p_17_port, MEM_WB_o(23) => 
                           s_wb_in_alu_res_p_16_port, MEM_WB_o(22) => 
                           s_wb_in_alu_res_p_15_port, MEM_WB_o(21) => 
                           s_wb_in_alu_res_p_14_port, MEM_WB_o(20) => 
                           s_wb_in_alu_res_p_13_port, MEM_WB_o(19) => 
                           s_wb_in_alu_res_p_12_port, MEM_WB_o(18) => 
                           s_wb_in_alu_res_p_11_port, MEM_WB_o(17) => 
                           s_wb_in_alu_res_p_10_port, MEM_WB_o(16) => 
                           s_wb_in_alu_res_p_9_port, MEM_WB_o(15) => 
                           s_wb_in_alu_res_p_8_port, MEM_WB_o(14) => 
                           s_wb_in_alu_res_p_7_port, MEM_WB_o(13) => 
                           s_wb_in_alu_res_p_6_port, MEM_WB_o(12) => 
                           s_wb_in_alu_res_p_5_port, MEM_WB_o(11) => 
                           s_wb_in_alu_res_p_4_port, MEM_WB_o(10) => 
                           s_wb_in_alu_res_p_3_port, MEM_WB_o(9) => 
                           s_wb_in_alu_res_p_2_port, MEM_WB_o(8) => 
                           s_wb_in_alu_res_p_1_port, MEM_WB_o(7) => 
                           s_wb_in_alu_res_p_0_port, MEM_WB_o(6) => 
                           s_wb_in_write_reg_p_4_port, MEM_WB_o(5) => 
                           s_wb_in_write_reg_p_3_port, MEM_WB_o(4) => 
                           s_wb_in_write_reg_p_2_port, MEM_WB_o(3) => 
                           s_wb_in_write_reg_p_1_port, MEM_WB_o(2) => 
                           s_wb_in_write_reg_p_0_port, MEM_WB_o(1) => 
                           s_wb_in_memtoReg_p, MEM_WB_o(0) => 
                           s_wb_in_regWrite_p);
   U2 : HS65_LHS_XNOR2X6 port map( A => s_forward_A_0_port, B => 
                           s_forward_A_1_port, Z => n1);
   U3 : HS65_LHS_XNOR2X6 port map( A => s_forward_B_0_port, B => 
                           s_forward_B_1_port, Z => n2);
   U4 : HS65_LH_AND2X4 port map( A => s_forward_A_1_port, B => n36, Z => n9);
   U5 : HS65_LH_AND2X4 port map( A => s_forward_B_1_port, B => n37, Z => n6);
   U6 : HS65_LH_BFX9 port map( A => n9, Z => n5);
   U7 : HS65_LH_BFX9 port map( A => n9, Z => n8);
   U8 : HS65_LH_BFX9 port map( A => n13, Z => n15);
   U9 : HS65_LH_BFX9 port map( A => n1, Z => n11);
   U10 : HS65_LH_BFX9 port map( A => n1, Z => n12);
   U11 : HS65_LH_BFX9 port map( A => n31, Z => n29);
   U12 : HS65_LH_BFX9 port map( A => n9, Z => n3);
   U13 : HS65_LH_BFX9 port map( A => n6, Z => n17);
   U14 : HS65_LH_BFX9 port map( A => n6, Z => n18);
   U15 : HS65_LH_BFX9 port map( A => n6, Z => n19);
   U16 : HS65_LH_BFX9 port map( A => n13, Z => n14);
   U17 : HS65_LH_BFX9 port map( A => n23, Z => n24);
   U18 : HS65_LH_BFX9 port map( A => n23, Z => n25);
   U19 : HS65_LH_BFX9 port map( A => n1, Z => n10);
   U20 : HS65_LH_BFX9 port map( A => n2, Z => n20);
   U21 : HS65_LH_BFX9 port map( A => n2, Z => n21);
   U22 : HS65_LH_IVX9 port map( A => n28, Z => n27);
   U23 : HS65_LH_BFX9 port map( A => n23, Z => n26);
   U24 : HS65_LH_BFX9 port map( A => n13, Z => n16);
   U25 : HS65_LH_BFX9 port map( A => n2, Z => n22);
   U26 : HS65_LH_BFX9 port map( A => n31, Z => n30);
   U27 : HS65_LH_IVX9 port map( A => s_forward_A_0_port, Z => n36);
   U28 : HS65_LH_BFX9 port map( A => n7, Z => n13);
   U29 : HS65_LH_NOR2X6 port map( A => n36, B => s_forward_A_1_port, Z => n7);
   U30 : HS65_LH_IVX9 port map( A => s_forward_B_0_port, Z => n37);
   U31 : HS65_LH_BFX9 port map( A => n31, Z => n28);
   U32 : HS65_LH_IVX9 port map( A => s_wb_in_memtoReg_p, Z => n31);
   U33 : HS65_LH_BFX9 port map( A => n4, Z => n23);
   U34 : HS65_LH_NOR2X6 port map( A => n37, B => s_forward_B_1_port, Z => n4);
   U35 : HS65_LH_BFX9 port map( A => n32, Z => n33);
   U36 : HS65_LH_BFX9 port map( A => n32, Z => n34);
   U37 : HS65_LH_BFX9 port map( A => n32, Z => n35);
   U38 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_2_port, C =>
                           s_exe_in_regB_p_2_port, D => n21, E => 
                           mini_mips_o_DMEM_ADDR_2_port, F => n18, Z => 
                           s_src_b_2_port);
   U39 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_0_port, C =>
                           s_exe_in_regB_p_0_port, D => n20, E => 
                           mini_mips_o_DMEM_ADDR_0_port, F => n17, Z => 
                           s_src_b_0_port);
   U40 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_1_port, B => n29, C =>
                           mini_mips_i(33), D => n27, Z => 
                           s_writeback_data_1_port);
   U41 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_2_port, B => n30, C =>
                           mini_mips_i(34), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_2_port);
   U42 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_4_port, B => n30, C =>
                           mini_mips_i(36), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_4_port);
   U43 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_3_port, B => n30, C =>
                           mini_mips_i(35), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_3_port);
   U44 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_5_port, B => n30, C =>
                           mini_mips_i(37), D => n27, Z => 
                           s_writeback_data_5_port);
   U45 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_8_port, B => n30, C =>
                           mini_mips_i(40), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_8_port);
   U46 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_0_port, B => n28, C =>
                           mini_mips_i(32), D => n27, Z => 
                           s_writeback_data_0_port);
   U47 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_1_port, C =>
                           s_exe_in_regA_p_1_port, D => n10, E => n3, F => 
                           mini_mips_o_DMEM_ADDR_1_port, Z => s_src_a_1_port);
   U48 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_2_port, C =>
                           s_exe_in_regA_p_2_port, D => n11, E => n5, F => 
                           mini_mips_o_DMEM_ADDR_2_port, Z => s_src_a_2_port);
   U49 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_4_port, C =>
                           s_exe_in_regA_p_4_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_4_port, Z => s_src_a_4_port);
   U50 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_3_port, C =>
                           s_exe_in_regA_p_3_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_3_port, Z => s_src_a_3_port);
   U51 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_5_port, C =>
                           s_exe_in_regA_p_5_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_5_port, Z => s_src_a_5_port);
   U52 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_8_port, C =>
                           s_exe_in_regA_p_8_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_8_port, Z => s_src_a_8_port);
   U53 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_0_port, C =>
                           s_exe_in_regA_p_0_port, D => n10, E => n3, F => 
                           mini_mips_o_DMEM_ADDR_0_port, Z => s_src_a_0_port);
   U54 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_16_port, C 
                           => s_exe_in_regA_p_16_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_16_port, Z => s_src_a_16_port);
   U55 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_15_port, C 
                           => s_exe_in_regA_p_15_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_15_port, Z => s_src_a_15_port);
   U56 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_13_port, C 
                           => s_exe_in_regA_p_13_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_13_port, Z => s_src_a_13_port);
   U57 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_14_port, C 
                           => s_exe_in_regA_p_14_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_14_port, Z => s_src_a_14_port);
   U58 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_17_port, C 
                           => s_exe_in_regA_p_17_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_17_port, Z => s_src_a_17_port);
   U59 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_20_port, C 
                           => s_exe_in_regA_p_20_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_20_port, Z => s_src_a_20_port);
   U60 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_3_port, C =>
                           s_exe_in_regB_p_3_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_3_port, F => n19, Z => 
                           s_src_b_3_port);
   U61 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_1_port, C =>
                           s_exe_in_regB_p_1_port, D => n20, E => 
                           mini_mips_o_DMEM_ADDR_1_port, F => n17, Z => 
                           s_src_b_1_port);
   U62 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_4_port, C =>
                           s_exe_in_regB_p_4_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_4_port, F => n19, Z => 
                           s_src_b_4_port);
   U63 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_5_port, C =>
                           s_exe_in_regB_p_5_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_5_port, F => n19, Z => 
                           s_src_b_5_port);
   U64 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_6_port, C =>
                           s_exe_in_regB_p_6_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_6_port, F => n19, Z => 
                           s_src_b_6_port);
   U65 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_7_port, C =>
                           s_exe_in_regB_p_7_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_7_port, F => n19, Z => 
                           s_src_b_7_port);
   U66 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_8_port, C =>
                           s_exe_in_regB_p_8_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_8_port, F => n19, Z => 
                           s_src_b_8_port);
   U67 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_20_port, B => n29, C 
                           => mini_mips_i(52), D => n27, Z => 
                           s_writeback_data_20_port);
   U68 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_14_port, B => n29, C 
                           => mini_mips_i(46), D => n27, Z => 
                           s_writeback_data_14_port);
   U69 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_17_port, B => n29, C 
                           => mini_mips_i(49), D => n27, Z => 
                           s_writeback_data_17_port);
   U70 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_6_port, B => n30, C =>
                           mini_mips_i(38), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_6_port);
   U71 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_7_port, B => n30, C =>
                           mini_mips_i(39), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_7_port);
   U72 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_9_port, B => n30, C =>
                           s_wb_in_memtoReg_p, D => mini_mips_i(41), Z => 
                           s_writeback_data_9_port);
   U73 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_10_port, B => n29, C 
                           => mini_mips_i(42), D => n27, Z => 
                           s_writeback_data_10_port);
   U74 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_11_port, B => n29, C 
                           => mini_mips_i(43), D => n27, Z => 
                           s_writeback_data_11_port);
   U75 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_12_port, B => n29, C 
                           => mini_mips_i(44), D => n27, Z => 
                           s_writeback_data_12_port);
   U76 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_13_port, B => n29, C 
                           => mini_mips_i(45), D => n27, Z => 
                           s_writeback_data_13_port);
   U77 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_15_port, B => n29, C 
                           => mini_mips_i(47), D => n27, Z => 
                           s_writeback_data_15_port);
   U78 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_16_port, B => n29, C 
                           => mini_mips_i(48), D => n27, Z => 
                           s_writeback_data_16_port);
   U79 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_18_port, B => n29, C 
                           => mini_mips_i(50), D => n27, Z => 
                           s_writeback_data_18_port);
   U80 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_6_port, C =>
                           s_exe_in_regA_p_6_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_6_port, Z => s_src_a_6_port);
   U81 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_7_port, C =>
                           s_exe_in_regA_p_7_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_7_port, Z => s_src_a_7_port);
   U82 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_9_port, C =>
                           s_exe_in_regA_p_9_port, D => n12, E => n8, F => 
                           mini_mips_o_DMEM_ADDR_9_port, Z => s_src_a_9_port);
   U83 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_10_port, C 
                           => s_exe_in_regA_p_10_port, D => n10, E => n3, F => 
                           mini_mips_o_DMEM_ADDR_10_port, Z => s_src_a_10_port)
                           ;
   U84 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_11_port, C 
                           => s_exe_in_regA_p_11_port, D => n10, E => n3, F => 
                           mini_mips_o_DMEM_ADDR_11_port, Z => s_src_a_11_port)
                           ;
   U85 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_12_port, C 
                           => s_exe_in_regA_p_12_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_12_port, Z => s_src_a_12_port);
   U86 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_18_port, C 
                           => s_exe_in_regA_p_18_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_18_port, Z => s_src_a_18_port);
   U87 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_28_port, C 
                           => s_exe_in_regA_p_28_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_28_port, Z => s_src_a_28_port);
   U88 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_22_port, C 
                           => s_exe_in_regA_p_22_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_22_port, Z => s_src_a_22_port);
   U89 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_24_port, C 
                           => s_exe_in_regA_p_24_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_24_port, Z => s_src_a_24_port);
   U90 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_21_port, C 
                           => s_exe_in_regA_p_21_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_21_port, Z => s_src_a_21_port);
   U91 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_27_port, C 
                           => s_exe_in_regA_p_27_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_27_port, Z => s_src_a_27_port);
   U92 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_25_port, C 
                           => s_exe_in_regA_p_25_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_25_port, Z => s_src_a_25_port);
   U93 : HS65_LH_AO222X4 port map( A => n14, B => s_writeback_data_19_port, C 
                           => s_exe_in_regA_p_19_port, D => n10, E => n3, F => 
                           s_mem_out_alu_res_p_19_port, Z => s_src_a_19_port);
   U94 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_23_port, C 
                           => s_exe_in_regA_p_23_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_23_port, Z => s_src_a_23_port);
   U95 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_26_port, C 
                           => s_exe_in_regA_p_26_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_26_port, Z => s_src_a_26_port);
   U96 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_9_port, C =>
                           s_exe_in_regB_p_9_port, D => n22, E => 
                           mini_mips_o_DMEM_ADDR_9_port, F => n19, Z => 
                           s_src_b_9_port);
   U97 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_10_port, C 
                           => s_exe_in_regB_p_10_port, D => n20, E => 
                           mini_mips_o_DMEM_ADDR_10_port, F => n17, Z => 
                           s_src_b_10_port);
   U98 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_11_port, C 
                           => s_exe_in_regB_p_11_port, D => n20, E => 
                           mini_mips_o_DMEM_ADDR_11_port, F => n17, Z => 
                           s_src_b_11_port);
   U99 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_12_port, C 
                           => s_exe_in_regB_p_12_port, D => n20, E => 
                           s_mem_out_alu_res_p_12_port, F => n17, Z => 
                           s_src_b_12_port);
   U100 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_13_port, C 
                           => s_exe_in_regB_p_13_port, D => n20, E => 
                           s_mem_out_alu_res_p_13_port, F => n17, Z => 
                           s_src_b_13_port);
   U101 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_14_port, C 
                           => s_exe_in_regB_p_14_port, D => n20, E => 
                           s_mem_out_alu_res_p_14_port, F => n17, Z => 
                           s_src_b_14_port);
   U102 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_27_port, B => n29, C 
                           => mini_mips_i(59), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_27_port);
   U103 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_23_port, B => n29, C 
                           => mini_mips_i(55), D => n27, Z => 
                           s_writeback_data_23_port);
   U104 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_26_port, B => n29, C 
                           => mini_mips_i(58), D => n27, Z => 
                           s_writeback_data_26_port);
   U105 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_29_port, B => n30, C 
                           => mini_mips_i(61), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_29_port);
   U106 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_28_port, B => n29, C 
                           => mini_mips_i(60), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_28_port);
   U107 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_19_port, B => n29, C 
                           => mini_mips_i(51), D => n27, Z => 
                           s_writeback_data_19_port);
   U108 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_21_port, B => n29, C 
                           => mini_mips_i(53), D => n27, Z => 
                           s_writeback_data_21_port);
   U109 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_22_port, B => n29, C 
                           => mini_mips_i(54), D => n27, Z => 
                           s_writeback_data_22_port);
   U110 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_24_port, B => n29, C 
                           => mini_mips_i(56), D => n27, Z => 
                           s_writeback_data_24_port);
   U111 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_25_port, B => n29, C 
                           => mini_mips_i(57), D => n27, Z => 
                           s_writeback_data_25_port);
   U112 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_29_port, C 
                           => s_exe_in_regA_p_29_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_29_port, Z => s_src_a_29_port);
   U113 : HS65_LH_AO222X4 port map( A => n15, B => s_writeback_data_30_port, C 
                           => s_exe_in_regA_p_30_port, D => n11, E => n5, F => 
                           s_mem_out_alu_res_p_30_port, Z => s_src_a_30_port);
   U114 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_15_port, C 
                           => s_exe_in_regB_p_15_port, D => n20, E => 
                           s_mem_out_alu_res_p_15_port, F => n17, Z => 
                           s_src_b_15_port);
   U115 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_16_port, C 
                           => s_exe_in_regB_p_16_port, D => n20, E => 
                           s_mem_out_alu_res_p_16_port, F => n17, Z => 
                           s_src_b_16_port);
   U116 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_17_port, C 
                           => s_exe_in_regB_p_17_port, D => n20, E => 
                           s_mem_out_alu_res_p_17_port, F => n17, Z => 
                           s_src_b_17_port);
   U117 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_18_port, C 
                           => s_exe_in_regB_p_18_port, D => n20, E => 
                           s_mem_out_alu_res_p_18_port, F => n17, Z => 
                           s_src_b_18_port);
   U118 : HS65_LH_AO222X4 port map( A => n24, B => s_writeback_data_19_port, C 
                           => s_exe_in_regB_p_19_port, D => n20, E => 
                           s_mem_out_alu_res_p_19_port, F => n17, Z => 
                           s_src_b_19_port);
   U119 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_20_port, C 
                           => s_exe_in_regB_p_20_port, D => n21, E => 
                           s_mem_out_alu_res_p_20_port, F => n18, Z => 
                           s_src_b_20_port);
   U120 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_21_port, C 
                           => s_exe_in_regB_p_21_port, D => n21, E => 
                           s_mem_out_alu_res_p_21_port, F => n18, Z => 
                           s_src_b_21_port);
   U121 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_30_port, B => n30, C 
                           => mini_mips_i(62), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_30_port);
   U122 : HS65_LH_AO22X9 port map( A => s_wb_in_alu_res_p_31_port, B => n30, C 
                           => mini_mips_i(63), D => s_wb_in_memtoReg_p, Z => 
                           s_writeback_data_31_port);
   U123 : HS65_LH_AO222X4 port map( A => n16, B => s_writeback_data_31_port, C 
                           => s_exe_in_regA_p_31_port, D => n12, E => n8, F => 
                           s_mem_out_alu_res_p_31_port, Z => s_src_a_31_port);
   U124 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_28_port, C 
                           => s_exe_in_regB_p_28_port, D => n21, E => 
                           s_mem_out_alu_res_p_28_port, F => n18, Z => 
                           s_src_b_28_port);
   U125 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_22_port, C 
                           => s_exe_in_regB_p_22_port, D => n21, E => 
                           s_mem_out_alu_res_p_22_port, F => n18, Z => 
                           s_src_b_22_port);
   U126 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_23_port, C 
                           => s_exe_in_regB_p_23_port, D => n21, E => 
                           s_mem_out_alu_res_p_23_port, F => n18, Z => 
                           s_src_b_23_port);
   U127 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_24_port, C 
                           => s_exe_in_regB_p_24_port, D => n21, E => 
                           s_mem_out_alu_res_p_24_port, F => n18, Z => 
                           s_src_b_24_port);
   U128 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_25_port, C 
                           => s_exe_in_regB_p_25_port, D => n21, E => 
                           s_mem_out_alu_res_p_25_port, F => n18, Z => 
                           s_src_b_25_port);
   U129 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_26_port, C 
                           => s_exe_in_regB_p_26_port, D => n21, E => 
                           s_mem_out_alu_res_p_26_port, F => n18, Z => 
                           s_src_b_26_port);
   U130 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_27_port, C 
                           => s_exe_in_regB_p_27_port, D => n21, E => 
                           s_mem_out_alu_res_p_27_port, F => n18, Z => 
                           s_src_b_27_port);
   U131 : HS65_LH_AO222X4 port map( A => n26, B => s_writeback_data_31_port, C 
                           => s_exe_in_regB_p_31_port, D => n22, E => 
                           s_mem_out_alu_res_p_31_port, F => n19, Z => 
                           s_src_b_31_port);
   U132 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_29_port, C 
                           => s_exe_in_regB_p_29_port, D => n21, E => 
                           s_mem_out_alu_res_p_29_port, F => n18, Z => 
                           s_src_b_29_port);
   U133 : HS65_LH_AO222X4 port map( A => n25, B => s_writeback_data_30_port, C 
                           => s_exe_in_regB_p_30_port, D => n21, E => 
                           s_mem_out_alu_res_p_30_port, F => n18, Z => 
                           s_src_b_30_port);
   U134 : HS65_LH_BFX9 port map( A => rst_n, Z => n32);
   s_ctrl_out_cALU_OP_p_3_port <= '0';

end SYN_Behavioral;

library IEEE,IO65LPHVT_SF_1V8_50A_7M4X0Y2Z,CORE65LPHVT;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity mini_mips_p is

   port( clk, rst_n : inout std_logic);

end mini_mips_p;

architecture SYN_Behavioral of mini_mips_p is

   component mini_mips_pipeline
      port( clk, rst_n : in std_logic;  mini_mips_i : in std_logic_vector (63 
            downto 0);  mini_mips_o : out std_logic_vector (56 downto 0));
   end component;
   
   component BD2SCARUDQP_1V8_SF_LIN
      port( A, TA, TM, EN, TEN : in std_logic;  IO : inout std_logic;  HYST, 
            PDN, PUN : in std_logic;  ZI : out std_logic);
   end component;
   
   component ST_SPHDL_4096x32m8_L
      port( A : in std_logic_vector (11 downto 0);  D : in std_logic_vector (31
            downto 0);  Q : out std_logic_vector (31 downto 0);  CK, CSN : in 
            std_logic;  RY : out std_logic;  TBYPASS, WEN : in std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, clk_i, rst_n_i, 
      s_mini_mips_i_DMEM_DATA_31_port, s_mini_mips_i_DMEM_DATA_30_port, 
      s_mini_mips_i_DMEM_DATA_29_port, s_mini_mips_i_DMEM_DATA_28_port, 
      s_mini_mips_i_DMEM_DATA_27_port, s_mini_mips_i_DMEM_DATA_26_port, 
      s_mini_mips_i_DMEM_DATA_25_port, s_mini_mips_i_DMEM_DATA_24_port, 
      s_mini_mips_i_DMEM_DATA_23_port, s_mini_mips_i_DMEM_DATA_22_port, 
      s_mini_mips_i_DMEM_DATA_21_port, s_mini_mips_i_DMEM_DATA_20_port, 
      s_mini_mips_i_DMEM_DATA_19_port, s_mini_mips_i_DMEM_DATA_18_port, 
      s_mini_mips_i_DMEM_DATA_17_port, s_mini_mips_i_DMEM_DATA_16_port, 
      s_mini_mips_i_DMEM_DATA_15_port, s_mini_mips_i_DMEM_DATA_14_port, 
      s_mini_mips_i_DMEM_DATA_13_port, s_mini_mips_i_DMEM_DATA_12_port, 
      s_mini_mips_i_DMEM_DATA_11_port, s_mini_mips_i_DMEM_DATA_10_port, 
      s_mini_mips_i_DMEM_DATA_9_port, s_mini_mips_i_DMEM_DATA_8_port, 
      s_mini_mips_i_DMEM_DATA_7_port, s_mini_mips_i_DMEM_DATA_6_port, 
      s_mini_mips_i_DMEM_DATA_5_port, s_mini_mips_i_DMEM_DATA_4_port, 
      s_mini_mips_i_DMEM_DATA_3_port, s_mini_mips_i_DMEM_DATA_2_port, 
      s_mini_mips_i_DMEM_DATA_1_port, s_mini_mips_i_DMEM_DATA_0_port, 
      s_mini_mips_i_IMEM_DATA_31_port, s_mini_mips_i_IMEM_DATA_30_port, 
      s_mini_mips_i_IMEM_DATA_29_port, s_mini_mips_i_IMEM_DATA_28_port, 
      s_mini_mips_i_IMEM_DATA_27_port, s_mini_mips_i_IMEM_DATA_26_port, 
      s_mini_mips_i_IMEM_DATA_25_port, s_mini_mips_i_IMEM_DATA_24_port, 
      s_mini_mips_i_IMEM_DATA_23_port, s_mini_mips_i_IMEM_DATA_22_port, 
      s_mini_mips_i_IMEM_DATA_21_port, s_mini_mips_i_IMEM_DATA_20_port, 
      s_mini_mips_i_IMEM_DATA_19_port, s_mini_mips_i_IMEM_DATA_18_port, 
      s_mini_mips_i_IMEM_DATA_17_port, s_mini_mips_i_IMEM_DATA_16_port, 
      s_mini_mips_i_IMEM_DATA_15_port, s_mini_mips_i_IMEM_DATA_14_port, 
      s_mini_mips_i_IMEM_DATA_13_port, s_mini_mips_i_IMEM_DATA_12_port, 
      s_mini_mips_i_IMEM_DATA_11_port, s_mini_mips_i_IMEM_DATA_10_port, 
      s_mini_mips_i_IMEM_DATA_9_port, s_mini_mips_i_IMEM_DATA_8_port, 
      s_mini_mips_i_IMEM_DATA_7_port, s_mini_mips_i_IMEM_DATA_6_port, 
      s_mini_mips_i_IMEM_DATA_5_port, s_mini_mips_i_IMEM_DATA_4_port, 
      s_mini_mips_i_IMEM_DATA_3_port, s_mini_mips_i_IMEM_DATA_2_port, 
      s_mini_mips_i_IMEM_DATA_1_port, s_mini_mips_i_IMEM_DATA_0_port, 
      s_mini_mips_o_DMEM_ADDR_11_port, s_mini_mips_o_DMEM_ADDR_10_port, 
      s_mini_mips_o_DMEM_ADDR_9_port, s_mini_mips_o_DMEM_ADDR_8_port, 
      s_mini_mips_o_DMEM_ADDR_7_port, s_mini_mips_o_DMEM_ADDR_6_port, 
      s_mini_mips_o_DMEM_ADDR_5_port, s_mini_mips_o_DMEM_ADDR_4_port, 
      s_mini_mips_o_DMEM_ADDR_3_port, s_mini_mips_o_DMEM_ADDR_2_port, 
      s_mini_mips_o_DMEM_ADDR_1_port, s_mini_mips_o_DMEM_ADDR_0_port, 
      s_mini_mips_o_IMEM_ADDR_11_port, s_mini_mips_o_IMEM_ADDR_10_port, 
      s_mini_mips_o_IMEM_ADDR_9_port, s_mini_mips_o_IMEM_ADDR_8_port, 
      s_mini_mips_o_IMEM_ADDR_7_port, s_mini_mips_o_IMEM_ADDR_6_port, 
      s_mini_mips_o_IMEM_ADDR_5_port, s_mini_mips_o_IMEM_ADDR_4_port, 
      s_mini_mips_o_IMEM_ADDR_3_port, s_mini_mips_o_IMEM_ADDR_2_port, 
      s_mini_mips_o_IMEM_ADDR_1_port, s_mini_mips_o_IMEM_ADDR_0_port, 
      s_mini_mips_o_DMEM_WEN_N_port, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056 : std_logic;

begin
   
   imem_inst : ST_SPHDL_4096x32m8_L port map( A(11) => 
                           s_mini_mips_o_IMEM_ADDR_11_port, A(10) => 
                           s_mini_mips_o_IMEM_ADDR_10_port, A(9) => 
                           s_mini_mips_o_IMEM_ADDR_9_port, A(8) => 
                           s_mini_mips_o_IMEM_ADDR_8_port, A(7) => 
                           s_mini_mips_o_IMEM_ADDR_7_port, A(6) => 
                           s_mini_mips_o_IMEM_ADDR_6_port, A(5) => 
                           s_mini_mips_o_IMEM_ADDR_5_port, A(4) => 
                           s_mini_mips_o_IMEM_ADDR_4_port, A(3) => 
                           s_mini_mips_o_IMEM_ADDR_3_port, A(2) => 
                           s_mini_mips_o_IMEM_ADDR_2_port, A(1) => 
                           s_mini_mips_o_IMEM_ADDR_1_port, A(0) => 
                           s_mini_mips_o_IMEM_ADDR_0_port, D(31) => 
                           X_Logic0_port, D(30) => X_Logic0_port, D(29) => 
                           X_Logic0_port, D(28) => X_Logic0_port, D(27) => 
                           X_Logic0_port, D(26) => X_Logic0_port, D(25) => 
                           X_Logic0_port, D(24) => X_Logic0_port, D(23) => 
                           X_Logic0_port, D(22) => X_Logic0_port, D(21) => 
                           X_Logic0_port, D(20) => X_Logic0_port, D(19) => 
                           X_Logic0_port, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, Q(31) => 
                           s_mini_mips_i_IMEM_DATA_31_port, Q(30) => 
                           s_mini_mips_i_IMEM_DATA_30_port, Q(29) => 
                           s_mini_mips_i_IMEM_DATA_29_port, Q(28) => 
                           s_mini_mips_i_IMEM_DATA_28_port, Q(27) => 
                           s_mini_mips_i_IMEM_DATA_27_port, Q(26) => 
                           s_mini_mips_i_IMEM_DATA_26_port, Q(25) => 
                           s_mini_mips_i_IMEM_DATA_25_port, Q(24) => 
                           s_mini_mips_i_IMEM_DATA_24_port, Q(23) => 
                           s_mini_mips_i_IMEM_DATA_23_port, Q(22) => 
                           s_mini_mips_i_IMEM_DATA_22_port, Q(21) => 
                           s_mini_mips_i_IMEM_DATA_21_port, Q(20) => 
                           s_mini_mips_i_IMEM_DATA_20_port, Q(19) => 
                           s_mini_mips_i_IMEM_DATA_19_port, Q(18) => 
                           s_mini_mips_i_IMEM_DATA_18_port, Q(17) => 
                           s_mini_mips_i_IMEM_DATA_17_port, Q(16) => 
                           s_mini_mips_i_IMEM_DATA_16_port, Q(15) => 
                           s_mini_mips_i_IMEM_DATA_15_port, Q(14) => 
                           s_mini_mips_i_IMEM_DATA_14_port, Q(13) => 
                           s_mini_mips_i_IMEM_DATA_13_port, Q(12) => 
                           s_mini_mips_i_IMEM_DATA_12_port, Q(11) => 
                           s_mini_mips_i_IMEM_DATA_11_port, Q(10) => 
                           s_mini_mips_i_IMEM_DATA_10_port, Q(9) => 
                           s_mini_mips_i_IMEM_DATA_9_port, Q(8) => 
                           s_mini_mips_i_IMEM_DATA_8_port, Q(7) => 
                           s_mini_mips_i_IMEM_DATA_7_port, Q(6) => 
                           s_mini_mips_i_IMEM_DATA_6_port, Q(5) => 
                           s_mini_mips_i_IMEM_DATA_5_port, Q(4) => 
                           s_mini_mips_i_IMEM_DATA_4_port, Q(3) => 
                           s_mini_mips_i_IMEM_DATA_3_port, Q(2) => 
                           s_mini_mips_i_IMEM_DATA_2_port, Q(1) => 
                           s_mini_mips_i_IMEM_DATA_1_port, Q(0) => 
                           s_mini_mips_i_IMEM_DATA_0_port, CK => clk_i, CSN => 
                           X_Logic0_port, RY => n_1023, TBYPASS => 
                           X_Logic0_port, WEN => X_Logic1_port);
   dmem_inst : ST_SPHDL_4096x32m8_L port map( A(11) => 
                           s_mini_mips_o_DMEM_ADDR_11_port, A(10) => 
                           s_mini_mips_o_DMEM_ADDR_10_port, A(9) => 
                           s_mini_mips_o_DMEM_ADDR_9_port, A(8) => 
                           s_mini_mips_o_DMEM_ADDR_8_port, A(7) => 
                           s_mini_mips_o_DMEM_ADDR_7_port, A(6) => 
                           s_mini_mips_o_DMEM_ADDR_6_port, A(5) => 
                           s_mini_mips_o_DMEM_ADDR_5_port, A(4) => 
                           s_mini_mips_o_DMEM_ADDR_4_port, A(3) => 
                           s_mini_mips_o_DMEM_ADDR_3_port, A(2) => 
                           s_mini_mips_o_DMEM_ADDR_2_port, A(1) => 
                           s_mini_mips_o_DMEM_ADDR_1_port, A(0) => 
                           s_mini_mips_o_DMEM_ADDR_0_port, D(31) => 
                           s_mini_mips_i_DMEM_DATA_31_port, D(30) => 
                           s_mini_mips_i_DMEM_DATA_30_port, D(29) => 
                           s_mini_mips_i_DMEM_DATA_29_port, D(28) => 
                           s_mini_mips_i_DMEM_DATA_28_port, D(27) => 
                           s_mini_mips_i_DMEM_DATA_27_port, D(26) => 
                           s_mini_mips_i_DMEM_DATA_26_port, D(25) => 
                           s_mini_mips_i_DMEM_DATA_25_port, D(24) => 
                           s_mini_mips_i_DMEM_DATA_24_port, D(23) => 
                           s_mini_mips_i_DMEM_DATA_23_port, D(22) => 
                           s_mini_mips_i_DMEM_DATA_22_port, D(21) => 
                           s_mini_mips_i_DMEM_DATA_21_port, D(20) => 
                           s_mini_mips_i_DMEM_DATA_20_port, D(19) => 
                           s_mini_mips_i_DMEM_DATA_19_port, D(18) => 
                           s_mini_mips_i_DMEM_DATA_18_port, D(17) => 
                           s_mini_mips_i_DMEM_DATA_17_port, D(16) => 
                           s_mini_mips_i_DMEM_DATA_16_port, D(15) => 
                           s_mini_mips_i_DMEM_DATA_15_port, D(14) => 
                           s_mini_mips_i_DMEM_DATA_14_port, D(13) => 
                           s_mini_mips_i_DMEM_DATA_13_port, D(12) => 
                           s_mini_mips_i_DMEM_DATA_12_port, D(11) => 
                           s_mini_mips_i_DMEM_DATA_11_port, D(10) => 
                           s_mini_mips_i_DMEM_DATA_10_port, D(9) => 
                           s_mini_mips_i_DMEM_DATA_9_port, D(8) => 
                           s_mini_mips_i_DMEM_DATA_8_port, D(7) => 
                           s_mini_mips_i_DMEM_DATA_7_port, D(6) => 
                           s_mini_mips_i_DMEM_DATA_6_port, D(5) => 
                           s_mini_mips_i_DMEM_DATA_5_port, D(4) => 
                           s_mini_mips_i_DMEM_DATA_4_port, D(3) => 
                           s_mini_mips_i_DMEM_DATA_3_port, D(2) => 
                           s_mini_mips_i_DMEM_DATA_2_port, D(1) => 
                           s_mini_mips_i_DMEM_DATA_1_port, D(0) => 
                           s_mini_mips_i_DMEM_DATA_0_port, Q(31) => 
                           s_mini_mips_i_DMEM_DATA_31_port, Q(30) => 
                           s_mini_mips_i_DMEM_DATA_30_port, Q(29) => 
                           s_mini_mips_i_DMEM_DATA_29_port, Q(28) => 
                           s_mini_mips_i_DMEM_DATA_28_port, Q(27) => 
                           s_mini_mips_i_DMEM_DATA_27_port, Q(26) => 
                           s_mini_mips_i_DMEM_DATA_26_port, Q(25) => 
                           s_mini_mips_i_DMEM_DATA_25_port, Q(24) => 
                           s_mini_mips_i_DMEM_DATA_24_port, Q(23) => 
                           s_mini_mips_i_DMEM_DATA_23_port, Q(22) => 
                           s_mini_mips_i_DMEM_DATA_22_port, Q(21) => 
                           s_mini_mips_i_DMEM_DATA_21_port, Q(20) => 
                           s_mini_mips_i_DMEM_DATA_20_port, Q(19) => 
                           s_mini_mips_i_DMEM_DATA_19_port, Q(18) => 
                           s_mini_mips_i_DMEM_DATA_18_port, Q(17) => 
                           s_mini_mips_i_DMEM_DATA_17_port, Q(16) => 
                           s_mini_mips_i_DMEM_DATA_16_port, Q(15) => 
                           s_mini_mips_i_DMEM_DATA_15_port, Q(14) => 
                           s_mini_mips_i_DMEM_DATA_14_port, Q(13) => 
                           s_mini_mips_i_DMEM_DATA_13_port, Q(12) => 
                           s_mini_mips_i_DMEM_DATA_12_port, Q(11) => 
                           s_mini_mips_i_DMEM_DATA_11_port, Q(10) => 
                           s_mini_mips_i_DMEM_DATA_10_port, Q(9) => 
                           s_mini_mips_i_DMEM_DATA_9_port, Q(8) => 
                           s_mini_mips_i_DMEM_DATA_8_port, Q(7) => 
                           s_mini_mips_i_DMEM_DATA_7_port, Q(6) => 
                           s_mini_mips_i_DMEM_DATA_6_port, Q(5) => 
                           s_mini_mips_i_DMEM_DATA_5_port, Q(4) => 
                           s_mini_mips_i_DMEM_DATA_4_port, Q(3) => 
                           s_mini_mips_i_DMEM_DATA_3_port, Q(2) => 
                           s_mini_mips_i_DMEM_DATA_2_port, Q(1) => 
                           s_mini_mips_i_DMEM_DATA_1_port, Q(0) => 
                           s_mini_mips_i_DMEM_DATA_0_port, CK => clk_i, CSN => 
                           X_Logic0_port, RY => n_1024, TBYPASS => 
                           X_Logic0_port, WEN => s_mini_mips_o_DMEM_WEN_N_port)
                           ;
   clk_pad_in : BD2SCARUDQP_1V8_SF_LIN port map( A => X_Logic0_port, TA => 
                           X_Logic0_port, TM => X_Logic0_port, EN => 
                           X_Logic1_port, TEN => X_Logic1_port, IO => clk, HYST
                           => X_Logic0_port, PDN => X_Logic0_port, PUN => 
                           X_Logic0_port, ZI => clk_i);
   rst_n_pad_in : BD2SCARUDQP_1V8_SF_LIN port map( A => X_Logic0_port, TA => 
                           X_Logic0_port, TM => X_Logic0_port, EN => 
                           X_Logic1_port, TEN => X_Logic1_port, IO => rst_n, 
                           HYST => X_Logic0_port, PDN => X_Logic0_port, PUN => 
                           X_Logic0_port, ZI => rst_n_i);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   mini_mips_inst : mini_mips_pipeline port map( clk => clk_i, rst_n => rst_n_i
                           , mini_mips_i(63) => s_mini_mips_i_DMEM_DATA_31_port
                           , mini_mips_i(62) => s_mini_mips_i_DMEM_DATA_30_port
                           , mini_mips_i(61) => s_mini_mips_i_DMEM_DATA_29_port
                           , mini_mips_i(60) => s_mini_mips_i_DMEM_DATA_28_port
                           , mini_mips_i(59) => s_mini_mips_i_DMEM_DATA_27_port
                           , mini_mips_i(58) => s_mini_mips_i_DMEM_DATA_26_port
                           , mini_mips_i(57) => s_mini_mips_i_DMEM_DATA_25_port
                           , mini_mips_i(56) => s_mini_mips_i_DMEM_DATA_24_port
                           , mini_mips_i(55) => s_mini_mips_i_DMEM_DATA_23_port
                           , mini_mips_i(54) => s_mini_mips_i_DMEM_DATA_22_port
                           , mini_mips_i(53) => s_mini_mips_i_DMEM_DATA_21_port
                           , mini_mips_i(52) => s_mini_mips_i_DMEM_DATA_20_port
                           , mini_mips_i(51) => s_mini_mips_i_DMEM_DATA_19_port
                           , mini_mips_i(50) => s_mini_mips_i_DMEM_DATA_18_port
                           , mini_mips_i(49) => s_mini_mips_i_DMEM_DATA_17_port
                           , mini_mips_i(48) => s_mini_mips_i_DMEM_DATA_16_port
                           , mini_mips_i(47) => s_mini_mips_i_DMEM_DATA_15_port
                           , mini_mips_i(46) => s_mini_mips_i_DMEM_DATA_14_port
                           , mini_mips_i(45) => s_mini_mips_i_DMEM_DATA_13_port
                           , mini_mips_i(44) => s_mini_mips_i_DMEM_DATA_12_port
                           , mini_mips_i(43) => s_mini_mips_i_DMEM_DATA_11_port
                           , mini_mips_i(42) => s_mini_mips_i_DMEM_DATA_10_port
                           , mini_mips_i(41) => s_mini_mips_i_DMEM_DATA_9_port,
                           mini_mips_i(40) => s_mini_mips_i_DMEM_DATA_8_port, 
                           mini_mips_i(39) => s_mini_mips_i_DMEM_DATA_7_port, 
                           mini_mips_i(38) => s_mini_mips_i_DMEM_DATA_6_port, 
                           mini_mips_i(37) => s_mini_mips_i_DMEM_DATA_5_port, 
                           mini_mips_i(36) => s_mini_mips_i_DMEM_DATA_4_port, 
                           mini_mips_i(35) => s_mini_mips_i_DMEM_DATA_3_port, 
                           mini_mips_i(34) => s_mini_mips_i_DMEM_DATA_2_port, 
                           mini_mips_i(33) => s_mini_mips_i_DMEM_DATA_1_port, 
                           mini_mips_i(32) => s_mini_mips_i_DMEM_DATA_0_port, 
                           mini_mips_i(31) => s_mini_mips_i_IMEM_DATA_31_port, 
                           mini_mips_i(30) => s_mini_mips_i_IMEM_DATA_30_port, 
                           mini_mips_i(29) => s_mini_mips_i_IMEM_DATA_29_port, 
                           mini_mips_i(28) => s_mini_mips_i_IMEM_DATA_28_port, 
                           mini_mips_i(27) => s_mini_mips_i_IMEM_DATA_27_port, 
                           mini_mips_i(26) => s_mini_mips_i_IMEM_DATA_26_port, 
                           mini_mips_i(25) => s_mini_mips_i_IMEM_DATA_25_port, 
                           mini_mips_i(24) => s_mini_mips_i_IMEM_DATA_24_port, 
                           mini_mips_i(23) => s_mini_mips_i_IMEM_DATA_23_port, 
                           mini_mips_i(22) => s_mini_mips_i_IMEM_DATA_22_port, 
                           mini_mips_i(21) => s_mini_mips_i_IMEM_DATA_21_port, 
                           mini_mips_i(20) => s_mini_mips_i_IMEM_DATA_20_port, 
                           mini_mips_i(19) => s_mini_mips_i_IMEM_DATA_19_port, 
                           mini_mips_i(18) => s_mini_mips_i_IMEM_DATA_18_port, 
                           mini_mips_i(17) => s_mini_mips_i_IMEM_DATA_17_port, 
                           mini_mips_i(16) => s_mini_mips_i_IMEM_DATA_16_port, 
                           mini_mips_i(15) => s_mini_mips_i_IMEM_DATA_15_port, 
                           mini_mips_i(14) => s_mini_mips_i_IMEM_DATA_14_port, 
                           mini_mips_i(13) => s_mini_mips_i_IMEM_DATA_13_port, 
                           mini_mips_i(12) => s_mini_mips_i_IMEM_DATA_12_port, 
                           mini_mips_i(11) => s_mini_mips_i_IMEM_DATA_11_port, 
                           mini_mips_i(10) => s_mini_mips_i_IMEM_DATA_10_port, 
                           mini_mips_i(9) => s_mini_mips_i_IMEM_DATA_9_port, 
                           mini_mips_i(8) => s_mini_mips_i_IMEM_DATA_8_port, 
                           mini_mips_i(7) => s_mini_mips_i_IMEM_DATA_7_port, 
                           mini_mips_i(6) => s_mini_mips_i_IMEM_DATA_6_port, 
                           mini_mips_i(5) => s_mini_mips_i_IMEM_DATA_5_port, 
                           mini_mips_i(4) => s_mini_mips_i_IMEM_DATA_4_port, 
                           mini_mips_i(3) => s_mini_mips_i_IMEM_DATA_3_port, 
                           mini_mips_i(2) => s_mini_mips_i_IMEM_DATA_2_port, 
                           mini_mips_i(1) => s_mini_mips_i_IMEM_DATA_1_port, 
                           mini_mips_i(0) => s_mini_mips_i_IMEM_DATA_0_port, 
                           mini_mips_o(56) => s_mini_mips_o_DMEM_ADDR_11_port, 
                           mini_mips_o(55) => s_mini_mips_o_DMEM_ADDR_10_port, 
                           mini_mips_o(54) => s_mini_mips_o_DMEM_ADDR_9_port, 
                           mini_mips_o(53) => s_mini_mips_o_DMEM_ADDR_8_port, 
                           mini_mips_o(52) => s_mini_mips_o_DMEM_ADDR_7_port, 
                           mini_mips_o(51) => s_mini_mips_o_DMEM_ADDR_6_port, 
                           mini_mips_o(50) => s_mini_mips_o_DMEM_ADDR_5_port, 
                           mini_mips_o(49) => s_mini_mips_o_DMEM_ADDR_4_port, 
                           mini_mips_o(48) => s_mini_mips_o_DMEM_ADDR_3_port, 
                           mini_mips_o(47) => s_mini_mips_o_DMEM_ADDR_2_port, 
                           mini_mips_o(46) => s_mini_mips_o_DMEM_ADDR_1_port, 
                           mini_mips_o(45) => s_mini_mips_o_DMEM_ADDR_0_port, 
                           mini_mips_o(44) => n_1025, mini_mips_o(43) => n_1026
                           , mini_mips_o(42) => n_1027, mini_mips_o(41) => 
                           n_1028, mini_mips_o(40) => n_1029, mini_mips_o(39) 
                           => n_1030, mini_mips_o(38) => n_1031, 
                           mini_mips_o(37) => n_1032, mini_mips_o(36) => n_1033
                           , mini_mips_o(35) => n_1034, mini_mips_o(34) => 
                           n_1035, mini_mips_o(33) => n_1036, mini_mips_o(32) 
                           => n_1037, mini_mips_o(31) => n_1038, 
                           mini_mips_o(30) => n_1039, mini_mips_o(29) => n_1040
                           , mini_mips_o(28) => n_1041, mini_mips_o(27) => 
                           n_1042, mini_mips_o(26) => n_1043, mini_mips_o(25) 
                           => n_1044, mini_mips_o(24) => n_1045, 
                           mini_mips_o(23) => n_1046, mini_mips_o(22) => n_1047
                           , mini_mips_o(21) => n_1048, mini_mips_o(20) => 
                           n_1049, mini_mips_o(19) => n_1050, mini_mips_o(18) 
                           => n_1051, mini_mips_o(17) => n_1052, 
                           mini_mips_o(16) => n_1053, mini_mips_o(15) => n_1054
                           , mini_mips_o(14) => n_1055, mini_mips_o(13) => 
                           n_1056, mini_mips_o(12) => 
                           s_mini_mips_o_IMEM_ADDR_11_port, mini_mips_o(11) => 
                           s_mini_mips_o_IMEM_ADDR_10_port, mini_mips_o(10) => 
                           s_mini_mips_o_IMEM_ADDR_9_port, mini_mips_o(9) => 
                           s_mini_mips_o_IMEM_ADDR_8_port, mini_mips_o(8) => 
                           s_mini_mips_o_IMEM_ADDR_7_port, mini_mips_o(7) => 
                           s_mini_mips_o_IMEM_ADDR_6_port, mini_mips_o(6) => 
                           s_mini_mips_o_IMEM_ADDR_5_port, mini_mips_o(5) => 
                           s_mini_mips_o_IMEM_ADDR_4_port, mini_mips_o(4) => 
                           s_mini_mips_o_IMEM_ADDR_3_port, mini_mips_o(3) => 
                           s_mini_mips_o_IMEM_ADDR_2_port, mini_mips_o(2) => 
                           s_mini_mips_o_IMEM_ADDR_1_port, mini_mips_o(1) => 
                           s_mini_mips_o_IMEM_ADDR_0_port, mini_mips_o(0) => 
                           s_mini_mips_o_DMEM_WEN_N_port);

end SYN_Behavioral;
